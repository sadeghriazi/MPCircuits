
module psi_BMR_b10000_n4 ( p_input, o );
  input [39999:0] p_input;
  output [9999:0] o;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972,
         n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982,
         n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992,
         n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002,
         n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
         n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022,
         n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032,
         n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042,
         n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052,
         n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062,
         n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072,
         n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082,
         n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092,
         n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102,
         n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112,
         n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122,
         n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132,
         n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142,
         n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152,
         n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162,
         n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172,
         n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182,
         n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192,
         n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202,
         n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212,
         n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222,
         n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232,
         n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242,
         n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252,
         n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262,
         n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272,
         n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282,
         n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292,
         n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302,
         n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312,
         n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322,
         n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332,
         n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342,
         n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352,
         n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362,
         n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372,
         n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382,
         n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392,
         n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402,
         n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412,
         n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422,
         n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432,
         n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442,
         n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452,
         n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
         n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
         n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
         n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
         n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
         n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612,
         n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622,
         n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632,
         n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
         n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652,
         n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662,
         n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672,
         n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682,
         n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692,
         n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702,
         n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712,
         n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722,
         n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732,
         n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742,
         n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752,
         n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762,
         n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772,
         n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782,
         n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792,
         n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802,
         n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812,
         n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822,
         n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832,
         n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842,
         n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852,
         n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862,
         n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872,
         n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882,
         n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892,
         n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902,
         n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912,
         n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922,
         n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932,
         n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942,
         n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952,
         n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962,
         n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972,
         n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982,
         n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992,
         n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002,
         n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012,
         n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022,
         n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032,
         n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042,
         n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052,
         n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062,
         n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072,
         n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082,
         n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092,
         n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102,
         n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112,
         n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122,
         n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132,
         n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142,
         n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152,
         n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162,
         n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172,
         n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182,
         n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192,
         n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202,
         n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212,
         n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222,
         n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232,
         n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242,
         n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252,
         n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262,
         n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272,
         n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282,
         n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292,
         n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302,
         n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312,
         n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322,
         n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332,
         n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342,
         n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352,
         n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362,
         n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372,
         n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382,
         n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392,
         n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402,
         n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412,
         n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422,
         n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432,
         n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442,
         n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452,
         n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462,
         n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472,
         n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482,
         n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492,
         n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502,
         n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512,
         n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522,
         n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532,
         n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542,
         n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552,
         n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562,
         n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572,
         n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582,
         n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592,
         n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602,
         n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612,
         n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622,
         n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632,
         n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642,
         n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652,
         n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662,
         n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672,
         n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682,
         n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692,
         n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702,
         n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712,
         n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722,
         n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732,
         n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742,
         n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752,
         n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762,
         n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772,
         n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782,
         n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792,
         n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802,
         n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812,
         n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822,
         n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832,
         n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842,
         n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852,
         n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862,
         n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872,
         n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882,
         n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892,
         n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902,
         n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912,
         n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922,
         n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932,
         n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942,
         n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952,
         n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962,
         n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972,
         n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982,
         n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992,
         n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002,
         n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012,
         n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022,
         n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032,
         n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042,
         n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052,
         n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062,
         n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072,
         n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082,
         n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092,
         n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102,
         n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112,
         n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122,
         n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132,
         n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142,
         n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152,
         n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162,
         n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172,
         n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182,
         n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192,
         n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202,
         n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212,
         n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222,
         n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232,
         n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242,
         n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252,
         n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262,
         n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272,
         n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282,
         n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292,
         n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302,
         n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312,
         n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322,
         n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332,
         n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342,
         n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352,
         n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362,
         n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372,
         n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382,
         n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392,
         n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402,
         n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412,
         n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422,
         n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432,
         n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442,
         n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452,
         n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462,
         n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472,
         n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482,
         n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492,
         n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502,
         n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512,
         n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522,
         n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532,
         n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542,
         n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552,
         n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562,
         n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572,
         n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582,
         n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592,
         n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602,
         n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612,
         n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622,
         n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632,
         n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642,
         n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652,
         n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662,
         n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672,
         n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682,
         n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692,
         n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702,
         n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712,
         n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722,
         n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732,
         n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742,
         n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752,
         n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762,
         n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772,
         n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782,
         n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792,
         n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802,
         n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812,
         n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822,
         n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832,
         n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842,
         n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852,
         n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862,
         n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872,
         n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882,
         n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892,
         n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902,
         n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912,
         n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922,
         n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932,
         n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942,
         n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952,
         n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962,
         n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972,
         n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982,
         n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992,
         n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002,
         n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012,
         n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022,
         n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032,
         n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042,
         n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052,
         n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062,
         n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072,
         n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082,
         n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092,
         n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102,
         n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112,
         n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122,
         n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132,
         n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142,
         n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152,
         n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162,
         n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172,
         n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182,
         n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192,
         n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202,
         n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212,
         n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222,
         n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232,
         n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242,
         n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252,
         n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262,
         n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272,
         n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282,
         n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292,
         n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302,
         n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312,
         n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322,
         n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332,
         n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342,
         n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352,
         n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362,
         n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372,
         n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382,
         n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392,
         n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402,
         n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412,
         n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422,
         n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432,
         n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442,
         n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452,
         n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462,
         n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472,
         n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482,
         n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492,
         n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502,
         n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512,
         n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522,
         n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532,
         n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542,
         n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552,
         n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562,
         n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572,
         n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582,
         n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592,
         n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602,
         n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612,
         n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622,
         n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632,
         n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642,
         n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652,
         n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662,
         n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672,
         n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682,
         n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692,
         n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702,
         n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712,
         n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722,
         n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732,
         n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742,
         n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752,
         n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762,
         n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772,
         n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782,
         n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792,
         n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802,
         n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812,
         n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822,
         n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832,
         n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842,
         n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852,
         n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862,
         n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872,
         n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882,
         n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892,
         n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902,
         n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912,
         n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922,
         n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932,
         n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942,
         n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952,
         n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962,
         n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972,
         n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982,
         n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992,
         n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002,
         n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012,
         n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022,
         n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032,
         n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042,
         n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052,
         n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062,
         n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072,
         n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082,
         n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092,
         n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102,
         n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112,
         n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122,
         n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132,
         n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142,
         n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152,
         n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162,
         n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172,
         n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182,
         n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192,
         n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202,
         n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212,
         n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222,
         n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232,
         n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242,
         n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252,
         n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262,
         n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272,
         n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282,
         n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292,
         n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302,
         n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312,
         n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322,
         n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332,
         n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342,
         n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352,
         n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362,
         n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372,
         n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382,
         n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392,
         n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402,
         n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412,
         n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422,
         n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432,
         n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442,
         n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452,
         n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462,
         n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472,
         n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482,
         n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492,
         n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502,
         n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512,
         n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522,
         n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532,
         n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542,
         n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552,
         n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562,
         n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572,
         n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582,
         n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592,
         n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602,
         n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612,
         n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622,
         n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632,
         n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642,
         n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652,
         n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662,
         n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672,
         n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682,
         n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692,
         n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702,
         n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712,
         n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722,
         n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732,
         n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742,
         n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752,
         n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762,
         n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772,
         n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782,
         n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792,
         n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802,
         n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812,
         n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822,
         n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832,
         n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842,
         n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852,
         n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862,
         n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872,
         n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882,
         n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892,
         n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902,
         n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912,
         n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922,
         n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932,
         n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942,
         n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952,
         n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962,
         n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972,
         n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982,
         n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992,
         n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002,
         n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012,
         n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022,
         n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032,
         n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042,
         n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052,
         n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062,
         n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072,
         n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082,
         n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092,
         n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102,
         n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112,
         n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122,
         n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132,
         n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142,
         n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152,
         n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162,
         n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172,
         n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182,
         n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192,
         n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202,
         n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212,
         n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222,
         n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232,
         n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242,
         n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252,
         n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262,
         n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272,
         n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282,
         n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292,
         n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302,
         n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312,
         n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322,
         n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332,
         n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342,
         n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352,
         n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362,
         n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372,
         n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382,
         n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392,
         n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402,
         n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412,
         n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422,
         n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432,
         n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442,
         n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452,
         n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462,
         n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472,
         n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482,
         n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492,
         n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502,
         n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512,
         n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522,
         n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532,
         n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542,
         n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552,
         n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562,
         n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572,
         n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582,
         n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592,
         n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602,
         n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612,
         n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622,
         n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632,
         n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642,
         n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652,
         n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662,
         n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672,
         n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682,
         n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692,
         n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702,
         n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712,
         n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722,
         n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732,
         n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742,
         n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752,
         n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762,
         n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772,
         n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782,
         n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792,
         n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802,
         n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812,
         n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822,
         n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832,
         n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842,
         n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852,
         n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862,
         n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872,
         n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882,
         n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892,
         n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902,
         n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912,
         n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922,
         n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932,
         n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942,
         n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952,
         n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962,
         n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972,
         n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982,
         n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992,
         n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001,
         n10002, n10003, n10004, n10005, n10006, n10007, n10008, n10009,
         n10010, n10011, n10012, n10013, n10014, n10015, n10016, n10017,
         n10018, n10019, n10020, n10021, n10022, n10023, n10024, n10025,
         n10026, n10027, n10028, n10029, n10030, n10031, n10032, n10033,
         n10034, n10035, n10036, n10037, n10038, n10039, n10040, n10041,
         n10042, n10043, n10044, n10045, n10046, n10047, n10048, n10049,
         n10050, n10051, n10052, n10053, n10054, n10055, n10056, n10057,
         n10058, n10059, n10060, n10061, n10062, n10063, n10064, n10065,
         n10066, n10067, n10068, n10069, n10070, n10071, n10072, n10073,
         n10074, n10075, n10076, n10077, n10078, n10079, n10080, n10081,
         n10082, n10083, n10084, n10085, n10086, n10087, n10088, n10089,
         n10090, n10091, n10092, n10093, n10094, n10095, n10096, n10097,
         n10098, n10099, n10100, n10101, n10102, n10103, n10104, n10105,
         n10106, n10107, n10108, n10109, n10110, n10111, n10112, n10113,
         n10114, n10115, n10116, n10117, n10118, n10119, n10120, n10121,
         n10122, n10123, n10124, n10125, n10126, n10127, n10128, n10129,
         n10130, n10131, n10132, n10133, n10134, n10135, n10136, n10137,
         n10138, n10139, n10140, n10141, n10142, n10143, n10144, n10145,
         n10146, n10147, n10148, n10149, n10150, n10151, n10152, n10153,
         n10154, n10155, n10156, n10157, n10158, n10159, n10160, n10161,
         n10162, n10163, n10164, n10165, n10166, n10167, n10168, n10169,
         n10170, n10171, n10172, n10173, n10174, n10175, n10176, n10177,
         n10178, n10179, n10180, n10181, n10182, n10183, n10184, n10185,
         n10186, n10187, n10188, n10189, n10190, n10191, n10192, n10193,
         n10194, n10195, n10196, n10197, n10198, n10199, n10200, n10201,
         n10202, n10203, n10204, n10205, n10206, n10207, n10208, n10209,
         n10210, n10211, n10212, n10213, n10214, n10215, n10216, n10217,
         n10218, n10219, n10220, n10221, n10222, n10223, n10224, n10225,
         n10226, n10227, n10228, n10229, n10230, n10231, n10232, n10233,
         n10234, n10235, n10236, n10237, n10238, n10239, n10240, n10241,
         n10242, n10243, n10244, n10245, n10246, n10247, n10248, n10249,
         n10250, n10251, n10252, n10253, n10254, n10255, n10256, n10257,
         n10258, n10259, n10260, n10261, n10262, n10263, n10264, n10265,
         n10266, n10267, n10268, n10269, n10270, n10271, n10272, n10273,
         n10274, n10275, n10276, n10277, n10278, n10279, n10280, n10281,
         n10282, n10283, n10284, n10285, n10286, n10287, n10288, n10289,
         n10290, n10291, n10292, n10293, n10294, n10295, n10296, n10297,
         n10298, n10299, n10300, n10301, n10302, n10303, n10304, n10305,
         n10306, n10307, n10308, n10309, n10310, n10311, n10312, n10313,
         n10314, n10315, n10316, n10317, n10318, n10319, n10320, n10321,
         n10322, n10323, n10324, n10325, n10326, n10327, n10328, n10329,
         n10330, n10331, n10332, n10333, n10334, n10335, n10336, n10337,
         n10338, n10339, n10340, n10341, n10342, n10343, n10344, n10345,
         n10346, n10347, n10348, n10349, n10350, n10351, n10352, n10353,
         n10354, n10355, n10356, n10357, n10358, n10359, n10360, n10361,
         n10362, n10363, n10364, n10365, n10366, n10367, n10368, n10369,
         n10370, n10371, n10372, n10373, n10374, n10375, n10376, n10377,
         n10378, n10379, n10380, n10381, n10382, n10383, n10384, n10385,
         n10386, n10387, n10388, n10389, n10390, n10391, n10392, n10393,
         n10394, n10395, n10396, n10397, n10398, n10399, n10400, n10401,
         n10402, n10403, n10404, n10405, n10406, n10407, n10408, n10409,
         n10410, n10411, n10412, n10413, n10414, n10415, n10416, n10417,
         n10418, n10419, n10420, n10421, n10422, n10423, n10424, n10425,
         n10426, n10427, n10428, n10429, n10430, n10431, n10432, n10433,
         n10434, n10435, n10436, n10437, n10438, n10439, n10440, n10441,
         n10442, n10443, n10444, n10445, n10446, n10447, n10448, n10449,
         n10450, n10451, n10452, n10453, n10454, n10455, n10456, n10457,
         n10458, n10459, n10460, n10461, n10462, n10463, n10464, n10465,
         n10466, n10467, n10468, n10469, n10470, n10471, n10472, n10473,
         n10474, n10475, n10476, n10477, n10478, n10479, n10480, n10481,
         n10482, n10483, n10484, n10485, n10486, n10487, n10488, n10489,
         n10490, n10491, n10492, n10493, n10494, n10495, n10496, n10497,
         n10498, n10499, n10500, n10501, n10502, n10503, n10504, n10505,
         n10506, n10507, n10508, n10509, n10510, n10511, n10512, n10513,
         n10514, n10515, n10516, n10517, n10518, n10519, n10520, n10521,
         n10522, n10523, n10524, n10525, n10526, n10527, n10528, n10529,
         n10530, n10531, n10532, n10533, n10534, n10535, n10536, n10537,
         n10538, n10539, n10540, n10541, n10542, n10543, n10544, n10545,
         n10546, n10547, n10548, n10549, n10550, n10551, n10552, n10553,
         n10554, n10555, n10556, n10557, n10558, n10559, n10560, n10561,
         n10562, n10563, n10564, n10565, n10566, n10567, n10568, n10569,
         n10570, n10571, n10572, n10573, n10574, n10575, n10576, n10577,
         n10578, n10579, n10580, n10581, n10582, n10583, n10584, n10585,
         n10586, n10587, n10588, n10589, n10590, n10591, n10592, n10593,
         n10594, n10595, n10596, n10597, n10598, n10599, n10600, n10601,
         n10602, n10603, n10604, n10605, n10606, n10607, n10608, n10609,
         n10610, n10611, n10612, n10613, n10614, n10615, n10616, n10617,
         n10618, n10619, n10620, n10621, n10622, n10623, n10624, n10625,
         n10626, n10627, n10628, n10629, n10630, n10631, n10632, n10633,
         n10634, n10635, n10636, n10637, n10638, n10639, n10640, n10641,
         n10642, n10643, n10644, n10645, n10646, n10647, n10648, n10649,
         n10650, n10651, n10652, n10653, n10654, n10655, n10656, n10657,
         n10658, n10659, n10660, n10661, n10662, n10663, n10664, n10665,
         n10666, n10667, n10668, n10669, n10670, n10671, n10672, n10673,
         n10674, n10675, n10676, n10677, n10678, n10679, n10680, n10681,
         n10682, n10683, n10684, n10685, n10686, n10687, n10688, n10689,
         n10690, n10691, n10692, n10693, n10694, n10695, n10696, n10697,
         n10698, n10699, n10700, n10701, n10702, n10703, n10704, n10705,
         n10706, n10707, n10708, n10709, n10710, n10711, n10712, n10713,
         n10714, n10715, n10716, n10717, n10718, n10719, n10720, n10721,
         n10722, n10723, n10724, n10725, n10726, n10727, n10728, n10729,
         n10730, n10731, n10732, n10733, n10734, n10735, n10736, n10737,
         n10738, n10739, n10740, n10741, n10742, n10743, n10744, n10745,
         n10746, n10747, n10748, n10749, n10750, n10751, n10752, n10753,
         n10754, n10755, n10756, n10757, n10758, n10759, n10760, n10761,
         n10762, n10763, n10764, n10765, n10766, n10767, n10768, n10769,
         n10770, n10771, n10772, n10773, n10774, n10775, n10776, n10777,
         n10778, n10779, n10780, n10781, n10782, n10783, n10784, n10785,
         n10786, n10787, n10788, n10789, n10790, n10791, n10792, n10793,
         n10794, n10795, n10796, n10797, n10798, n10799, n10800, n10801,
         n10802, n10803, n10804, n10805, n10806, n10807, n10808, n10809,
         n10810, n10811, n10812, n10813, n10814, n10815, n10816, n10817,
         n10818, n10819, n10820, n10821, n10822, n10823, n10824, n10825,
         n10826, n10827, n10828, n10829, n10830, n10831, n10832, n10833,
         n10834, n10835, n10836, n10837, n10838, n10839, n10840, n10841,
         n10842, n10843, n10844, n10845, n10846, n10847, n10848, n10849,
         n10850, n10851, n10852, n10853, n10854, n10855, n10856, n10857,
         n10858, n10859, n10860, n10861, n10862, n10863, n10864, n10865,
         n10866, n10867, n10868, n10869, n10870, n10871, n10872, n10873,
         n10874, n10875, n10876, n10877, n10878, n10879, n10880, n10881,
         n10882, n10883, n10884, n10885, n10886, n10887, n10888, n10889,
         n10890, n10891, n10892, n10893, n10894, n10895, n10896, n10897,
         n10898, n10899, n10900, n10901, n10902, n10903, n10904, n10905,
         n10906, n10907, n10908, n10909, n10910, n10911, n10912, n10913,
         n10914, n10915, n10916, n10917, n10918, n10919, n10920, n10921,
         n10922, n10923, n10924, n10925, n10926, n10927, n10928, n10929,
         n10930, n10931, n10932, n10933, n10934, n10935, n10936, n10937,
         n10938, n10939, n10940, n10941, n10942, n10943, n10944, n10945,
         n10946, n10947, n10948, n10949, n10950, n10951, n10952, n10953,
         n10954, n10955, n10956, n10957, n10958, n10959, n10960, n10961,
         n10962, n10963, n10964, n10965, n10966, n10967, n10968, n10969,
         n10970, n10971, n10972, n10973, n10974, n10975, n10976, n10977,
         n10978, n10979, n10980, n10981, n10982, n10983, n10984, n10985,
         n10986, n10987, n10988, n10989, n10990, n10991, n10992, n10993,
         n10994, n10995, n10996, n10997, n10998, n10999, n11000, n11001,
         n11002, n11003, n11004, n11005, n11006, n11007, n11008, n11009,
         n11010, n11011, n11012, n11013, n11014, n11015, n11016, n11017,
         n11018, n11019, n11020, n11021, n11022, n11023, n11024, n11025,
         n11026, n11027, n11028, n11029, n11030, n11031, n11032, n11033,
         n11034, n11035, n11036, n11037, n11038, n11039, n11040, n11041,
         n11042, n11043, n11044, n11045, n11046, n11047, n11048, n11049,
         n11050, n11051, n11052, n11053, n11054, n11055, n11056, n11057,
         n11058, n11059, n11060, n11061, n11062, n11063, n11064, n11065,
         n11066, n11067, n11068, n11069, n11070, n11071, n11072, n11073,
         n11074, n11075, n11076, n11077, n11078, n11079, n11080, n11081,
         n11082, n11083, n11084, n11085, n11086, n11087, n11088, n11089,
         n11090, n11091, n11092, n11093, n11094, n11095, n11096, n11097,
         n11098, n11099, n11100, n11101, n11102, n11103, n11104, n11105,
         n11106, n11107, n11108, n11109, n11110, n11111, n11112, n11113,
         n11114, n11115, n11116, n11117, n11118, n11119, n11120, n11121,
         n11122, n11123, n11124, n11125, n11126, n11127, n11128, n11129,
         n11130, n11131, n11132, n11133, n11134, n11135, n11136, n11137,
         n11138, n11139, n11140, n11141, n11142, n11143, n11144, n11145,
         n11146, n11147, n11148, n11149, n11150, n11151, n11152, n11153,
         n11154, n11155, n11156, n11157, n11158, n11159, n11160, n11161,
         n11162, n11163, n11164, n11165, n11166, n11167, n11168, n11169,
         n11170, n11171, n11172, n11173, n11174, n11175, n11176, n11177,
         n11178, n11179, n11180, n11181, n11182, n11183, n11184, n11185,
         n11186, n11187, n11188, n11189, n11190, n11191, n11192, n11193,
         n11194, n11195, n11196, n11197, n11198, n11199, n11200, n11201,
         n11202, n11203, n11204, n11205, n11206, n11207, n11208, n11209,
         n11210, n11211, n11212, n11213, n11214, n11215, n11216, n11217,
         n11218, n11219, n11220, n11221, n11222, n11223, n11224, n11225,
         n11226, n11227, n11228, n11229, n11230, n11231, n11232, n11233,
         n11234, n11235, n11236, n11237, n11238, n11239, n11240, n11241,
         n11242, n11243, n11244, n11245, n11246, n11247, n11248, n11249,
         n11250, n11251, n11252, n11253, n11254, n11255, n11256, n11257,
         n11258, n11259, n11260, n11261, n11262, n11263, n11264, n11265,
         n11266, n11267, n11268, n11269, n11270, n11271, n11272, n11273,
         n11274, n11275, n11276, n11277, n11278, n11279, n11280, n11281,
         n11282, n11283, n11284, n11285, n11286, n11287, n11288, n11289,
         n11290, n11291, n11292, n11293, n11294, n11295, n11296, n11297,
         n11298, n11299, n11300, n11301, n11302, n11303, n11304, n11305,
         n11306, n11307, n11308, n11309, n11310, n11311, n11312, n11313,
         n11314, n11315, n11316, n11317, n11318, n11319, n11320, n11321,
         n11322, n11323, n11324, n11325, n11326, n11327, n11328, n11329,
         n11330, n11331, n11332, n11333, n11334, n11335, n11336, n11337,
         n11338, n11339, n11340, n11341, n11342, n11343, n11344, n11345,
         n11346, n11347, n11348, n11349, n11350, n11351, n11352, n11353,
         n11354, n11355, n11356, n11357, n11358, n11359, n11360, n11361,
         n11362, n11363, n11364, n11365, n11366, n11367, n11368, n11369,
         n11370, n11371, n11372, n11373, n11374, n11375, n11376, n11377,
         n11378, n11379, n11380, n11381, n11382, n11383, n11384, n11385,
         n11386, n11387, n11388, n11389, n11390, n11391, n11392, n11393,
         n11394, n11395, n11396, n11397, n11398, n11399, n11400, n11401,
         n11402, n11403, n11404, n11405, n11406, n11407, n11408, n11409,
         n11410, n11411, n11412, n11413, n11414, n11415, n11416, n11417,
         n11418, n11419, n11420, n11421, n11422, n11423, n11424, n11425,
         n11426, n11427, n11428, n11429, n11430, n11431, n11432, n11433,
         n11434, n11435, n11436, n11437, n11438, n11439, n11440, n11441,
         n11442, n11443, n11444, n11445, n11446, n11447, n11448, n11449,
         n11450, n11451, n11452, n11453, n11454, n11455, n11456, n11457,
         n11458, n11459, n11460, n11461, n11462, n11463, n11464, n11465,
         n11466, n11467, n11468, n11469, n11470, n11471, n11472, n11473,
         n11474, n11475, n11476, n11477, n11478, n11479, n11480, n11481,
         n11482, n11483, n11484, n11485, n11486, n11487, n11488, n11489,
         n11490, n11491, n11492, n11493, n11494, n11495, n11496, n11497,
         n11498, n11499, n11500, n11501, n11502, n11503, n11504, n11505,
         n11506, n11507, n11508, n11509, n11510, n11511, n11512, n11513,
         n11514, n11515, n11516, n11517, n11518, n11519, n11520, n11521,
         n11522, n11523, n11524, n11525, n11526, n11527, n11528, n11529,
         n11530, n11531, n11532, n11533, n11534, n11535, n11536, n11537,
         n11538, n11539, n11540, n11541, n11542, n11543, n11544, n11545,
         n11546, n11547, n11548, n11549, n11550, n11551, n11552, n11553,
         n11554, n11555, n11556, n11557, n11558, n11559, n11560, n11561,
         n11562, n11563, n11564, n11565, n11566, n11567, n11568, n11569,
         n11570, n11571, n11572, n11573, n11574, n11575, n11576, n11577,
         n11578, n11579, n11580, n11581, n11582, n11583, n11584, n11585,
         n11586, n11587, n11588, n11589, n11590, n11591, n11592, n11593,
         n11594, n11595, n11596, n11597, n11598, n11599, n11600, n11601,
         n11602, n11603, n11604, n11605, n11606, n11607, n11608, n11609,
         n11610, n11611, n11612, n11613, n11614, n11615, n11616, n11617,
         n11618, n11619, n11620, n11621, n11622, n11623, n11624, n11625,
         n11626, n11627, n11628, n11629, n11630, n11631, n11632, n11633,
         n11634, n11635, n11636, n11637, n11638, n11639, n11640, n11641,
         n11642, n11643, n11644, n11645, n11646, n11647, n11648, n11649,
         n11650, n11651, n11652, n11653, n11654, n11655, n11656, n11657,
         n11658, n11659, n11660, n11661, n11662, n11663, n11664, n11665,
         n11666, n11667, n11668, n11669, n11670, n11671, n11672, n11673,
         n11674, n11675, n11676, n11677, n11678, n11679, n11680, n11681,
         n11682, n11683, n11684, n11685, n11686, n11687, n11688, n11689,
         n11690, n11691, n11692, n11693, n11694, n11695, n11696, n11697,
         n11698, n11699, n11700, n11701, n11702, n11703, n11704, n11705,
         n11706, n11707, n11708, n11709, n11710, n11711, n11712, n11713,
         n11714, n11715, n11716, n11717, n11718, n11719, n11720, n11721,
         n11722, n11723, n11724, n11725, n11726, n11727, n11728, n11729,
         n11730, n11731, n11732, n11733, n11734, n11735, n11736, n11737,
         n11738, n11739, n11740, n11741, n11742, n11743, n11744, n11745,
         n11746, n11747, n11748, n11749, n11750, n11751, n11752, n11753,
         n11754, n11755, n11756, n11757, n11758, n11759, n11760, n11761,
         n11762, n11763, n11764, n11765, n11766, n11767, n11768, n11769,
         n11770, n11771, n11772, n11773, n11774, n11775, n11776, n11777,
         n11778, n11779, n11780, n11781, n11782, n11783, n11784, n11785,
         n11786, n11787, n11788, n11789, n11790, n11791, n11792, n11793,
         n11794, n11795, n11796, n11797, n11798, n11799, n11800, n11801,
         n11802, n11803, n11804, n11805, n11806, n11807, n11808, n11809,
         n11810, n11811, n11812, n11813, n11814, n11815, n11816, n11817,
         n11818, n11819, n11820, n11821, n11822, n11823, n11824, n11825,
         n11826, n11827, n11828, n11829, n11830, n11831, n11832, n11833,
         n11834, n11835, n11836, n11837, n11838, n11839, n11840, n11841,
         n11842, n11843, n11844, n11845, n11846, n11847, n11848, n11849,
         n11850, n11851, n11852, n11853, n11854, n11855, n11856, n11857,
         n11858, n11859, n11860, n11861, n11862, n11863, n11864, n11865,
         n11866, n11867, n11868, n11869, n11870, n11871, n11872, n11873,
         n11874, n11875, n11876, n11877, n11878, n11879, n11880, n11881,
         n11882, n11883, n11884, n11885, n11886, n11887, n11888, n11889,
         n11890, n11891, n11892, n11893, n11894, n11895, n11896, n11897,
         n11898, n11899, n11900, n11901, n11902, n11903, n11904, n11905,
         n11906, n11907, n11908, n11909, n11910, n11911, n11912, n11913,
         n11914, n11915, n11916, n11917, n11918, n11919, n11920, n11921,
         n11922, n11923, n11924, n11925, n11926, n11927, n11928, n11929,
         n11930, n11931, n11932, n11933, n11934, n11935, n11936, n11937,
         n11938, n11939, n11940, n11941, n11942, n11943, n11944, n11945,
         n11946, n11947, n11948, n11949, n11950, n11951, n11952, n11953,
         n11954, n11955, n11956, n11957, n11958, n11959, n11960, n11961,
         n11962, n11963, n11964, n11965, n11966, n11967, n11968, n11969,
         n11970, n11971, n11972, n11973, n11974, n11975, n11976, n11977,
         n11978, n11979, n11980, n11981, n11982, n11983, n11984, n11985,
         n11986, n11987, n11988, n11989, n11990, n11991, n11992, n11993,
         n11994, n11995, n11996, n11997, n11998, n11999, n12000, n12001,
         n12002, n12003, n12004, n12005, n12006, n12007, n12008, n12009,
         n12010, n12011, n12012, n12013, n12014, n12015, n12016, n12017,
         n12018, n12019, n12020, n12021, n12022, n12023, n12024, n12025,
         n12026, n12027, n12028, n12029, n12030, n12031, n12032, n12033,
         n12034, n12035, n12036, n12037, n12038, n12039, n12040, n12041,
         n12042, n12043, n12044, n12045, n12046, n12047, n12048, n12049,
         n12050, n12051, n12052, n12053, n12054, n12055, n12056, n12057,
         n12058, n12059, n12060, n12061, n12062, n12063, n12064, n12065,
         n12066, n12067, n12068, n12069, n12070, n12071, n12072, n12073,
         n12074, n12075, n12076, n12077, n12078, n12079, n12080, n12081,
         n12082, n12083, n12084, n12085, n12086, n12087, n12088, n12089,
         n12090, n12091, n12092, n12093, n12094, n12095, n12096, n12097,
         n12098, n12099, n12100, n12101, n12102, n12103, n12104, n12105,
         n12106, n12107, n12108, n12109, n12110, n12111, n12112, n12113,
         n12114, n12115, n12116, n12117, n12118, n12119, n12120, n12121,
         n12122, n12123, n12124, n12125, n12126, n12127, n12128, n12129,
         n12130, n12131, n12132, n12133, n12134, n12135, n12136, n12137,
         n12138, n12139, n12140, n12141, n12142, n12143, n12144, n12145,
         n12146, n12147, n12148, n12149, n12150, n12151, n12152, n12153,
         n12154, n12155, n12156, n12157, n12158, n12159, n12160, n12161,
         n12162, n12163, n12164, n12165, n12166, n12167, n12168, n12169,
         n12170, n12171, n12172, n12173, n12174, n12175, n12176, n12177,
         n12178, n12179, n12180, n12181, n12182, n12183, n12184, n12185,
         n12186, n12187, n12188, n12189, n12190, n12191, n12192, n12193,
         n12194, n12195, n12196, n12197, n12198, n12199, n12200, n12201,
         n12202, n12203, n12204, n12205, n12206, n12207, n12208, n12209,
         n12210, n12211, n12212, n12213, n12214, n12215, n12216, n12217,
         n12218, n12219, n12220, n12221, n12222, n12223, n12224, n12225,
         n12226, n12227, n12228, n12229, n12230, n12231, n12232, n12233,
         n12234, n12235, n12236, n12237, n12238, n12239, n12240, n12241,
         n12242, n12243, n12244, n12245, n12246, n12247, n12248, n12249,
         n12250, n12251, n12252, n12253, n12254, n12255, n12256, n12257,
         n12258, n12259, n12260, n12261, n12262, n12263, n12264, n12265,
         n12266, n12267, n12268, n12269, n12270, n12271, n12272, n12273,
         n12274, n12275, n12276, n12277, n12278, n12279, n12280, n12281,
         n12282, n12283, n12284, n12285, n12286, n12287, n12288, n12289,
         n12290, n12291, n12292, n12293, n12294, n12295, n12296, n12297,
         n12298, n12299, n12300, n12301, n12302, n12303, n12304, n12305,
         n12306, n12307, n12308, n12309, n12310, n12311, n12312, n12313,
         n12314, n12315, n12316, n12317, n12318, n12319, n12320, n12321,
         n12322, n12323, n12324, n12325, n12326, n12327, n12328, n12329,
         n12330, n12331, n12332, n12333, n12334, n12335, n12336, n12337,
         n12338, n12339, n12340, n12341, n12342, n12343, n12344, n12345,
         n12346, n12347, n12348, n12349, n12350, n12351, n12352, n12353,
         n12354, n12355, n12356, n12357, n12358, n12359, n12360, n12361,
         n12362, n12363, n12364, n12365, n12366, n12367, n12368, n12369,
         n12370, n12371, n12372, n12373, n12374, n12375, n12376, n12377,
         n12378, n12379, n12380, n12381, n12382, n12383, n12384, n12385,
         n12386, n12387, n12388, n12389, n12390, n12391, n12392, n12393,
         n12394, n12395, n12396, n12397, n12398, n12399, n12400, n12401,
         n12402, n12403, n12404, n12405, n12406, n12407, n12408, n12409,
         n12410, n12411, n12412, n12413, n12414, n12415, n12416, n12417,
         n12418, n12419, n12420, n12421, n12422, n12423, n12424, n12425,
         n12426, n12427, n12428, n12429, n12430, n12431, n12432, n12433,
         n12434, n12435, n12436, n12437, n12438, n12439, n12440, n12441,
         n12442, n12443, n12444, n12445, n12446, n12447, n12448, n12449,
         n12450, n12451, n12452, n12453, n12454, n12455, n12456, n12457,
         n12458, n12459, n12460, n12461, n12462, n12463, n12464, n12465,
         n12466, n12467, n12468, n12469, n12470, n12471, n12472, n12473,
         n12474, n12475, n12476, n12477, n12478, n12479, n12480, n12481,
         n12482, n12483, n12484, n12485, n12486, n12487, n12488, n12489,
         n12490, n12491, n12492, n12493, n12494, n12495, n12496, n12497,
         n12498, n12499, n12500, n12501, n12502, n12503, n12504, n12505,
         n12506, n12507, n12508, n12509, n12510, n12511, n12512, n12513,
         n12514, n12515, n12516, n12517, n12518, n12519, n12520, n12521,
         n12522, n12523, n12524, n12525, n12526, n12527, n12528, n12529,
         n12530, n12531, n12532, n12533, n12534, n12535, n12536, n12537,
         n12538, n12539, n12540, n12541, n12542, n12543, n12544, n12545,
         n12546, n12547, n12548, n12549, n12550, n12551, n12552, n12553,
         n12554, n12555, n12556, n12557, n12558, n12559, n12560, n12561,
         n12562, n12563, n12564, n12565, n12566, n12567, n12568, n12569,
         n12570, n12571, n12572, n12573, n12574, n12575, n12576, n12577,
         n12578, n12579, n12580, n12581, n12582, n12583, n12584, n12585,
         n12586, n12587, n12588, n12589, n12590, n12591, n12592, n12593,
         n12594, n12595, n12596, n12597, n12598, n12599, n12600, n12601,
         n12602, n12603, n12604, n12605, n12606, n12607, n12608, n12609,
         n12610, n12611, n12612, n12613, n12614, n12615, n12616, n12617,
         n12618, n12619, n12620, n12621, n12622, n12623, n12624, n12625,
         n12626, n12627, n12628, n12629, n12630, n12631, n12632, n12633,
         n12634, n12635, n12636, n12637, n12638, n12639, n12640, n12641,
         n12642, n12643, n12644, n12645, n12646, n12647, n12648, n12649,
         n12650, n12651, n12652, n12653, n12654, n12655, n12656, n12657,
         n12658, n12659, n12660, n12661, n12662, n12663, n12664, n12665,
         n12666, n12667, n12668, n12669, n12670, n12671, n12672, n12673,
         n12674, n12675, n12676, n12677, n12678, n12679, n12680, n12681,
         n12682, n12683, n12684, n12685, n12686, n12687, n12688, n12689,
         n12690, n12691, n12692, n12693, n12694, n12695, n12696, n12697,
         n12698, n12699, n12700, n12701, n12702, n12703, n12704, n12705,
         n12706, n12707, n12708, n12709, n12710, n12711, n12712, n12713,
         n12714, n12715, n12716, n12717, n12718, n12719, n12720, n12721,
         n12722, n12723, n12724, n12725, n12726, n12727, n12728, n12729,
         n12730, n12731, n12732, n12733, n12734, n12735, n12736, n12737,
         n12738, n12739, n12740, n12741, n12742, n12743, n12744, n12745,
         n12746, n12747, n12748, n12749, n12750, n12751, n12752, n12753,
         n12754, n12755, n12756, n12757, n12758, n12759, n12760, n12761,
         n12762, n12763, n12764, n12765, n12766, n12767, n12768, n12769,
         n12770, n12771, n12772, n12773, n12774, n12775, n12776, n12777,
         n12778, n12779, n12780, n12781, n12782, n12783, n12784, n12785,
         n12786, n12787, n12788, n12789, n12790, n12791, n12792, n12793,
         n12794, n12795, n12796, n12797, n12798, n12799, n12800, n12801,
         n12802, n12803, n12804, n12805, n12806, n12807, n12808, n12809,
         n12810, n12811, n12812, n12813, n12814, n12815, n12816, n12817,
         n12818, n12819, n12820, n12821, n12822, n12823, n12824, n12825,
         n12826, n12827, n12828, n12829, n12830, n12831, n12832, n12833,
         n12834, n12835, n12836, n12837, n12838, n12839, n12840, n12841,
         n12842, n12843, n12844, n12845, n12846, n12847, n12848, n12849,
         n12850, n12851, n12852, n12853, n12854, n12855, n12856, n12857,
         n12858, n12859, n12860, n12861, n12862, n12863, n12864, n12865,
         n12866, n12867, n12868, n12869, n12870, n12871, n12872, n12873,
         n12874, n12875, n12876, n12877, n12878, n12879, n12880, n12881,
         n12882, n12883, n12884, n12885, n12886, n12887, n12888, n12889,
         n12890, n12891, n12892, n12893, n12894, n12895, n12896, n12897,
         n12898, n12899, n12900, n12901, n12902, n12903, n12904, n12905,
         n12906, n12907, n12908, n12909, n12910, n12911, n12912, n12913,
         n12914, n12915, n12916, n12917, n12918, n12919, n12920, n12921,
         n12922, n12923, n12924, n12925, n12926, n12927, n12928, n12929,
         n12930, n12931, n12932, n12933, n12934, n12935, n12936, n12937,
         n12938, n12939, n12940, n12941, n12942, n12943, n12944, n12945,
         n12946, n12947, n12948, n12949, n12950, n12951, n12952, n12953,
         n12954, n12955, n12956, n12957, n12958, n12959, n12960, n12961,
         n12962, n12963, n12964, n12965, n12966, n12967, n12968, n12969,
         n12970, n12971, n12972, n12973, n12974, n12975, n12976, n12977,
         n12978, n12979, n12980, n12981, n12982, n12983, n12984, n12985,
         n12986, n12987, n12988, n12989, n12990, n12991, n12992, n12993,
         n12994, n12995, n12996, n12997, n12998, n12999, n13000, n13001,
         n13002, n13003, n13004, n13005, n13006, n13007, n13008, n13009,
         n13010, n13011, n13012, n13013, n13014, n13015, n13016, n13017,
         n13018, n13019, n13020, n13021, n13022, n13023, n13024, n13025,
         n13026, n13027, n13028, n13029, n13030, n13031, n13032, n13033,
         n13034, n13035, n13036, n13037, n13038, n13039, n13040, n13041,
         n13042, n13043, n13044, n13045, n13046, n13047, n13048, n13049,
         n13050, n13051, n13052, n13053, n13054, n13055, n13056, n13057,
         n13058, n13059, n13060, n13061, n13062, n13063, n13064, n13065,
         n13066, n13067, n13068, n13069, n13070, n13071, n13072, n13073,
         n13074, n13075, n13076, n13077, n13078, n13079, n13080, n13081,
         n13082, n13083, n13084, n13085, n13086, n13087, n13088, n13089,
         n13090, n13091, n13092, n13093, n13094, n13095, n13096, n13097,
         n13098, n13099, n13100, n13101, n13102, n13103, n13104, n13105,
         n13106, n13107, n13108, n13109, n13110, n13111, n13112, n13113,
         n13114, n13115, n13116, n13117, n13118, n13119, n13120, n13121,
         n13122, n13123, n13124, n13125, n13126, n13127, n13128, n13129,
         n13130, n13131, n13132, n13133, n13134, n13135, n13136, n13137,
         n13138, n13139, n13140, n13141, n13142, n13143, n13144, n13145,
         n13146, n13147, n13148, n13149, n13150, n13151, n13152, n13153,
         n13154, n13155, n13156, n13157, n13158, n13159, n13160, n13161,
         n13162, n13163, n13164, n13165, n13166, n13167, n13168, n13169,
         n13170, n13171, n13172, n13173, n13174, n13175, n13176, n13177,
         n13178, n13179, n13180, n13181, n13182, n13183, n13184, n13185,
         n13186, n13187, n13188, n13189, n13190, n13191, n13192, n13193,
         n13194, n13195, n13196, n13197, n13198, n13199, n13200, n13201,
         n13202, n13203, n13204, n13205, n13206, n13207, n13208, n13209,
         n13210, n13211, n13212, n13213, n13214, n13215, n13216, n13217,
         n13218, n13219, n13220, n13221, n13222, n13223, n13224, n13225,
         n13226, n13227, n13228, n13229, n13230, n13231, n13232, n13233,
         n13234, n13235, n13236, n13237, n13238, n13239, n13240, n13241,
         n13242, n13243, n13244, n13245, n13246, n13247, n13248, n13249,
         n13250, n13251, n13252, n13253, n13254, n13255, n13256, n13257,
         n13258, n13259, n13260, n13261, n13262, n13263, n13264, n13265,
         n13266, n13267, n13268, n13269, n13270, n13271, n13272, n13273,
         n13274, n13275, n13276, n13277, n13278, n13279, n13280, n13281,
         n13282, n13283, n13284, n13285, n13286, n13287, n13288, n13289,
         n13290, n13291, n13292, n13293, n13294, n13295, n13296, n13297,
         n13298, n13299, n13300, n13301, n13302, n13303, n13304, n13305,
         n13306, n13307, n13308, n13309, n13310, n13311, n13312, n13313,
         n13314, n13315, n13316, n13317, n13318, n13319, n13320, n13321,
         n13322, n13323, n13324, n13325, n13326, n13327, n13328, n13329,
         n13330, n13331, n13332, n13333, n13334, n13335, n13336, n13337,
         n13338, n13339, n13340, n13341, n13342, n13343, n13344, n13345,
         n13346, n13347, n13348, n13349, n13350, n13351, n13352, n13353,
         n13354, n13355, n13356, n13357, n13358, n13359, n13360, n13361,
         n13362, n13363, n13364, n13365, n13366, n13367, n13368, n13369,
         n13370, n13371, n13372, n13373, n13374, n13375, n13376, n13377,
         n13378, n13379, n13380, n13381, n13382, n13383, n13384, n13385,
         n13386, n13387, n13388, n13389, n13390, n13391, n13392, n13393,
         n13394, n13395, n13396, n13397, n13398, n13399, n13400, n13401,
         n13402, n13403, n13404, n13405, n13406, n13407, n13408, n13409,
         n13410, n13411, n13412, n13413, n13414, n13415, n13416, n13417,
         n13418, n13419, n13420, n13421, n13422, n13423, n13424, n13425,
         n13426, n13427, n13428, n13429, n13430, n13431, n13432, n13433,
         n13434, n13435, n13436, n13437, n13438, n13439, n13440, n13441,
         n13442, n13443, n13444, n13445, n13446, n13447, n13448, n13449,
         n13450, n13451, n13452, n13453, n13454, n13455, n13456, n13457,
         n13458, n13459, n13460, n13461, n13462, n13463, n13464, n13465,
         n13466, n13467, n13468, n13469, n13470, n13471, n13472, n13473,
         n13474, n13475, n13476, n13477, n13478, n13479, n13480, n13481,
         n13482, n13483, n13484, n13485, n13486, n13487, n13488, n13489,
         n13490, n13491, n13492, n13493, n13494, n13495, n13496, n13497,
         n13498, n13499, n13500, n13501, n13502, n13503, n13504, n13505,
         n13506, n13507, n13508, n13509, n13510, n13511, n13512, n13513,
         n13514, n13515, n13516, n13517, n13518, n13519, n13520, n13521,
         n13522, n13523, n13524, n13525, n13526, n13527, n13528, n13529,
         n13530, n13531, n13532, n13533, n13534, n13535, n13536, n13537,
         n13538, n13539, n13540, n13541, n13542, n13543, n13544, n13545,
         n13546, n13547, n13548, n13549, n13550, n13551, n13552, n13553,
         n13554, n13555, n13556, n13557, n13558, n13559, n13560, n13561,
         n13562, n13563, n13564, n13565, n13566, n13567, n13568, n13569,
         n13570, n13571, n13572, n13573, n13574, n13575, n13576, n13577,
         n13578, n13579, n13580, n13581, n13582, n13583, n13584, n13585,
         n13586, n13587, n13588, n13589, n13590, n13591, n13592, n13593,
         n13594, n13595, n13596, n13597, n13598, n13599, n13600, n13601,
         n13602, n13603, n13604, n13605, n13606, n13607, n13608, n13609,
         n13610, n13611, n13612, n13613, n13614, n13615, n13616, n13617,
         n13618, n13619, n13620, n13621, n13622, n13623, n13624, n13625,
         n13626, n13627, n13628, n13629, n13630, n13631, n13632, n13633,
         n13634, n13635, n13636, n13637, n13638, n13639, n13640, n13641,
         n13642, n13643, n13644, n13645, n13646, n13647, n13648, n13649,
         n13650, n13651, n13652, n13653, n13654, n13655, n13656, n13657,
         n13658, n13659, n13660, n13661, n13662, n13663, n13664, n13665,
         n13666, n13667, n13668, n13669, n13670, n13671, n13672, n13673,
         n13674, n13675, n13676, n13677, n13678, n13679, n13680, n13681,
         n13682, n13683, n13684, n13685, n13686, n13687, n13688, n13689,
         n13690, n13691, n13692, n13693, n13694, n13695, n13696, n13697,
         n13698, n13699, n13700, n13701, n13702, n13703, n13704, n13705,
         n13706, n13707, n13708, n13709, n13710, n13711, n13712, n13713,
         n13714, n13715, n13716, n13717, n13718, n13719, n13720, n13721,
         n13722, n13723, n13724, n13725, n13726, n13727, n13728, n13729,
         n13730, n13731, n13732, n13733, n13734, n13735, n13736, n13737,
         n13738, n13739, n13740, n13741, n13742, n13743, n13744, n13745,
         n13746, n13747, n13748, n13749, n13750, n13751, n13752, n13753,
         n13754, n13755, n13756, n13757, n13758, n13759, n13760, n13761,
         n13762, n13763, n13764, n13765, n13766, n13767, n13768, n13769,
         n13770, n13771, n13772, n13773, n13774, n13775, n13776, n13777,
         n13778, n13779, n13780, n13781, n13782, n13783, n13784, n13785,
         n13786, n13787, n13788, n13789, n13790, n13791, n13792, n13793,
         n13794, n13795, n13796, n13797, n13798, n13799, n13800, n13801,
         n13802, n13803, n13804, n13805, n13806, n13807, n13808, n13809,
         n13810, n13811, n13812, n13813, n13814, n13815, n13816, n13817,
         n13818, n13819, n13820, n13821, n13822, n13823, n13824, n13825,
         n13826, n13827, n13828, n13829, n13830, n13831, n13832, n13833,
         n13834, n13835, n13836, n13837, n13838, n13839, n13840, n13841,
         n13842, n13843, n13844, n13845, n13846, n13847, n13848, n13849,
         n13850, n13851, n13852, n13853, n13854, n13855, n13856, n13857,
         n13858, n13859, n13860, n13861, n13862, n13863, n13864, n13865,
         n13866, n13867, n13868, n13869, n13870, n13871, n13872, n13873,
         n13874, n13875, n13876, n13877, n13878, n13879, n13880, n13881,
         n13882, n13883, n13884, n13885, n13886, n13887, n13888, n13889,
         n13890, n13891, n13892, n13893, n13894, n13895, n13896, n13897,
         n13898, n13899, n13900, n13901, n13902, n13903, n13904, n13905,
         n13906, n13907, n13908, n13909, n13910, n13911, n13912, n13913,
         n13914, n13915, n13916, n13917, n13918, n13919, n13920, n13921,
         n13922, n13923, n13924, n13925, n13926, n13927, n13928, n13929,
         n13930, n13931, n13932, n13933, n13934, n13935, n13936, n13937,
         n13938, n13939, n13940, n13941, n13942, n13943, n13944, n13945,
         n13946, n13947, n13948, n13949, n13950, n13951, n13952, n13953,
         n13954, n13955, n13956, n13957, n13958, n13959, n13960, n13961,
         n13962, n13963, n13964, n13965, n13966, n13967, n13968, n13969,
         n13970, n13971, n13972, n13973, n13974, n13975, n13976, n13977,
         n13978, n13979, n13980, n13981, n13982, n13983, n13984, n13985,
         n13986, n13987, n13988, n13989, n13990, n13991, n13992, n13993,
         n13994, n13995, n13996, n13997, n13998, n13999, n14000, n14001,
         n14002, n14003, n14004, n14005, n14006, n14007, n14008, n14009,
         n14010, n14011, n14012, n14013, n14014, n14015, n14016, n14017,
         n14018, n14019, n14020, n14021, n14022, n14023, n14024, n14025,
         n14026, n14027, n14028, n14029, n14030, n14031, n14032, n14033,
         n14034, n14035, n14036, n14037, n14038, n14039, n14040, n14041,
         n14042, n14043, n14044, n14045, n14046, n14047, n14048, n14049,
         n14050, n14051, n14052, n14053, n14054, n14055, n14056, n14057,
         n14058, n14059, n14060, n14061, n14062, n14063, n14064, n14065,
         n14066, n14067, n14068, n14069, n14070, n14071, n14072, n14073,
         n14074, n14075, n14076, n14077, n14078, n14079, n14080, n14081,
         n14082, n14083, n14084, n14085, n14086, n14087, n14088, n14089,
         n14090, n14091, n14092, n14093, n14094, n14095, n14096, n14097,
         n14098, n14099, n14100, n14101, n14102, n14103, n14104, n14105,
         n14106, n14107, n14108, n14109, n14110, n14111, n14112, n14113,
         n14114, n14115, n14116, n14117, n14118, n14119, n14120, n14121,
         n14122, n14123, n14124, n14125, n14126, n14127, n14128, n14129,
         n14130, n14131, n14132, n14133, n14134, n14135, n14136, n14137,
         n14138, n14139, n14140, n14141, n14142, n14143, n14144, n14145,
         n14146, n14147, n14148, n14149, n14150, n14151, n14152, n14153,
         n14154, n14155, n14156, n14157, n14158, n14159, n14160, n14161,
         n14162, n14163, n14164, n14165, n14166, n14167, n14168, n14169,
         n14170, n14171, n14172, n14173, n14174, n14175, n14176, n14177,
         n14178, n14179, n14180, n14181, n14182, n14183, n14184, n14185,
         n14186, n14187, n14188, n14189, n14190, n14191, n14192, n14193,
         n14194, n14195, n14196, n14197, n14198, n14199, n14200, n14201,
         n14202, n14203, n14204, n14205, n14206, n14207, n14208, n14209,
         n14210, n14211, n14212, n14213, n14214, n14215, n14216, n14217,
         n14218, n14219, n14220, n14221, n14222, n14223, n14224, n14225,
         n14226, n14227, n14228, n14229, n14230, n14231, n14232, n14233,
         n14234, n14235, n14236, n14237, n14238, n14239, n14240, n14241,
         n14242, n14243, n14244, n14245, n14246, n14247, n14248, n14249,
         n14250, n14251, n14252, n14253, n14254, n14255, n14256, n14257,
         n14258, n14259, n14260, n14261, n14262, n14263, n14264, n14265,
         n14266, n14267, n14268, n14269, n14270, n14271, n14272, n14273,
         n14274, n14275, n14276, n14277, n14278, n14279, n14280, n14281,
         n14282, n14283, n14284, n14285, n14286, n14287, n14288, n14289,
         n14290, n14291, n14292, n14293, n14294, n14295, n14296, n14297,
         n14298, n14299, n14300, n14301, n14302, n14303, n14304, n14305,
         n14306, n14307, n14308, n14309, n14310, n14311, n14312, n14313,
         n14314, n14315, n14316, n14317, n14318, n14319, n14320, n14321,
         n14322, n14323, n14324, n14325, n14326, n14327, n14328, n14329,
         n14330, n14331, n14332, n14333, n14334, n14335, n14336, n14337,
         n14338, n14339, n14340, n14341, n14342, n14343, n14344, n14345,
         n14346, n14347, n14348, n14349, n14350, n14351, n14352, n14353,
         n14354, n14355, n14356, n14357, n14358, n14359, n14360, n14361,
         n14362, n14363, n14364, n14365, n14366, n14367, n14368, n14369,
         n14370, n14371, n14372, n14373, n14374, n14375, n14376, n14377,
         n14378, n14379, n14380, n14381, n14382, n14383, n14384, n14385,
         n14386, n14387, n14388, n14389, n14390, n14391, n14392, n14393,
         n14394, n14395, n14396, n14397, n14398, n14399, n14400, n14401,
         n14402, n14403, n14404, n14405, n14406, n14407, n14408, n14409,
         n14410, n14411, n14412, n14413, n14414, n14415, n14416, n14417,
         n14418, n14419, n14420, n14421, n14422, n14423, n14424, n14425,
         n14426, n14427, n14428, n14429, n14430, n14431, n14432, n14433,
         n14434, n14435, n14436, n14437, n14438, n14439, n14440, n14441,
         n14442, n14443, n14444, n14445, n14446, n14447, n14448, n14449,
         n14450, n14451, n14452, n14453, n14454, n14455, n14456, n14457,
         n14458, n14459, n14460, n14461, n14462, n14463, n14464, n14465,
         n14466, n14467, n14468, n14469, n14470, n14471, n14472, n14473,
         n14474, n14475, n14476, n14477, n14478, n14479, n14480, n14481,
         n14482, n14483, n14484, n14485, n14486, n14487, n14488, n14489,
         n14490, n14491, n14492, n14493, n14494, n14495, n14496, n14497,
         n14498, n14499, n14500, n14501, n14502, n14503, n14504, n14505,
         n14506, n14507, n14508, n14509, n14510, n14511, n14512, n14513,
         n14514, n14515, n14516, n14517, n14518, n14519, n14520, n14521,
         n14522, n14523, n14524, n14525, n14526, n14527, n14528, n14529,
         n14530, n14531, n14532, n14533, n14534, n14535, n14536, n14537,
         n14538, n14539, n14540, n14541, n14542, n14543, n14544, n14545,
         n14546, n14547, n14548, n14549, n14550, n14551, n14552, n14553,
         n14554, n14555, n14556, n14557, n14558, n14559, n14560, n14561,
         n14562, n14563, n14564, n14565, n14566, n14567, n14568, n14569,
         n14570, n14571, n14572, n14573, n14574, n14575, n14576, n14577,
         n14578, n14579, n14580, n14581, n14582, n14583, n14584, n14585,
         n14586, n14587, n14588, n14589, n14590, n14591, n14592, n14593,
         n14594, n14595, n14596, n14597, n14598, n14599, n14600, n14601,
         n14602, n14603, n14604, n14605, n14606, n14607, n14608, n14609,
         n14610, n14611, n14612, n14613, n14614, n14615, n14616, n14617,
         n14618, n14619, n14620, n14621, n14622, n14623, n14624, n14625,
         n14626, n14627, n14628, n14629, n14630, n14631, n14632, n14633,
         n14634, n14635, n14636, n14637, n14638, n14639, n14640, n14641,
         n14642, n14643, n14644, n14645, n14646, n14647, n14648, n14649,
         n14650, n14651, n14652, n14653, n14654, n14655, n14656, n14657,
         n14658, n14659, n14660, n14661, n14662, n14663, n14664, n14665,
         n14666, n14667, n14668, n14669, n14670, n14671, n14672, n14673,
         n14674, n14675, n14676, n14677, n14678, n14679, n14680, n14681,
         n14682, n14683, n14684, n14685, n14686, n14687, n14688, n14689,
         n14690, n14691, n14692, n14693, n14694, n14695, n14696, n14697,
         n14698, n14699, n14700, n14701, n14702, n14703, n14704, n14705,
         n14706, n14707, n14708, n14709, n14710, n14711, n14712, n14713,
         n14714, n14715, n14716, n14717, n14718, n14719, n14720, n14721,
         n14722, n14723, n14724, n14725, n14726, n14727, n14728, n14729,
         n14730, n14731, n14732, n14733, n14734, n14735, n14736, n14737,
         n14738, n14739, n14740, n14741, n14742, n14743, n14744, n14745,
         n14746, n14747, n14748, n14749, n14750, n14751, n14752, n14753,
         n14754, n14755, n14756, n14757, n14758, n14759, n14760, n14761,
         n14762, n14763, n14764, n14765, n14766, n14767, n14768, n14769,
         n14770, n14771, n14772, n14773, n14774, n14775, n14776, n14777,
         n14778, n14779, n14780, n14781, n14782, n14783, n14784, n14785,
         n14786, n14787, n14788, n14789, n14790, n14791, n14792, n14793,
         n14794, n14795, n14796, n14797, n14798, n14799, n14800, n14801,
         n14802, n14803, n14804, n14805, n14806, n14807, n14808, n14809,
         n14810, n14811, n14812, n14813, n14814, n14815, n14816, n14817,
         n14818, n14819, n14820, n14821, n14822, n14823, n14824, n14825,
         n14826, n14827, n14828, n14829, n14830, n14831, n14832, n14833,
         n14834, n14835, n14836, n14837, n14838, n14839, n14840, n14841,
         n14842, n14843, n14844, n14845, n14846, n14847, n14848, n14849,
         n14850, n14851, n14852, n14853, n14854, n14855, n14856, n14857,
         n14858, n14859, n14860, n14861, n14862, n14863, n14864, n14865,
         n14866, n14867, n14868, n14869, n14870, n14871, n14872, n14873,
         n14874, n14875, n14876, n14877, n14878, n14879, n14880, n14881,
         n14882, n14883, n14884, n14885, n14886, n14887, n14888, n14889,
         n14890, n14891, n14892, n14893, n14894, n14895, n14896, n14897,
         n14898, n14899, n14900, n14901, n14902, n14903, n14904, n14905,
         n14906, n14907, n14908, n14909, n14910, n14911, n14912, n14913,
         n14914, n14915, n14916, n14917, n14918, n14919, n14920, n14921,
         n14922, n14923, n14924, n14925, n14926, n14927, n14928, n14929,
         n14930, n14931, n14932, n14933, n14934, n14935, n14936, n14937,
         n14938, n14939, n14940, n14941, n14942, n14943, n14944, n14945,
         n14946, n14947, n14948, n14949, n14950, n14951, n14952, n14953,
         n14954, n14955, n14956, n14957, n14958, n14959, n14960, n14961,
         n14962, n14963, n14964, n14965, n14966, n14967, n14968, n14969,
         n14970, n14971, n14972, n14973, n14974, n14975, n14976, n14977,
         n14978, n14979, n14980, n14981, n14982, n14983, n14984, n14985,
         n14986, n14987, n14988, n14989, n14990, n14991, n14992, n14993,
         n14994, n14995, n14996, n14997, n14998, n14999, n15000, n15001,
         n15002, n15003, n15004, n15005, n15006, n15007, n15008, n15009,
         n15010, n15011, n15012, n15013, n15014, n15015, n15016, n15017,
         n15018, n15019, n15020, n15021, n15022, n15023, n15024, n15025,
         n15026, n15027, n15028, n15029, n15030, n15031, n15032, n15033,
         n15034, n15035, n15036, n15037, n15038, n15039, n15040, n15041,
         n15042, n15043, n15044, n15045, n15046, n15047, n15048, n15049,
         n15050, n15051, n15052, n15053, n15054, n15055, n15056, n15057,
         n15058, n15059, n15060, n15061, n15062, n15063, n15064, n15065,
         n15066, n15067, n15068, n15069, n15070, n15071, n15072, n15073,
         n15074, n15075, n15076, n15077, n15078, n15079, n15080, n15081,
         n15082, n15083, n15084, n15085, n15086, n15087, n15088, n15089,
         n15090, n15091, n15092, n15093, n15094, n15095, n15096, n15097,
         n15098, n15099, n15100, n15101, n15102, n15103, n15104, n15105,
         n15106, n15107, n15108, n15109, n15110, n15111, n15112, n15113,
         n15114, n15115, n15116, n15117, n15118, n15119, n15120, n15121,
         n15122, n15123, n15124, n15125, n15126, n15127, n15128, n15129,
         n15130, n15131, n15132, n15133, n15134, n15135, n15136, n15137,
         n15138, n15139, n15140, n15141, n15142, n15143, n15144, n15145,
         n15146, n15147, n15148, n15149, n15150, n15151, n15152, n15153,
         n15154, n15155, n15156, n15157, n15158, n15159, n15160, n15161,
         n15162, n15163, n15164, n15165, n15166, n15167, n15168, n15169,
         n15170, n15171, n15172, n15173, n15174, n15175, n15176, n15177,
         n15178, n15179, n15180, n15181, n15182, n15183, n15184, n15185,
         n15186, n15187, n15188, n15189, n15190, n15191, n15192, n15193,
         n15194, n15195, n15196, n15197, n15198, n15199, n15200, n15201,
         n15202, n15203, n15204, n15205, n15206, n15207, n15208, n15209,
         n15210, n15211, n15212, n15213, n15214, n15215, n15216, n15217,
         n15218, n15219, n15220, n15221, n15222, n15223, n15224, n15225,
         n15226, n15227, n15228, n15229, n15230, n15231, n15232, n15233,
         n15234, n15235, n15236, n15237, n15238, n15239, n15240, n15241,
         n15242, n15243, n15244, n15245, n15246, n15247, n15248, n15249,
         n15250, n15251, n15252, n15253, n15254, n15255, n15256, n15257,
         n15258, n15259, n15260, n15261, n15262, n15263, n15264, n15265,
         n15266, n15267, n15268, n15269, n15270, n15271, n15272, n15273,
         n15274, n15275, n15276, n15277, n15278, n15279, n15280, n15281,
         n15282, n15283, n15284, n15285, n15286, n15287, n15288, n15289,
         n15290, n15291, n15292, n15293, n15294, n15295, n15296, n15297,
         n15298, n15299, n15300, n15301, n15302, n15303, n15304, n15305,
         n15306, n15307, n15308, n15309, n15310, n15311, n15312, n15313,
         n15314, n15315, n15316, n15317, n15318, n15319, n15320, n15321,
         n15322, n15323, n15324, n15325, n15326, n15327, n15328, n15329,
         n15330, n15331, n15332, n15333, n15334, n15335, n15336, n15337,
         n15338, n15339, n15340, n15341, n15342, n15343, n15344, n15345,
         n15346, n15347, n15348, n15349, n15350, n15351, n15352, n15353,
         n15354, n15355, n15356, n15357, n15358, n15359, n15360, n15361,
         n15362, n15363, n15364, n15365, n15366, n15367, n15368, n15369,
         n15370, n15371, n15372, n15373, n15374, n15375, n15376, n15377,
         n15378, n15379, n15380, n15381, n15382, n15383, n15384, n15385,
         n15386, n15387, n15388, n15389, n15390, n15391, n15392, n15393,
         n15394, n15395, n15396, n15397, n15398, n15399, n15400, n15401,
         n15402, n15403, n15404, n15405, n15406, n15407, n15408, n15409,
         n15410, n15411, n15412, n15413, n15414, n15415, n15416, n15417,
         n15418, n15419, n15420, n15421, n15422, n15423, n15424, n15425,
         n15426, n15427, n15428, n15429, n15430, n15431, n15432, n15433,
         n15434, n15435, n15436, n15437, n15438, n15439, n15440, n15441,
         n15442, n15443, n15444, n15445, n15446, n15447, n15448, n15449,
         n15450, n15451, n15452, n15453, n15454, n15455, n15456, n15457,
         n15458, n15459, n15460, n15461, n15462, n15463, n15464, n15465,
         n15466, n15467, n15468, n15469, n15470, n15471, n15472, n15473,
         n15474, n15475, n15476, n15477, n15478, n15479, n15480, n15481,
         n15482, n15483, n15484, n15485, n15486, n15487, n15488, n15489,
         n15490, n15491, n15492, n15493, n15494, n15495, n15496, n15497,
         n15498, n15499, n15500, n15501, n15502, n15503, n15504, n15505,
         n15506, n15507, n15508, n15509, n15510, n15511, n15512, n15513,
         n15514, n15515, n15516, n15517, n15518, n15519, n15520, n15521,
         n15522, n15523, n15524, n15525, n15526, n15527, n15528, n15529,
         n15530, n15531, n15532, n15533, n15534, n15535, n15536, n15537,
         n15538, n15539, n15540, n15541, n15542, n15543, n15544, n15545,
         n15546, n15547, n15548, n15549, n15550, n15551, n15552, n15553,
         n15554, n15555, n15556, n15557, n15558, n15559, n15560, n15561,
         n15562, n15563, n15564, n15565, n15566, n15567, n15568, n15569,
         n15570, n15571, n15572, n15573, n15574, n15575, n15576, n15577,
         n15578, n15579, n15580, n15581, n15582, n15583, n15584, n15585,
         n15586, n15587, n15588, n15589, n15590, n15591, n15592, n15593,
         n15594, n15595, n15596, n15597, n15598, n15599, n15600, n15601,
         n15602, n15603, n15604, n15605, n15606, n15607, n15608, n15609,
         n15610, n15611, n15612, n15613, n15614, n15615, n15616, n15617,
         n15618, n15619, n15620, n15621, n15622, n15623, n15624, n15625,
         n15626, n15627, n15628, n15629, n15630, n15631, n15632, n15633,
         n15634, n15635, n15636, n15637, n15638, n15639, n15640, n15641,
         n15642, n15643, n15644, n15645, n15646, n15647, n15648, n15649,
         n15650, n15651, n15652, n15653, n15654, n15655, n15656, n15657,
         n15658, n15659, n15660, n15661, n15662, n15663, n15664, n15665,
         n15666, n15667, n15668, n15669, n15670, n15671, n15672, n15673,
         n15674, n15675, n15676, n15677, n15678, n15679, n15680, n15681,
         n15682, n15683, n15684, n15685, n15686, n15687, n15688, n15689,
         n15690, n15691, n15692, n15693, n15694, n15695, n15696, n15697,
         n15698, n15699, n15700, n15701, n15702, n15703, n15704, n15705,
         n15706, n15707, n15708, n15709, n15710, n15711, n15712, n15713,
         n15714, n15715, n15716, n15717, n15718, n15719, n15720, n15721,
         n15722, n15723, n15724, n15725, n15726, n15727, n15728, n15729,
         n15730, n15731, n15732, n15733, n15734, n15735, n15736, n15737,
         n15738, n15739, n15740, n15741, n15742, n15743, n15744, n15745,
         n15746, n15747, n15748, n15749, n15750, n15751, n15752, n15753,
         n15754, n15755, n15756, n15757, n15758, n15759, n15760, n15761,
         n15762, n15763, n15764, n15765, n15766, n15767, n15768, n15769,
         n15770, n15771, n15772, n15773, n15774, n15775, n15776, n15777,
         n15778, n15779, n15780, n15781, n15782, n15783, n15784, n15785,
         n15786, n15787, n15788, n15789, n15790, n15791, n15792, n15793,
         n15794, n15795, n15796, n15797, n15798, n15799, n15800, n15801,
         n15802, n15803, n15804, n15805, n15806, n15807, n15808, n15809,
         n15810, n15811, n15812, n15813, n15814, n15815, n15816, n15817,
         n15818, n15819, n15820, n15821, n15822, n15823, n15824, n15825,
         n15826, n15827, n15828, n15829, n15830, n15831, n15832, n15833,
         n15834, n15835, n15836, n15837, n15838, n15839, n15840, n15841,
         n15842, n15843, n15844, n15845, n15846, n15847, n15848, n15849,
         n15850, n15851, n15852, n15853, n15854, n15855, n15856, n15857,
         n15858, n15859, n15860, n15861, n15862, n15863, n15864, n15865,
         n15866, n15867, n15868, n15869, n15870, n15871, n15872, n15873,
         n15874, n15875, n15876, n15877, n15878, n15879, n15880, n15881,
         n15882, n15883, n15884, n15885, n15886, n15887, n15888, n15889,
         n15890, n15891, n15892, n15893, n15894, n15895, n15896, n15897,
         n15898, n15899, n15900, n15901, n15902, n15903, n15904, n15905,
         n15906, n15907, n15908, n15909, n15910, n15911, n15912, n15913,
         n15914, n15915, n15916, n15917, n15918, n15919, n15920, n15921,
         n15922, n15923, n15924, n15925, n15926, n15927, n15928, n15929,
         n15930, n15931, n15932, n15933, n15934, n15935, n15936, n15937,
         n15938, n15939, n15940, n15941, n15942, n15943, n15944, n15945,
         n15946, n15947, n15948, n15949, n15950, n15951, n15952, n15953,
         n15954, n15955, n15956, n15957, n15958, n15959, n15960, n15961,
         n15962, n15963, n15964, n15965, n15966, n15967, n15968, n15969,
         n15970, n15971, n15972, n15973, n15974, n15975, n15976, n15977,
         n15978, n15979, n15980, n15981, n15982, n15983, n15984, n15985,
         n15986, n15987, n15988, n15989, n15990, n15991, n15992, n15993,
         n15994, n15995, n15996, n15997, n15998, n15999, n16000, n16001,
         n16002, n16003, n16004, n16005, n16006, n16007, n16008, n16009,
         n16010, n16011, n16012, n16013, n16014, n16015, n16016, n16017,
         n16018, n16019, n16020, n16021, n16022, n16023, n16024, n16025,
         n16026, n16027, n16028, n16029, n16030, n16031, n16032, n16033,
         n16034, n16035, n16036, n16037, n16038, n16039, n16040, n16041,
         n16042, n16043, n16044, n16045, n16046, n16047, n16048, n16049,
         n16050, n16051, n16052, n16053, n16054, n16055, n16056, n16057,
         n16058, n16059, n16060, n16061, n16062, n16063, n16064, n16065,
         n16066, n16067, n16068, n16069, n16070, n16071, n16072, n16073,
         n16074, n16075, n16076, n16077, n16078, n16079, n16080, n16081,
         n16082, n16083, n16084, n16085, n16086, n16087, n16088, n16089,
         n16090, n16091, n16092, n16093, n16094, n16095, n16096, n16097,
         n16098, n16099, n16100, n16101, n16102, n16103, n16104, n16105,
         n16106, n16107, n16108, n16109, n16110, n16111, n16112, n16113,
         n16114, n16115, n16116, n16117, n16118, n16119, n16120, n16121,
         n16122, n16123, n16124, n16125, n16126, n16127, n16128, n16129,
         n16130, n16131, n16132, n16133, n16134, n16135, n16136, n16137,
         n16138, n16139, n16140, n16141, n16142, n16143, n16144, n16145,
         n16146, n16147, n16148, n16149, n16150, n16151, n16152, n16153,
         n16154, n16155, n16156, n16157, n16158, n16159, n16160, n16161,
         n16162, n16163, n16164, n16165, n16166, n16167, n16168, n16169,
         n16170, n16171, n16172, n16173, n16174, n16175, n16176, n16177,
         n16178, n16179, n16180, n16181, n16182, n16183, n16184, n16185,
         n16186, n16187, n16188, n16189, n16190, n16191, n16192, n16193,
         n16194, n16195, n16196, n16197, n16198, n16199, n16200, n16201,
         n16202, n16203, n16204, n16205, n16206, n16207, n16208, n16209,
         n16210, n16211, n16212, n16213, n16214, n16215, n16216, n16217,
         n16218, n16219, n16220, n16221, n16222, n16223, n16224, n16225,
         n16226, n16227, n16228, n16229, n16230, n16231, n16232, n16233,
         n16234, n16235, n16236, n16237, n16238, n16239, n16240, n16241,
         n16242, n16243, n16244, n16245, n16246, n16247, n16248, n16249,
         n16250, n16251, n16252, n16253, n16254, n16255, n16256, n16257,
         n16258, n16259, n16260, n16261, n16262, n16263, n16264, n16265,
         n16266, n16267, n16268, n16269, n16270, n16271, n16272, n16273,
         n16274, n16275, n16276, n16277, n16278, n16279, n16280, n16281,
         n16282, n16283, n16284, n16285, n16286, n16287, n16288, n16289,
         n16290, n16291, n16292, n16293, n16294, n16295, n16296, n16297,
         n16298, n16299, n16300, n16301, n16302, n16303, n16304, n16305,
         n16306, n16307, n16308, n16309, n16310, n16311, n16312, n16313,
         n16314, n16315, n16316, n16317, n16318, n16319, n16320, n16321,
         n16322, n16323, n16324, n16325, n16326, n16327, n16328, n16329,
         n16330, n16331, n16332, n16333, n16334, n16335, n16336, n16337,
         n16338, n16339, n16340, n16341, n16342, n16343, n16344, n16345,
         n16346, n16347, n16348, n16349, n16350, n16351, n16352, n16353,
         n16354, n16355, n16356, n16357, n16358, n16359, n16360, n16361,
         n16362, n16363, n16364, n16365, n16366, n16367, n16368, n16369,
         n16370, n16371, n16372, n16373, n16374, n16375, n16376, n16377,
         n16378, n16379, n16380, n16381, n16382, n16383, n16384, n16385,
         n16386, n16387, n16388, n16389, n16390, n16391, n16392, n16393,
         n16394, n16395, n16396, n16397, n16398, n16399, n16400, n16401,
         n16402, n16403, n16404, n16405, n16406, n16407, n16408, n16409,
         n16410, n16411, n16412, n16413, n16414, n16415, n16416, n16417,
         n16418, n16419, n16420, n16421, n16422, n16423, n16424, n16425,
         n16426, n16427, n16428, n16429, n16430, n16431, n16432, n16433,
         n16434, n16435, n16436, n16437, n16438, n16439, n16440, n16441,
         n16442, n16443, n16444, n16445, n16446, n16447, n16448, n16449,
         n16450, n16451, n16452, n16453, n16454, n16455, n16456, n16457,
         n16458, n16459, n16460, n16461, n16462, n16463, n16464, n16465,
         n16466, n16467, n16468, n16469, n16470, n16471, n16472, n16473,
         n16474, n16475, n16476, n16477, n16478, n16479, n16480, n16481,
         n16482, n16483, n16484, n16485, n16486, n16487, n16488, n16489,
         n16490, n16491, n16492, n16493, n16494, n16495, n16496, n16497,
         n16498, n16499, n16500, n16501, n16502, n16503, n16504, n16505,
         n16506, n16507, n16508, n16509, n16510, n16511, n16512, n16513,
         n16514, n16515, n16516, n16517, n16518, n16519, n16520, n16521,
         n16522, n16523, n16524, n16525, n16526, n16527, n16528, n16529,
         n16530, n16531, n16532, n16533, n16534, n16535, n16536, n16537,
         n16538, n16539, n16540, n16541, n16542, n16543, n16544, n16545,
         n16546, n16547, n16548, n16549, n16550, n16551, n16552, n16553,
         n16554, n16555, n16556, n16557, n16558, n16559, n16560, n16561,
         n16562, n16563, n16564, n16565, n16566, n16567, n16568, n16569,
         n16570, n16571, n16572, n16573, n16574, n16575, n16576, n16577,
         n16578, n16579, n16580, n16581, n16582, n16583, n16584, n16585,
         n16586, n16587, n16588, n16589, n16590, n16591, n16592, n16593,
         n16594, n16595, n16596, n16597, n16598, n16599, n16600, n16601,
         n16602, n16603, n16604, n16605, n16606, n16607, n16608, n16609,
         n16610, n16611, n16612, n16613, n16614, n16615, n16616, n16617,
         n16618, n16619, n16620, n16621, n16622, n16623, n16624, n16625,
         n16626, n16627, n16628, n16629, n16630, n16631, n16632, n16633,
         n16634, n16635, n16636, n16637, n16638, n16639, n16640, n16641,
         n16642, n16643, n16644, n16645, n16646, n16647, n16648, n16649,
         n16650, n16651, n16652, n16653, n16654, n16655, n16656, n16657,
         n16658, n16659, n16660, n16661, n16662, n16663, n16664, n16665,
         n16666, n16667, n16668, n16669, n16670, n16671, n16672, n16673,
         n16674, n16675, n16676, n16677, n16678, n16679, n16680, n16681,
         n16682, n16683, n16684, n16685, n16686, n16687, n16688, n16689,
         n16690, n16691, n16692, n16693, n16694, n16695, n16696, n16697,
         n16698, n16699, n16700, n16701, n16702, n16703, n16704, n16705,
         n16706, n16707, n16708, n16709, n16710, n16711, n16712, n16713,
         n16714, n16715, n16716, n16717, n16718, n16719, n16720, n16721,
         n16722, n16723, n16724, n16725, n16726, n16727, n16728, n16729,
         n16730, n16731, n16732, n16733, n16734, n16735, n16736, n16737,
         n16738, n16739, n16740, n16741, n16742, n16743, n16744, n16745,
         n16746, n16747, n16748, n16749, n16750, n16751, n16752, n16753,
         n16754, n16755, n16756, n16757, n16758, n16759, n16760, n16761,
         n16762, n16763, n16764, n16765, n16766, n16767, n16768, n16769,
         n16770, n16771, n16772, n16773, n16774, n16775, n16776, n16777,
         n16778, n16779, n16780, n16781, n16782, n16783, n16784, n16785,
         n16786, n16787, n16788, n16789, n16790, n16791, n16792, n16793,
         n16794, n16795, n16796, n16797, n16798, n16799, n16800, n16801,
         n16802, n16803, n16804, n16805, n16806, n16807, n16808, n16809,
         n16810, n16811, n16812, n16813, n16814, n16815, n16816, n16817,
         n16818, n16819, n16820, n16821, n16822, n16823, n16824, n16825,
         n16826, n16827, n16828, n16829, n16830, n16831, n16832, n16833,
         n16834, n16835, n16836, n16837, n16838, n16839, n16840, n16841,
         n16842, n16843, n16844, n16845, n16846, n16847, n16848, n16849,
         n16850, n16851, n16852, n16853, n16854, n16855, n16856, n16857,
         n16858, n16859, n16860, n16861, n16862, n16863, n16864, n16865,
         n16866, n16867, n16868, n16869, n16870, n16871, n16872, n16873,
         n16874, n16875, n16876, n16877, n16878, n16879, n16880, n16881,
         n16882, n16883, n16884, n16885, n16886, n16887, n16888, n16889,
         n16890, n16891, n16892, n16893, n16894, n16895, n16896, n16897,
         n16898, n16899, n16900, n16901, n16902, n16903, n16904, n16905,
         n16906, n16907, n16908, n16909, n16910, n16911, n16912, n16913,
         n16914, n16915, n16916, n16917, n16918, n16919, n16920, n16921,
         n16922, n16923, n16924, n16925, n16926, n16927, n16928, n16929,
         n16930, n16931, n16932, n16933, n16934, n16935, n16936, n16937,
         n16938, n16939, n16940, n16941, n16942, n16943, n16944, n16945,
         n16946, n16947, n16948, n16949, n16950, n16951, n16952, n16953,
         n16954, n16955, n16956, n16957, n16958, n16959, n16960, n16961,
         n16962, n16963, n16964, n16965, n16966, n16967, n16968, n16969,
         n16970, n16971, n16972, n16973, n16974, n16975, n16976, n16977,
         n16978, n16979, n16980, n16981, n16982, n16983, n16984, n16985,
         n16986, n16987, n16988, n16989, n16990, n16991, n16992, n16993,
         n16994, n16995, n16996, n16997, n16998, n16999, n17000, n17001,
         n17002, n17003, n17004, n17005, n17006, n17007, n17008, n17009,
         n17010, n17011, n17012, n17013, n17014, n17015, n17016, n17017,
         n17018, n17019, n17020, n17021, n17022, n17023, n17024, n17025,
         n17026, n17027, n17028, n17029, n17030, n17031, n17032, n17033,
         n17034, n17035, n17036, n17037, n17038, n17039, n17040, n17041,
         n17042, n17043, n17044, n17045, n17046, n17047, n17048, n17049,
         n17050, n17051, n17052, n17053, n17054, n17055, n17056, n17057,
         n17058, n17059, n17060, n17061, n17062, n17063, n17064, n17065,
         n17066, n17067, n17068, n17069, n17070, n17071, n17072, n17073,
         n17074, n17075, n17076, n17077, n17078, n17079, n17080, n17081,
         n17082, n17083, n17084, n17085, n17086, n17087, n17088, n17089,
         n17090, n17091, n17092, n17093, n17094, n17095, n17096, n17097,
         n17098, n17099, n17100, n17101, n17102, n17103, n17104, n17105,
         n17106, n17107, n17108, n17109, n17110, n17111, n17112, n17113,
         n17114, n17115, n17116, n17117, n17118, n17119, n17120, n17121,
         n17122, n17123, n17124, n17125, n17126, n17127, n17128, n17129,
         n17130, n17131, n17132, n17133, n17134, n17135, n17136, n17137,
         n17138, n17139, n17140, n17141, n17142, n17143, n17144, n17145,
         n17146, n17147, n17148, n17149, n17150, n17151, n17152, n17153,
         n17154, n17155, n17156, n17157, n17158, n17159, n17160, n17161,
         n17162, n17163, n17164, n17165, n17166, n17167, n17168, n17169,
         n17170, n17171, n17172, n17173, n17174, n17175, n17176, n17177,
         n17178, n17179, n17180, n17181, n17182, n17183, n17184, n17185,
         n17186, n17187, n17188, n17189, n17190, n17191, n17192, n17193,
         n17194, n17195, n17196, n17197, n17198, n17199, n17200, n17201,
         n17202, n17203, n17204, n17205, n17206, n17207, n17208, n17209,
         n17210, n17211, n17212, n17213, n17214, n17215, n17216, n17217,
         n17218, n17219, n17220, n17221, n17222, n17223, n17224, n17225,
         n17226, n17227, n17228, n17229, n17230, n17231, n17232, n17233,
         n17234, n17235, n17236, n17237, n17238, n17239, n17240, n17241,
         n17242, n17243, n17244, n17245, n17246, n17247, n17248, n17249,
         n17250, n17251, n17252, n17253, n17254, n17255, n17256, n17257,
         n17258, n17259, n17260, n17261, n17262, n17263, n17264, n17265,
         n17266, n17267, n17268, n17269, n17270, n17271, n17272, n17273,
         n17274, n17275, n17276, n17277, n17278, n17279, n17280, n17281,
         n17282, n17283, n17284, n17285, n17286, n17287, n17288, n17289,
         n17290, n17291, n17292, n17293, n17294, n17295, n17296, n17297,
         n17298, n17299, n17300, n17301, n17302, n17303, n17304, n17305,
         n17306, n17307, n17308, n17309, n17310, n17311, n17312, n17313,
         n17314, n17315, n17316, n17317, n17318, n17319, n17320, n17321,
         n17322, n17323, n17324, n17325, n17326, n17327, n17328, n17329,
         n17330, n17331, n17332, n17333, n17334, n17335, n17336, n17337,
         n17338, n17339, n17340, n17341, n17342, n17343, n17344, n17345,
         n17346, n17347, n17348, n17349, n17350, n17351, n17352, n17353,
         n17354, n17355, n17356, n17357, n17358, n17359, n17360, n17361,
         n17362, n17363, n17364, n17365, n17366, n17367, n17368, n17369,
         n17370, n17371, n17372, n17373, n17374, n17375, n17376, n17377,
         n17378, n17379, n17380, n17381, n17382, n17383, n17384, n17385,
         n17386, n17387, n17388, n17389, n17390, n17391, n17392, n17393,
         n17394, n17395, n17396, n17397, n17398, n17399, n17400, n17401,
         n17402, n17403, n17404, n17405, n17406, n17407, n17408, n17409,
         n17410, n17411, n17412, n17413, n17414, n17415, n17416, n17417,
         n17418, n17419, n17420, n17421, n17422, n17423, n17424, n17425,
         n17426, n17427, n17428, n17429, n17430, n17431, n17432, n17433,
         n17434, n17435, n17436, n17437, n17438, n17439, n17440, n17441,
         n17442, n17443, n17444, n17445, n17446, n17447, n17448, n17449,
         n17450, n17451, n17452, n17453, n17454, n17455, n17456, n17457,
         n17458, n17459, n17460, n17461, n17462, n17463, n17464, n17465,
         n17466, n17467, n17468, n17469, n17470, n17471, n17472, n17473,
         n17474, n17475, n17476, n17477, n17478, n17479, n17480, n17481,
         n17482, n17483, n17484, n17485, n17486, n17487, n17488, n17489,
         n17490, n17491, n17492, n17493, n17494, n17495, n17496, n17497,
         n17498, n17499, n17500, n17501, n17502, n17503, n17504, n17505,
         n17506, n17507, n17508, n17509, n17510, n17511, n17512, n17513,
         n17514, n17515, n17516, n17517, n17518, n17519, n17520, n17521,
         n17522, n17523, n17524, n17525, n17526, n17527, n17528, n17529,
         n17530, n17531, n17532, n17533, n17534, n17535, n17536, n17537,
         n17538, n17539, n17540, n17541, n17542, n17543, n17544, n17545,
         n17546, n17547, n17548, n17549, n17550, n17551, n17552, n17553,
         n17554, n17555, n17556, n17557, n17558, n17559, n17560, n17561,
         n17562, n17563, n17564, n17565, n17566, n17567, n17568, n17569,
         n17570, n17571, n17572, n17573, n17574, n17575, n17576, n17577,
         n17578, n17579, n17580, n17581, n17582, n17583, n17584, n17585,
         n17586, n17587, n17588, n17589, n17590, n17591, n17592, n17593,
         n17594, n17595, n17596, n17597, n17598, n17599, n17600, n17601,
         n17602, n17603, n17604, n17605, n17606, n17607, n17608, n17609,
         n17610, n17611, n17612, n17613, n17614, n17615, n17616, n17617,
         n17618, n17619, n17620, n17621, n17622, n17623, n17624, n17625,
         n17626, n17627, n17628, n17629, n17630, n17631, n17632, n17633,
         n17634, n17635, n17636, n17637, n17638, n17639, n17640, n17641,
         n17642, n17643, n17644, n17645, n17646, n17647, n17648, n17649,
         n17650, n17651, n17652, n17653, n17654, n17655, n17656, n17657,
         n17658, n17659, n17660, n17661, n17662, n17663, n17664, n17665,
         n17666, n17667, n17668, n17669, n17670, n17671, n17672, n17673,
         n17674, n17675, n17676, n17677, n17678, n17679, n17680, n17681,
         n17682, n17683, n17684, n17685, n17686, n17687, n17688, n17689,
         n17690, n17691, n17692, n17693, n17694, n17695, n17696, n17697,
         n17698, n17699, n17700, n17701, n17702, n17703, n17704, n17705,
         n17706, n17707, n17708, n17709, n17710, n17711, n17712, n17713,
         n17714, n17715, n17716, n17717, n17718, n17719, n17720, n17721,
         n17722, n17723, n17724, n17725, n17726, n17727, n17728, n17729,
         n17730, n17731, n17732, n17733, n17734, n17735, n17736, n17737,
         n17738, n17739, n17740, n17741, n17742, n17743, n17744, n17745,
         n17746, n17747, n17748, n17749, n17750, n17751, n17752, n17753,
         n17754, n17755, n17756, n17757, n17758, n17759, n17760, n17761,
         n17762, n17763, n17764, n17765, n17766, n17767, n17768, n17769,
         n17770, n17771, n17772, n17773, n17774, n17775, n17776, n17777,
         n17778, n17779, n17780, n17781, n17782, n17783, n17784, n17785,
         n17786, n17787, n17788, n17789, n17790, n17791, n17792, n17793,
         n17794, n17795, n17796, n17797, n17798, n17799, n17800, n17801,
         n17802, n17803, n17804, n17805, n17806, n17807, n17808, n17809,
         n17810, n17811, n17812, n17813, n17814, n17815, n17816, n17817,
         n17818, n17819, n17820, n17821, n17822, n17823, n17824, n17825,
         n17826, n17827, n17828, n17829, n17830, n17831, n17832, n17833,
         n17834, n17835, n17836, n17837, n17838, n17839, n17840, n17841,
         n17842, n17843, n17844, n17845, n17846, n17847, n17848, n17849,
         n17850, n17851, n17852, n17853, n17854, n17855, n17856, n17857,
         n17858, n17859, n17860, n17861, n17862, n17863, n17864, n17865,
         n17866, n17867, n17868, n17869, n17870, n17871, n17872, n17873,
         n17874, n17875, n17876, n17877, n17878, n17879, n17880, n17881,
         n17882, n17883, n17884, n17885, n17886, n17887, n17888, n17889,
         n17890, n17891, n17892, n17893, n17894, n17895, n17896, n17897,
         n17898, n17899, n17900, n17901, n17902, n17903, n17904, n17905,
         n17906, n17907, n17908, n17909, n17910, n17911, n17912, n17913,
         n17914, n17915, n17916, n17917, n17918, n17919, n17920, n17921,
         n17922, n17923, n17924, n17925, n17926, n17927, n17928, n17929,
         n17930, n17931, n17932, n17933, n17934, n17935, n17936, n17937,
         n17938, n17939, n17940, n17941, n17942, n17943, n17944, n17945,
         n17946, n17947, n17948, n17949, n17950, n17951, n17952, n17953,
         n17954, n17955, n17956, n17957, n17958, n17959, n17960, n17961,
         n17962, n17963, n17964, n17965, n17966, n17967, n17968, n17969,
         n17970, n17971, n17972, n17973, n17974, n17975, n17976, n17977,
         n17978, n17979, n17980, n17981, n17982, n17983, n17984, n17985,
         n17986, n17987, n17988, n17989, n17990, n17991, n17992, n17993,
         n17994, n17995, n17996, n17997, n17998, n17999, n18000, n18001,
         n18002, n18003, n18004, n18005, n18006, n18007, n18008, n18009,
         n18010, n18011, n18012, n18013, n18014, n18015, n18016, n18017,
         n18018, n18019, n18020, n18021, n18022, n18023, n18024, n18025,
         n18026, n18027, n18028, n18029, n18030, n18031, n18032, n18033,
         n18034, n18035, n18036, n18037, n18038, n18039, n18040, n18041,
         n18042, n18043, n18044, n18045, n18046, n18047, n18048, n18049,
         n18050, n18051, n18052, n18053, n18054, n18055, n18056, n18057,
         n18058, n18059, n18060, n18061, n18062, n18063, n18064, n18065,
         n18066, n18067, n18068, n18069, n18070, n18071, n18072, n18073,
         n18074, n18075, n18076, n18077, n18078, n18079, n18080, n18081,
         n18082, n18083, n18084, n18085, n18086, n18087, n18088, n18089,
         n18090, n18091, n18092, n18093, n18094, n18095, n18096, n18097,
         n18098, n18099, n18100, n18101, n18102, n18103, n18104, n18105,
         n18106, n18107, n18108, n18109, n18110, n18111, n18112, n18113,
         n18114, n18115, n18116, n18117, n18118, n18119, n18120, n18121,
         n18122, n18123, n18124, n18125, n18126, n18127, n18128, n18129,
         n18130, n18131, n18132, n18133, n18134, n18135, n18136, n18137,
         n18138, n18139, n18140, n18141, n18142, n18143, n18144, n18145,
         n18146, n18147, n18148, n18149, n18150, n18151, n18152, n18153,
         n18154, n18155, n18156, n18157, n18158, n18159, n18160, n18161,
         n18162, n18163, n18164, n18165, n18166, n18167, n18168, n18169,
         n18170, n18171, n18172, n18173, n18174, n18175, n18176, n18177,
         n18178, n18179, n18180, n18181, n18182, n18183, n18184, n18185,
         n18186, n18187, n18188, n18189, n18190, n18191, n18192, n18193,
         n18194, n18195, n18196, n18197, n18198, n18199, n18200, n18201,
         n18202, n18203, n18204, n18205, n18206, n18207, n18208, n18209,
         n18210, n18211, n18212, n18213, n18214, n18215, n18216, n18217,
         n18218, n18219, n18220, n18221, n18222, n18223, n18224, n18225,
         n18226, n18227, n18228, n18229, n18230, n18231, n18232, n18233,
         n18234, n18235, n18236, n18237, n18238, n18239, n18240, n18241,
         n18242, n18243, n18244, n18245, n18246, n18247, n18248, n18249,
         n18250, n18251, n18252, n18253, n18254, n18255, n18256, n18257,
         n18258, n18259, n18260, n18261, n18262, n18263, n18264, n18265,
         n18266, n18267, n18268, n18269, n18270, n18271, n18272, n18273,
         n18274, n18275, n18276, n18277, n18278, n18279, n18280, n18281,
         n18282, n18283, n18284, n18285, n18286, n18287, n18288, n18289,
         n18290, n18291, n18292, n18293, n18294, n18295, n18296, n18297,
         n18298, n18299, n18300, n18301, n18302, n18303, n18304, n18305,
         n18306, n18307, n18308, n18309, n18310, n18311, n18312, n18313,
         n18314, n18315, n18316, n18317, n18318, n18319, n18320, n18321,
         n18322, n18323, n18324, n18325, n18326, n18327, n18328, n18329,
         n18330, n18331, n18332, n18333, n18334, n18335, n18336, n18337,
         n18338, n18339, n18340, n18341, n18342, n18343, n18344, n18345,
         n18346, n18347, n18348, n18349, n18350, n18351, n18352, n18353,
         n18354, n18355, n18356, n18357, n18358, n18359, n18360, n18361,
         n18362, n18363, n18364, n18365, n18366, n18367, n18368, n18369,
         n18370, n18371, n18372, n18373, n18374, n18375, n18376, n18377,
         n18378, n18379, n18380, n18381, n18382, n18383, n18384, n18385,
         n18386, n18387, n18388, n18389, n18390, n18391, n18392, n18393,
         n18394, n18395, n18396, n18397, n18398, n18399, n18400, n18401,
         n18402, n18403, n18404, n18405, n18406, n18407, n18408, n18409,
         n18410, n18411, n18412, n18413, n18414, n18415, n18416, n18417,
         n18418, n18419, n18420, n18421, n18422, n18423, n18424, n18425,
         n18426, n18427, n18428, n18429, n18430, n18431, n18432, n18433,
         n18434, n18435, n18436, n18437, n18438, n18439, n18440, n18441,
         n18442, n18443, n18444, n18445, n18446, n18447, n18448, n18449,
         n18450, n18451, n18452, n18453, n18454, n18455, n18456, n18457,
         n18458, n18459, n18460, n18461, n18462, n18463, n18464, n18465,
         n18466, n18467, n18468, n18469, n18470, n18471, n18472, n18473,
         n18474, n18475, n18476, n18477, n18478, n18479, n18480, n18481,
         n18482, n18483, n18484, n18485, n18486, n18487, n18488, n18489,
         n18490, n18491, n18492, n18493, n18494, n18495, n18496, n18497,
         n18498, n18499, n18500, n18501, n18502, n18503, n18504, n18505,
         n18506, n18507, n18508, n18509, n18510, n18511, n18512, n18513,
         n18514, n18515, n18516, n18517, n18518, n18519, n18520, n18521,
         n18522, n18523, n18524, n18525, n18526, n18527, n18528, n18529,
         n18530, n18531, n18532, n18533, n18534, n18535, n18536, n18537,
         n18538, n18539, n18540, n18541, n18542, n18543, n18544, n18545,
         n18546, n18547, n18548, n18549, n18550, n18551, n18552, n18553,
         n18554, n18555, n18556, n18557, n18558, n18559, n18560, n18561,
         n18562, n18563, n18564, n18565, n18566, n18567, n18568, n18569,
         n18570, n18571, n18572, n18573, n18574, n18575, n18576, n18577,
         n18578, n18579, n18580, n18581, n18582, n18583, n18584, n18585,
         n18586, n18587, n18588, n18589, n18590, n18591, n18592, n18593,
         n18594, n18595, n18596, n18597, n18598, n18599, n18600, n18601,
         n18602, n18603, n18604, n18605, n18606, n18607, n18608, n18609,
         n18610, n18611, n18612, n18613, n18614, n18615, n18616, n18617,
         n18618, n18619, n18620, n18621, n18622, n18623, n18624, n18625,
         n18626, n18627, n18628, n18629, n18630, n18631, n18632, n18633,
         n18634, n18635, n18636, n18637, n18638, n18639, n18640, n18641,
         n18642, n18643, n18644, n18645, n18646, n18647, n18648, n18649,
         n18650, n18651, n18652, n18653, n18654, n18655, n18656, n18657,
         n18658, n18659, n18660, n18661, n18662, n18663, n18664, n18665,
         n18666, n18667, n18668, n18669, n18670, n18671, n18672, n18673,
         n18674, n18675, n18676, n18677, n18678, n18679, n18680, n18681,
         n18682, n18683, n18684, n18685, n18686, n18687, n18688, n18689,
         n18690, n18691, n18692, n18693, n18694, n18695, n18696, n18697,
         n18698, n18699, n18700, n18701, n18702, n18703, n18704, n18705,
         n18706, n18707, n18708, n18709, n18710, n18711, n18712, n18713,
         n18714, n18715, n18716, n18717, n18718, n18719, n18720, n18721,
         n18722, n18723, n18724, n18725, n18726, n18727, n18728, n18729,
         n18730, n18731, n18732, n18733, n18734, n18735, n18736, n18737,
         n18738, n18739, n18740, n18741, n18742, n18743, n18744, n18745,
         n18746, n18747, n18748, n18749, n18750, n18751, n18752, n18753,
         n18754, n18755, n18756, n18757, n18758, n18759, n18760, n18761,
         n18762, n18763, n18764, n18765, n18766, n18767, n18768, n18769,
         n18770, n18771, n18772, n18773, n18774, n18775, n18776, n18777,
         n18778, n18779, n18780, n18781, n18782, n18783, n18784, n18785,
         n18786, n18787, n18788, n18789, n18790, n18791, n18792, n18793,
         n18794, n18795, n18796, n18797, n18798, n18799, n18800, n18801,
         n18802, n18803, n18804, n18805, n18806, n18807, n18808, n18809,
         n18810, n18811, n18812, n18813, n18814, n18815, n18816, n18817,
         n18818, n18819, n18820, n18821, n18822, n18823, n18824, n18825,
         n18826, n18827, n18828, n18829, n18830, n18831, n18832, n18833,
         n18834, n18835, n18836, n18837, n18838, n18839, n18840, n18841,
         n18842, n18843, n18844, n18845, n18846, n18847, n18848, n18849,
         n18850, n18851, n18852, n18853, n18854, n18855, n18856, n18857,
         n18858, n18859, n18860, n18861, n18862, n18863, n18864, n18865,
         n18866, n18867, n18868, n18869, n18870, n18871, n18872, n18873,
         n18874, n18875, n18876, n18877, n18878, n18879, n18880, n18881,
         n18882, n18883, n18884, n18885, n18886, n18887, n18888, n18889,
         n18890, n18891, n18892, n18893, n18894, n18895, n18896, n18897,
         n18898, n18899, n18900, n18901, n18902, n18903, n18904, n18905,
         n18906, n18907, n18908, n18909, n18910, n18911, n18912, n18913,
         n18914, n18915, n18916, n18917, n18918, n18919, n18920, n18921,
         n18922, n18923, n18924, n18925, n18926, n18927, n18928, n18929,
         n18930, n18931, n18932, n18933, n18934, n18935, n18936, n18937,
         n18938, n18939, n18940, n18941, n18942, n18943, n18944, n18945,
         n18946, n18947, n18948, n18949, n18950, n18951, n18952, n18953,
         n18954, n18955, n18956, n18957, n18958, n18959, n18960, n18961,
         n18962, n18963, n18964, n18965, n18966, n18967, n18968, n18969,
         n18970, n18971, n18972, n18973, n18974, n18975, n18976, n18977,
         n18978, n18979, n18980, n18981, n18982, n18983, n18984, n18985,
         n18986, n18987, n18988, n18989, n18990, n18991, n18992, n18993,
         n18994, n18995, n18996, n18997, n18998, n18999, n19000, n19001,
         n19002, n19003, n19004, n19005, n19006, n19007, n19008, n19009,
         n19010, n19011, n19012, n19013, n19014, n19015, n19016, n19017,
         n19018, n19019, n19020, n19021, n19022, n19023, n19024, n19025,
         n19026, n19027, n19028, n19029, n19030, n19031, n19032, n19033,
         n19034, n19035, n19036, n19037, n19038, n19039, n19040, n19041,
         n19042, n19043, n19044, n19045, n19046, n19047, n19048, n19049,
         n19050, n19051, n19052, n19053, n19054, n19055, n19056, n19057,
         n19058, n19059, n19060, n19061, n19062, n19063, n19064, n19065,
         n19066, n19067, n19068, n19069, n19070, n19071, n19072, n19073,
         n19074, n19075, n19076, n19077, n19078, n19079, n19080, n19081,
         n19082, n19083, n19084, n19085, n19086, n19087, n19088, n19089,
         n19090, n19091, n19092, n19093, n19094, n19095, n19096, n19097,
         n19098, n19099, n19100, n19101, n19102, n19103, n19104, n19105,
         n19106, n19107, n19108, n19109, n19110, n19111, n19112, n19113,
         n19114, n19115, n19116, n19117, n19118, n19119, n19120, n19121,
         n19122, n19123, n19124, n19125, n19126, n19127, n19128, n19129,
         n19130, n19131, n19132, n19133, n19134, n19135, n19136, n19137,
         n19138, n19139, n19140, n19141, n19142, n19143, n19144, n19145,
         n19146, n19147, n19148, n19149, n19150, n19151, n19152, n19153,
         n19154, n19155, n19156, n19157, n19158, n19159, n19160, n19161,
         n19162, n19163, n19164, n19165, n19166, n19167, n19168, n19169,
         n19170, n19171, n19172, n19173, n19174, n19175, n19176, n19177,
         n19178, n19179, n19180, n19181, n19182, n19183, n19184, n19185,
         n19186, n19187, n19188, n19189, n19190, n19191, n19192, n19193,
         n19194, n19195, n19196, n19197, n19198, n19199, n19200, n19201,
         n19202, n19203, n19204, n19205, n19206, n19207, n19208, n19209,
         n19210, n19211, n19212, n19213, n19214, n19215, n19216, n19217,
         n19218, n19219, n19220, n19221, n19222, n19223, n19224, n19225,
         n19226, n19227, n19228, n19229, n19230, n19231, n19232, n19233,
         n19234, n19235, n19236, n19237, n19238, n19239, n19240, n19241,
         n19242, n19243, n19244, n19245, n19246, n19247, n19248, n19249,
         n19250, n19251, n19252, n19253, n19254, n19255, n19256, n19257,
         n19258, n19259, n19260, n19261, n19262, n19263, n19264, n19265,
         n19266, n19267, n19268, n19269, n19270, n19271, n19272, n19273,
         n19274, n19275, n19276, n19277, n19278, n19279, n19280, n19281,
         n19282, n19283, n19284, n19285, n19286, n19287, n19288, n19289,
         n19290, n19291, n19292, n19293, n19294, n19295, n19296, n19297,
         n19298, n19299, n19300, n19301, n19302, n19303, n19304, n19305,
         n19306, n19307, n19308, n19309, n19310, n19311, n19312, n19313,
         n19314, n19315, n19316, n19317, n19318, n19319, n19320, n19321,
         n19322, n19323, n19324, n19325, n19326, n19327, n19328, n19329,
         n19330, n19331, n19332, n19333, n19334, n19335, n19336, n19337,
         n19338, n19339, n19340, n19341, n19342, n19343, n19344, n19345,
         n19346, n19347, n19348, n19349, n19350, n19351, n19352, n19353,
         n19354, n19355, n19356, n19357, n19358, n19359, n19360, n19361,
         n19362, n19363, n19364, n19365, n19366, n19367, n19368, n19369,
         n19370, n19371, n19372, n19373, n19374, n19375, n19376, n19377,
         n19378, n19379, n19380, n19381, n19382, n19383, n19384, n19385,
         n19386, n19387, n19388, n19389, n19390, n19391, n19392, n19393,
         n19394, n19395, n19396, n19397, n19398, n19399, n19400, n19401,
         n19402, n19403, n19404, n19405, n19406, n19407, n19408, n19409,
         n19410, n19411, n19412, n19413, n19414, n19415, n19416, n19417,
         n19418, n19419, n19420, n19421, n19422, n19423, n19424, n19425,
         n19426, n19427, n19428, n19429, n19430, n19431, n19432, n19433,
         n19434, n19435, n19436, n19437, n19438, n19439, n19440, n19441,
         n19442, n19443, n19444, n19445, n19446, n19447, n19448, n19449,
         n19450, n19451, n19452, n19453, n19454, n19455, n19456, n19457,
         n19458, n19459, n19460, n19461, n19462, n19463, n19464, n19465,
         n19466, n19467, n19468, n19469, n19470, n19471, n19472, n19473,
         n19474, n19475, n19476, n19477, n19478, n19479, n19480, n19481,
         n19482, n19483, n19484, n19485, n19486, n19487, n19488, n19489,
         n19490, n19491, n19492, n19493, n19494, n19495, n19496, n19497,
         n19498, n19499, n19500, n19501, n19502, n19503, n19504, n19505,
         n19506, n19507, n19508, n19509, n19510, n19511, n19512, n19513,
         n19514, n19515, n19516, n19517, n19518, n19519, n19520, n19521,
         n19522, n19523, n19524, n19525, n19526, n19527, n19528, n19529,
         n19530, n19531, n19532, n19533, n19534, n19535, n19536, n19537,
         n19538, n19539, n19540, n19541, n19542, n19543, n19544, n19545,
         n19546, n19547, n19548, n19549, n19550, n19551, n19552, n19553,
         n19554, n19555, n19556, n19557, n19558, n19559, n19560, n19561,
         n19562, n19563, n19564, n19565, n19566, n19567, n19568, n19569,
         n19570, n19571, n19572, n19573, n19574, n19575, n19576, n19577,
         n19578, n19579, n19580, n19581, n19582, n19583, n19584, n19585,
         n19586, n19587, n19588, n19589, n19590, n19591, n19592, n19593,
         n19594, n19595, n19596, n19597, n19598, n19599, n19600, n19601,
         n19602, n19603, n19604, n19605, n19606, n19607, n19608, n19609,
         n19610, n19611, n19612, n19613, n19614, n19615, n19616, n19617,
         n19618, n19619, n19620, n19621, n19622, n19623, n19624, n19625,
         n19626, n19627, n19628, n19629, n19630, n19631, n19632, n19633,
         n19634, n19635, n19636, n19637, n19638, n19639, n19640, n19641,
         n19642, n19643, n19644, n19645, n19646, n19647, n19648, n19649,
         n19650, n19651, n19652, n19653, n19654, n19655, n19656, n19657,
         n19658, n19659, n19660, n19661, n19662, n19663, n19664, n19665,
         n19666, n19667, n19668, n19669, n19670, n19671, n19672, n19673,
         n19674, n19675, n19676, n19677, n19678, n19679, n19680, n19681,
         n19682, n19683, n19684, n19685, n19686, n19687, n19688, n19689,
         n19690, n19691, n19692, n19693, n19694, n19695, n19696, n19697,
         n19698, n19699, n19700, n19701, n19702, n19703, n19704, n19705,
         n19706, n19707, n19708, n19709, n19710, n19711, n19712, n19713,
         n19714, n19715, n19716, n19717, n19718, n19719, n19720, n19721,
         n19722, n19723, n19724, n19725, n19726, n19727, n19728, n19729,
         n19730, n19731, n19732, n19733, n19734, n19735, n19736, n19737,
         n19738, n19739, n19740, n19741, n19742, n19743, n19744, n19745,
         n19746, n19747, n19748, n19749, n19750, n19751, n19752, n19753,
         n19754, n19755, n19756, n19757, n19758, n19759, n19760, n19761,
         n19762, n19763, n19764, n19765, n19766, n19767, n19768, n19769,
         n19770, n19771, n19772, n19773, n19774, n19775, n19776, n19777,
         n19778, n19779, n19780, n19781, n19782, n19783, n19784, n19785,
         n19786, n19787, n19788, n19789, n19790, n19791, n19792, n19793,
         n19794, n19795, n19796, n19797, n19798, n19799, n19800, n19801,
         n19802, n19803, n19804, n19805, n19806, n19807, n19808, n19809,
         n19810, n19811, n19812, n19813, n19814, n19815, n19816, n19817,
         n19818, n19819, n19820, n19821, n19822, n19823, n19824, n19825,
         n19826, n19827, n19828, n19829, n19830, n19831, n19832, n19833,
         n19834, n19835, n19836, n19837, n19838, n19839, n19840, n19841,
         n19842, n19843, n19844, n19845, n19846, n19847, n19848, n19849,
         n19850, n19851, n19852, n19853, n19854, n19855, n19856, n19857,
         n19858, n19859, n19860, n19861, n19862, n19863, n19864, n19865,
         n19866, n19867, n19868, n19869, n19870, n19871, n19872, n19873,
         n19874, n19875, n19876, n19877, n19878, n19879, n19880, n19881,
         n19882, n19883, n19884, n19885, n19886, n19887, n19888, n19889,
         n19890, n19891, n19892, n19893, n19894, n19895, n19896, n19897,
         n19898, n19899, n19900, n19901, n19902, n19903, n19904, n19905,
         n19906, n19907, n19908, n19909, n19910, n19911, n19912, n19913,
         n19914, n19915, n19916, n19917, n19918, n19919, n19920, n19921,
         n19922, n19923, n19924, n19925, n19926, n19927, n19928, n19929,
         n19930, n19931, n19932, n19933, n19934, n19935, n19936, n19937,
         n19938, n19939, n19940, n19941, n19942, n19943, n19944, n19945,
         n19946, n19947, n19948, n19949, n19950, n19951, n19952, n19953,
         n19954, n19955, n19956, n19957, n19958, n19959, n19960, n19961,
         n19962, n19963, n19964, n19965, n19966, n19967, n19968, n19969,
         n19970, n19971, n19972, n19973, n19974, n19975, n19976, n19977,
         n19978, n19979, n19980, n19981, n19982, n19983, n19984, n19985,
         n19986, n19987, n19988, n19989, n19990, n19991, n19992, n19993,
         n19994, n19995, n19996, n19997, n19998, n19999, n20000;

  AND U1 ( .A(n1), .B(n2), .Z(o[9]) );
  AND U2 ( .A(p_input[20009]), .B(p_input[10009]), .Z(n2) );
  AND U3 ( .A(p_input[9]), .B(p_input[30009]), .Z(n1) );
  AND U4 ( .A(n3), .B(n4), .Z(o[99]) );
  AND U5 ( .A(p_input[20099]), .B(p_input[10099]), .Z(n4) );
  AND U6 ( .A(p_input[99]), .B(p_input[30099]), .Z(n3) );
  AND U7 ( .A(n5), .B(n6), .Z(o[999]) );
  AND U8 ( .A(p_input[20999]), .B(p_input[10999]), .Z(n6) );
  AND U9 ( .A(p_input[999]), .B(p_input[30999]), .Z(n5) );
  AND U10 ( .A(n7), .B(n8), .Z(o[9999]) );
  AND U11 ( .A(p_input[29999]), .B(p_input[19999]), .Z(n8) );
  AND U12 ( .A(p_input[9999]), .B(p_input[39999]), .Z(n7) );
  AND U13 ( .A(n9), .B(n10), .Z(o[9998]) );
  AND U14 ( .A(p_input[29998]), .B(p_input[19998]), .Z(n10) );
  AND U15 ( .A(p_input[9998]), .B(p_input[39998]), .Z(n9) );
  AND U16 ( .A(n11), .B(n12), .Z(o[9997]) );
  AND U17 ( .A(p_input[29997]), .B(p_input[19997]), .Z(n12) );
  AND U18 ( .A(p_input[9997]), .B(p_input[39997]), .Z(n11) );
  AND U19 ( .A(n13), .B(n14), .Z(o[9996]) );
  AND U20 ( .A(p_input[29996]), .B(p_input[19996]), .Z(n14) );
  AND U21 ( .A(p_input[9996]), .B(p_input[39996]), .Z(n13) );
  AND U22 ( .A(n15), .B(n16), .Z(o[9995]) );
  AND U23 ( .A(p_input[29995]), .B(p_input[19995]), .Z(n16) );
  AND U24 ( .A(p_input[9995]), .B(p_input[39995]), .Z(n15) );
  AND U25 ( .A(n17), .B(n18), .Z(o[9994]) );
  AND U26 ( .A(p_input[29994]), .B(p_input[19994]), .Z(n18) );
  AND U27 ( .A(p_input[9994]), .B(p_input[39994]), .Z(n17) );
  AND U28 ( .A(n19), .B(n20), .Z(o[9993]) );
  AND U29 ( .A(p_input[29993]), .B(p_input[19993]), .Z(n20) );
  AND U30 ( .A(p_input[9993]), .B(p_input[39993]), .Z(n19) );
  AND U31 ( .A(n21), .B(n22), .Z(o[9992]) );
  AND U32 ( .A(p_input[29992]), .B(p_input[19992]), .Z(n22) );
  AND U33 ( .A(p_input[9992]), .B(p_input[39992]), .Z(n21) );
  AND U34 ( .A(n23), .B(n24), .Z(o[9991]) );
  AND U35 ( .A(p_input[29991]), .B(p_input[19991]), .Z(n24) );
  AND U36 ( .A(p_input[9991]), .B(p_input[39991]), .Z(n23) );
  AND U37 ( .A(n25), .B(n26), .Z(o[9990]) );
  AND U38 ( .A(p_input[29990]), .B(p_input[19990]), .Z(n26) );
  AND U39 ( .A(p_input[9990]), .B(p_input[39990]), .Z(n25) );
  AND U40 ( .A(n27), .B(n28), .Z(o[998]) );
  AND U41 ( .A(p_input[20998]), .B(p_input[10998]), .Z(n28) );
  AND U42 ( .A(p_input[998]), .B(p_input[30998]), .Z(n27) );
  AND U43 ( .A(n29), .B(n30), .Z(o[9989]) );
  AND U44 ( .A(p_input[29989]), .B(p_input[19989]), .Z(n30) );
  AND U45 ( .A(p_input[9989]), .B(p_input[39989]), .Z(n29) );
  AND U46 ( .A(n31), .B(n32), .Z(o[9988]) );
  AND U47 ( .A(p_input[29988]), .B(p_input[19988]), .Z(n32) );
  AND U48 ( .A(p_input[9988]), .B(p_input[39988]), .Z(n31) );
  AND U49 ( .A(n33), .B(n34), .Z(o[9987]) );
  AND U50 ( .A(p_input[29987]), .B(p_input[19987]), .Z(n34) );
  AND U51 ( .A(p_input[9987]), .B(p_input[39987]), .Z(n33) );
  AND U52 ( .A(n35), .B(n36), .Z(o[9986]) );
  AND U53 ( .A(p_input[29986]), .B(p_input[19986]), .Z(n36) );
  AND U54 ( .A(p_input[9986]), .B(p_input[39986]), .Z(n35) );
  AND U55 ( .A(n37), .B(n38), .Z(o[9985]) );
  AND U56 ( .A(p_input[29985]), .B(p_input[19985]), .Z(n38) );
  AND U57 ( .A(p_input[9985]), .B(p_input[39985]), .Z(n37) );
  AND U58 ( .A(n39), .B(n40), .Z(o[9984]) );
  AND U59 ( .A(p_input[29984]), .B(p_input[19984]), .Z(n40) );
  AND U60 ( .A(p_input[9984]), .B(p_input[39984]), .Z(n39) );
  AND U61 ( .A(n41), .B(n42), .Z(o[9983]) );
  AND U62 ( .A(p_input[29983]), .B(p_input[19983]), .Z(n42) );
  AND U63 ( .A(p_input[9983]), .B(p_input[39983]), .Z(n41) );
  AND U64 ( .A(n43), .B(n44), .Z(o[9982]) );
  AND U65 ( .A(p_input[29982]), .B(p_input[19982]), .Z(n44) );
  AND U66 ( .A(p_input[9982]), .B(p_input[39982]), .Z(n43) );
  AND U67 ( .A(n45), .B(n46), .Z(o[9981]) );
  AND U68 ( .A(p_input[29981]), .B(p_input[19981]), .Z(n46) );
  AND U69 ( .A(p_input[9981]), .B(p_input[39981]), .Z(n45) );
  AND U70 ( .A(n47), .B(n48), .Z(o[9980]) );
  AND U71 ( .A(p_input[29980]), .B(p_input[19980]), .Z(n48) );
  AND U72 ( .A(p_input[9980]), .B(p_input[39980]), .Z(n47) );
  AND U73 ( .A(n49), .B(n50), .Z(o[997]) );
  AND U74 ( .A(p_input[20997]), .B(p_input[10997]), .Z(n50) );
  AND U75 ( .A(p_input[997]), .B(p_input[30997]), .Z(n49) );
  AND U76 ( .A(n51), .B(n52), .Z(o[9979]) );
  AND U77 ( .A(p_input[29979]), .B(p_input[19979]), .Z(n52) );
  AND U78 ( .A(p_input[9979]), .B(p_input[39979]), .Z(n51) );
  AND U79 ( .A(n53), .B(n54), .Z(o[9978]) );
  AND U80 ( .A(p_input[29978]), .B(p_input[19978]), .Z(n54) );
  AND U81 ( .A(p_input[9978]), .B(p_input[39978]), .Z(n53) );
  AND U82 ( .A(n55), .B(n56), .Z(o[9977]) );
  AND U83 ( .A(p_input[29977]), .B(p_input[19977]), .Z(n56) );
  AND U84 ( .A(p_input[9977]), .B(p_input[39977]), .Z(n55) );
  AND U85 ( .A(n57), .B(n58), .Z(o[9976]) );
  AND U86 ( .A(p_input[29976]), .B(p_input[19976]), .Z(n58) );
  AND U87 ( .A(p_input[9976]), .B(p_input[39976]), .Z(n57) );
  AND U88 ( .A(n59), .B(n60), .Z(o[9975]) );
  AND U89 ( .A(p_input[29975]), .B(p_input[19975]), .Z(n60) );
  AND U90 ( .A(p_input[9975]), .B(p_input[39975]), .Z(n59) );
  AND U91 ( .A(n61), .B(n62), .Z(o[9974]) );
  AND U92 ( .A(p_input[29974]), .B(p_input[19974]), .Z(n62) );
  AND U93 ( .A(p_input[9974]), .B(p_input[39974]), .Z(n61) );
  AND U94 ( .A(n63), .B(n64), .Z(o[9973]) );
  AND U95 ( .A(p_input[29973]), .B(p_input[19973]), .Z(n64) );
  AND U96 ( .A(p_input[9973]), .B(p_input[39973]), .Z(n63) );
  AND U97 ( .A(n65), .B(n66), .Z(o[9972]) );
  AND U98 ( .A(p_input[29972]), .B(p_input[19972]), .Z(n66) );
  AND U99 ( .A(p_input[9972]), .B(p_input[39972]), .Z(n65) );
  AND U100 ( .A(n67), .B(n68), .Z(o[9971]) );
  AND U101 ( .A(p_input[29971]), .B(p_input[19971]), .Z(n68) );
  AND U102 ( .A(p_input[9971]), .B(p_input[39971]), .Z(n67) );
  AND U103 ( .A(n69), .B(n70), .Z(o[9970]) );
  AND U104 ( .A(p_input[29970]), .B(p_input[19970]), .Z(n70) );
  AND U105 ( .A(p_input[9970]), .B(p_input[39970]), .Z(n69) );
  AND U106 ( .A(n71), .B(n72), .Z(o[996]) );
  AND U107 ( .A(p_input[20996]), .B(p_input[10996]), .Z(n72) );
  AND U108 ( .A(p_input[996]), .B(p_input[30996]), .Z(n71) );
  AND U109 ( .A(n73), .B(n74), .Z(o[9969]) );
  AND U110 ( .A(p_input[29969]), .B(p_input[19969]), .Z(n74) );
  AND U111 ( .A(p_input[9969]), .B(p_input[39969]), .Z(n73) );
  AND U112 ( .A(n75), .B(n76), .Z(o[9968]) );
  AND U113 ( .A(p_input[29968]), .B(p_input[19968]), .Z(n76) );
  AND U114 ( .A(p_input[9968]), .B(p_input[39968]), .Z(n75) );
  AND U115 ( .A(n77), .B(n78), .Z(o[9967]) );
  AND U116 ( .A(p_input[29967]), .B(p_input[19967]), .Z(n78) );
  AND U117 ( .A(p_input[9967]), .B(p_input[39967]), .Z(n77) );
  AND U118 ( .A(n79), .B(n80), .Z(o[9966]) );
  AND U119 ( .A(p_input[29966]), .B(p_input[19966]), .Z(n80) );
  AND U120 ( .A(p_input[9966]), .B(p_input[39966]), .Z(n79) );
  AND U121 ( .A(n81), .B(n82), .Z(o[9965]) );
  AND U122 ( .A(p_input[29965]), .B(p_input[19965]), .Z(n82) );
  AND U123 ( .A(p_input[9965]), .B(p_input[39965]), .Z(n81) );
  AND U124 ( .A(n83), .B(n84), .Z(o[9964]) );
  AND U125 ( .A(p_input[29964]), .B(p_input[19964]), .Z(n84) );
  AND U126 ( .A(p_input[9964]), .B(p_input[39964]), .Z(n83) );
  AND U127 ( .A(n85), .B(n86), .Z(o[9963]) );
  AND U128 ( .A(p_input[29963]), .B(p_input[19963]), .Z(n86) );
  AND U129 ( .A(p_input[9963]), .B(p_input[39963]), .Z(n85) );
  AND U130 ( .A(n87), .B(n88), .Z(o[9962]) );
  AND U131 ( .A(p_input[29962]), .B(p_input[19962]), .Z(n88) );
  AND U132 ( .A(p_input[9962]), .B(p_input[39962]), .Z(n87) );
  AND U133 ( .A(n89), .B(n90), .Z(o[9961]) );
  AND U134 ( .A(p_input[29961]), .B(p_input[19961]), .Z(n90) );
  AND U135 ( .A(p_input[9961]), .B(p_input[39961]), .Z(n89) );
  AND U136 ( .A(n91), .B(n92), .Z(o[9960]) );
  AND U137 ( .A(p_input[29960]), .B(p_input[19960]), .Z(n92) );
  AND U138 ( .A(p_input[9960]), .B(p_input[39960]), .Z(n91) );
  AND U139 ( .A(n93), .B(n94), .Z(o[995]) );
  AND U140 ( .A(p_input[20995]), .B(p_input[10995]), .Z(n94) );
  AND U141 ( .A(p_input[995]), .B(p_input[30995]), .Z(n93) );
  AND U142 ( .A(n95), .B(n96), .Z(o[9959]) );
  AND U143 ( .A(p_input[29959]), .B(p_input[19959]), .Z(n96) );
  AND U144 ( .A(p_input[9959]), .B(p_input[39959]), .Z(n95) );
  AND U145 ( .A(n97), .B(n98), .Z(o[9958]) );
  AND U146 ( .A(p_input[29958]), .B(p_input[19958]), .Z(n98) );
  AND U147 ( .A(p_input[9958]), .B(p_input[39958]), .Z(n97) );
  AND U148 ( .A(n99), .B(n100), .Z(o[9957]) );
  AND U149 ( .A(p_input[29957]), .B(p_input[19957]), .Z(n100) );
  AND U150 ( .A(p_input[9957]), .B(p_input[39957]), .Z(n99) );
  AND U151 ( .A(n101), .B(n102), .Z(o[9956]) );
  AND U152 ( .A(p_input[29956]), .B(p_input[19956]), .Z(n102) );
  AND U153 ( .A(p_input[9956]), .B(p_input[39956]), .Z(n101) );
  AND U154 ( .A(n103), .B(n104), .Z(o[9955]) );
  AND U155 ( .A(p_input[29955]), .B(p_input[19955]), .Z(n104) );
  AND U156 ( .A(p_input[9955]), .B(p_input[39955]), .Z(n103) );
  AND U157 ( .A(n105), .B(n106), .Z(o[9954]) );
  AND U158 ( .A(p_input[29954]), .B(p_input[19954]), .Z(n106) );
  AND U159 ( .A(p_input[9954]), .B(p_input[39954]), .Z(n105) );
  AND U160 ( .A(n107), .B(n108), .Z(o[9953]) );
  AND U161 ( .A(p_input[29953]), .B(p_input[19953]), .Z(n108) );
  AND U162 ( .A(p_input[9953]), .B(p_input[39953]), .Z(n107) );
  AND U163 ( .A(n109), .B(n110), .Z(o[9952]) );
  AND U164 ( .A(p_input[29952]), .B(p_input[19952]), .Z(n110) );
  AND U165 ( .A(p_input[9952]), .B(p_input[39952]), .Z(n109) );
  AND U166 ( .A(n111), .B(n112), .Z(o[9951]) );
  AND U167 ( .A(p_input[29951]), .B(p_input[19951]), .Z(n112) );
  AND U168 ( .A(p_input[9951]), .B(p_input[39951]), .Z(n111) );
  AND U169 ( .A(n113), .B(n114), .Z(o[9950]) );
  AND U170 ( .A(p_input[29950]), .B(p_input[19950]), .Z(n114) );
  AND U171 ( .A(p_input[9950]), .B(p_input[39950]), .Z(n113) );
  AND U172 ( .A(n115), .B(n116), .Z(o[994]) );
  AND U173 ( .A(p_input[20994]), .B(p_input[10994]), .Z(n116) );
  AND U174 ( .A(p_input[994]), .B(p_input[30994]), .Z(n115) );
  AND U175 ( .A(n117), .B(n118), .Z(o[9949]) );
  AND U176 ( .A(p_input[29949]), .B(p_input[19949]), .Z(n118) );
  AND U177 ( .A(p_input[9949]), .B(p_input[39949]), .Z(n117) );
  AND U178 ( .A(n119), .B(n120), .Z(o[9948]) );
  AND U179 ( .A(p_input[29948]), .B(p_input[19948]), .Z(n120) );
  AND U180 ( .A(p_input[9948]), .B(p_input[39948]), .Z(n119) );
  AND U181 ( .A(n121), .B(n122), .Z(o[9947]) );
  AND U182 ( .A(p_input[29947]), .B(p_input[19947]), .Z(n122) );
  AND U183 ( .A(p_input[9947]), .B(p_input[39947]), .Z(n121) );
  AND U184 ( .A(n123), .B(n124), .Z(o[9946]) );
  AND U185 ( .A(p_input[29946]), .B(p_input[19946]), .Z(n124) );
  AND U186 ( .A(p_input[9946]), .B(p_input[39946]), .Z(n123) );
  AND U187 ( .A(n125), .B(n126), .Z(o[9945]) );
  AND U188 ( .A(p_input[29945]), .B(p_input[19945]), .Z(n126) );
  AND U189 ( .A(p_input[9945]), .B(p_input[39945]), .Z(n125) );
  AND U190 ( .A(n127), .B(n128), .Z(o[9944]) );
  AND U191 ( .A(p_input[29944]), .B(p_input[19944]), .Z(n128) );
  AND U192 ( .A(p_input[9944]), .B(p_input[39944]), .Z(n127) );
  AND U193 ( .A(n129), .B(n130), .Z(o[9943]) );
  AND U194 ( .A(p_input[29943]), .B(p_input[19943]), .Z(n130) );
  AND U195 ( .A(p_input[9943]), .B(p_input[39943]), .Z(n129) );
  AND U196 ( .A(n131), .B(n132), .Z(o[9942]) );
  AND U197 ( .A(p_input[29942]), .B(p_input[19942]), .Z(n132) );
  AND U198 ( .A(p_input[9942]), .B(p_input[39942]), .Z(n131) );
  AND U199 ( .A(n133), .B(n134), .Z(o[9941]) );
  AND U200 ( .A(p_input[29941]), .B(p_input[19941]), .Z(n134) );
  AND U201 ( .A(p_input[9941]), .B(p_input[39941]), .Z(n133) );
  AND U202 ( .A(n135), .B(n136), .Z(o[9940]) );
  AND U203 ( .A(p_input[29940]), .B(p_input[19940]), .Z(n136) );
  AND U204 ( .A(p_input[9940]), .B(p_input[39940]), .Z(n135) );
  AND U205 ( .A(n137), .B(n138), .Z(o[993]) );
  AND U206 ( .A(p_input[20993]), .B(p_input[10993]), .Z(n138) );
  AND U207 ( .A(p_input[993]), .B(p_input[30993]), .Z(n137) );
  AND U208 ( .A(n139), .B(n140), .Z(o[9939]) );
  AND U209 ( .A(p_input[29939]), .B(p_input[19939]), .Z(n140) );
  AND U210 ( .A(p_input[9939]), .B(p_input[39939]), .Z(n139) );
  AND U211 ( .A(n141), .B(n142), .Z(o[9938]) );
  AND U212 ( .A(p_input[29938]), .B(p_input[19938]), .Z(n142) );
  AND U213 ( .A(p_input[9938]), .B(p_input[39938]), .Z(n141) );
  AND U214 ( .A(n143), .B(n144), .Z(o[9937]) );
  AND U215 ( .A(p_input[29937]), .B(p_input[19937]), .Z(n144) );
  AND U216 ( .A(p_input[9937]), .B(p_input[39937]), .Z(n143) );
  AND U217 ( .A(n145), .B(n146), .Z(o[9936]) );
  AND U218 ( .A(p_input[29936]), .B(p_input[19936]), .Z(n146) );
  AND U219 ( .A(p_input[9936]), .B(p_input[39936]), .Z(n145) );
  AND U220 ( .A(n147), .B(n148), .Z(o[9935]) );
  AND U221 ( .A(p_input[29935]), .B(p_input[19935]), .Z(n148) );
  AND U222 ( .A(p_input[9935]), .B(p_input[39935]), .Z(n147) );
  AND U223 ( .A(n149), .B(n150), .Z(o[9934]) );
  AND U224 ( .A(p_input[29934]), .B(p_input[19934]), .Z(n150) );
  AND U225 ( .A(p_input[9934]), .B(p_input[39934]), .Z(n149) );
  AND U226 ( .A(n151), .B(n152), .Z(o[9933]) );
  AND U227 ( .A(p_input[29933]), .B(p_input[19933]), .Z(n152) );
  AND U228 ( .A(p_input[9933]), .B(p_input[39933]), .Z(n151) );
  AND U229 ( .A(n153), .B(n154), .Z(o[9932]) );
  AND U230 ( .A(p_input[29932]), .B(p_input[19932]), .Z(n154) );
  AND U231 ( .A(p_input[9932]), .B(p_input[39932]), .Z(n153) );
  AND U232 ( .A(n155), .B(n156), .Z(o[9931]) );
  AND U233 ( .A(p_input[29931]), .B(p_input[19931]), .Z(n156) );
  AND U234 ( .A(p_input[9931]), .B(p_input[39931]), .Z(n155) );
  AND U235 ( .A(n157), .B(n158), .Z(o[9930]) );
  AND U236 ( .A(p_input[29930]), .B(p_input[19930]), .Z(n158) );
  AND U237 ( .A(p_input[9930]), .B(p_input[39930]), .Z(n157) );
  AND U238 ( .A(n159), .B(n160), .Z(o[992]) );
  AND U239 ( .A(p_input[20992]), .B(p_input[10992]), .Z(n160) );
  AND U240 ( .A(p_input[992]), .B(p_input[30992]), .Z(n159) );
  AND U241 ( .A(n161), .B(n162), .Z(o[9929]) );
  AND U242 ( .A(p_input[29929]), .B(p_input[19929]), .Z(n162) );
  AND U243 ( .A(p_input[9929]), .B(p_input[39929]), .Z(n161) );
  AND U244 ( .A(n163), .B(n164), .Z(o[9928]) );
  AND U245 ( .A(p_input[29928]), .B(p_input[19928]), .Z(n164) );
  AND U246 ( .A(p_input[9928]), .B(p_input[39928]), .Z(n163) );
  AND U247 ( .A(n165), .B(n166), .Z(o[9927]) );
  AND U248 ( .A(p_input[29927]), .B(p_input[19927]), .Z(n166) );
  AND U249 ( .A(p_input[9927]), .B(p_input[39927]), .Z(n165) );
  AND U250 ( .A(n167), .B(n168), .Z(o[9926]) );
  AND U251 ( .A(p_input[29926]), .B(p_input[19926]), .Z(n168) );
  AND U252 ( .A(p_input[9926]), .B(p_input[39926]), .Z(n167) );
  AND U253 ( .A(n169), .B(n170), .Z(o[9925]) );
  AND U254 ( .A(p_input[29925]), .B(p_input[19925]), .Z(n170) );
  AND U255 ( .A(p_input[9925]), .B(p_input[39925]), .Z(n169) );
  AND U256 ( .A(n171), .B(n172), .Z(o[9924]) );
  AND U257 ( .A(p_input[29924]), .B(p_input[19924]), .Z(n172) );
  AND U258 ( .A(p_input[9924]), .B(p_input[39924]), .Z(n171) );
  AND U259 ( .A(n173), .B(n174), .Z(o[9923]) );
  AND U260 ( .A(p_input[29923]), .B(p_input[19923]), .Z(n174) );
  AND U261 ( .A(p_input[9923]), .B(p_input[39923]), .Z(n173) );
  AND U262 ( .A(n175), .B(n176), .Z(o[9922]) );
  AND U263 ( .A(p_input[29922]), .B(p_input[19922]), .Z(n176) );
  AND U264 ( .A(p_input[9922]), .B(p_input[39922]), .Z(n175) );
  AND U265 ( .A(n177), .B(n178), .Z(o[9921]) );
  AND U266 ( .A(p_input[29921]), .B(p_input[19921]), .Z(n178) );
  AND U267 ( .A(p_input[9921]), .B(p_input[39921]), .Z(n177) );
  AND U268 ( .A(n179), .B(n180), .Z(o[9920]) );
  AND U269 ( .A(p_input[29920]), .B(p_input[19920]), .Z(n180) );
  AND U270 ( .A(p_input[9920]), .B(p_input[39920]), .Z(n179) );
  AND U271 ( .A(n181), .B(n182), .Z(o[991]) );
  AND U272 ( .A(p_input[20991]), .B(p_input[10991]), .Z(n182) );
  AND U273 ( .A(p_input[991]), .B(p_input[30991]), .Z(n181) );
  AND U274 ( .A(n183), .B(n184), .Z(o[9919]) );
  AND U275 ( .A(p_input[29919]), .B(p_input[19919]), .Z(n184) );
  AND U276 ( .A(p_input[9919]), .B(p_input[39919]), .Z(n183) );
  AND U277 ( .A(n185), .B(n186), .Z(o[9918]) );
  AND U278 ( .A(p_input[29918]), .B(p_input[19918]), .Z(n186) );
  AND U279 ( .A(p_input[9918]), .B(p_input[39918]), .Z(n185) );
  AND U280 ( .A(n187), .B(n188), .Z(o[9917]) );
  AND U281 ( .A(p_input[29917]), .B(p_input[19917]), .Z(n188) );
  AND U282 ( .A(p_input[9917]), .B(p_input[39917]), .Z(n187) );
  AND U283 ( .A(n189), .B(n190), .Z(o[9916]) );
  AND U284 ( .A(p_input[29916]), .B(p_input[19916]), .Z(n190) );
  AND U285 ( .A(p_input[9916]), .B(p_input[39916]), .Z(n189) );
  AND U286 ( .A(n191), .B(n192), .Z(o[9915]) );
  AND U287 ( .A(p_input[29915]), .B(p_input[19915]), .Z(n192) );
  AND U288 ( .A(p_input[9915]), .B(p_input[39915]), .Z(n191) );
  AND U289 ( .A(n193), .B(n194), .Z(o[9914]) );
  AND U290 ( .A(p_input[29914]), .B(p_input[19914]), .Z(n194) );
  AND U291 ( .A(p_input[9914]), .B(p_input[39914]), .Z(n193) );
  AND U292 ( .A(n195), .B(n196), .Z(o[9913]) );
  AND U293 ( .A(p_input[29913]), .B(p_input[19913]), .Z(n196) );
  AND U294 ( .A(p_input[9913]), .B(p_input[39913]), .Z(n195) );
  AND U295 ( .A(n197), .B(n198), .Z(o[9912]) );
  AND U296 ( .A(p_input[29912]), .B(p_input[19912]), .Z(n198) );
  AND U297 ( .A(p_input[9912]), .B(p_input[39912]), .Z(n197) );
  AND U298 ( .A(n199), .B(n200), .Z(o[9911]) );
  AND U299 ( .A(p_input[29911]), .B(p_input[19911]), .Z(n200) );
  AND U300 ( .A(p_input[9911]), .B(p_input[39911]), .Z(n199) );
  AND U301 ( .A(n201), .B(n202), .Z(o[9910]) );
  AND U302 ( .A(p_input[29910]), .B(p_input[19910]), .Z(n202) );
  AND U303 ( .A(p_input[9910]), .B(p_input[39910]), .Z(n201) );
  AND U304 ( .A(n203), .B(n204), .Z(o[990]) );
  AND U305 ( .A(p_input[20990]), .B(p_input[10990]), .Z(n204) );
  AND U306 ( .A(p_input[990]), .B(p_input[30990]), .Z(n203) );
  AND U307 ( .A(n205), .B(n206), .Z(o[9909]) );
  AND U308 ( .A(p_input[29909]), .B(p_input[19909]), .Z(n206) );
  AND U309 ( .A(p_input[9909]), .B(p_input[39909]), .Z(n205) );
  AND U310 ( .A(n207), .B(n208), .Z(o[9908]) );
  AND U311 ( .A(p_input[29908]), .B(p_input[19908]), .Z(n208) );
  AND U312 ( .A(p_input[9908]), .B(p_input[39908]), .Z(n207) );
  AND U313 ( .A(n209), .B(n210), .Z(o[9907]) );
  AND U314 ( .A(p_input[29907]), .B(p_input[19907]), .Z(n210) );
  AND U315 ( .A(p_input[9907]), .B(p_input[39907]), .Z(n209) );
  AND U316 ( .A(n211), .B(n212), .Z(o[9906]) );
  AND U317 ( .A(p_input[29906]), .B(p_input[19906]), .Z(n212) );
  AND U318 ( .A(p_input[9906]), .B(p_input[39906]), .Z(n211) );
  AND U319 ( .A(n213), .B(n214), .Z(o[9905]) );
  AND U320 ( .A(p_input[29905]), .B(p_input[19905]), .Z(n214) );
  AND U321 ( .A(p_input[9905]), .B(p_input[39905]), .Z(n213) );
  AND U322 ( .A(n215), .B(n216), .Z(o[9904]) );
  AND U323 ( .A(p_input[29904]), .B(p_input[19904]), .Z(n216) );
  AND U324 ( .A(p_input[9904]), .B(p_input[39904]), .Z(n215) );
  AND U325 ( .A(n217), .B(n218), .Z(o[9903]) );
  AND U326 ( .A(p_input[29903]), .B(p_input[19903]), .Z(n218) );
  AND U327 ( .A(p_input[9903]), .B(p_input[39903]), .Z(n217) );
  AND U328 ( .A(n219), .B(n220), .Z(o[9902]) );
  AND U329 ( .A(p_input[29902]), .B(p_input[19902]), .Z(n220) );
  AND U330 ( .A(p_input[9902]), .B(p_input[39902]), .Z(n219) );
  AND U331 ( .A(n221), .B(n222), .Z(o[9901]) );
  AND U332 ( .A(p_input[29901]), .B(p_input[19901]), .Z(n222) );
  AND U333 ( .A(p_input[9901]), .B(p_input[39901]), .Z(n221) );
  AND U334 ( .A(n223), .B(n224), .Z(o[9900]) );
  AND U335 ( .A(p_input[29900]), .B(p_input[19900]), .Z(n224) );
  AND U336 ( .A(p_input[9900]), .B(p_input[39900]), .Z(n223) );
  AND U337 ( .A(n225), .B(n226), .Z(o[98]) );
  AND U338 ( .A(p_input[20098]), .B(p_input[10098]), .Z(n226) );
  AND U339 ( .A(p_input[98]), .B(p_input[30098]), .Z(n225) );
  AND U340 ( .A(n227), .B(n228), .Z(o[989]) );
  AND U341 ( .A(p_input[20989]), .B(p_input[10989]), .Z(n228) );
  AND U342 ( .A(p_input[989]), .B(p_input[30989]), .Z(n227) );
  AND U343 ( .A(n229), .B(n230), .Z(o[9899]) );
  AND U344 ( .A(p_input[29899]), .B(p_input[19899]), .Z(n230) );
  AND U345 ( .A(p_input[9899]), .B(p_input[39899]), .Z(n229) );
  AND U346 ( .A(n231), .B(n232), .Z(o[9898]) );
  AND U347 ( .A(p_input[29898]), .B(p_input[19898]), .Z(n232) );
  AND U348 ( .A(p_input[9898]), .B(p_input[39898]), .Z(n231) );
  AND U349 ( .A(n233), .B(n234), .Z(o[9897]) );
  AND U350 ( .A(p_input[29897]), .B(p_input[19897]), .Z(n234) );
  AND U351 ( .A(p_input[9897]), .B(p_input[39897]), .Z(n233) );
  AND U352 ( .A(n235), .B(n236), .Z(o[9896]) );
  AND U353 ( .A(p_input[29896]), .B(p_input[19896]), .Z(n236) );
  AND U354 ( .A(p_input[9896]), .B(p_input[39896]), .Z(n235) );
  AND U355 ( .A(n237), .B(n238), .Z(o[9895]) );
  AND U356 ( .A(p_input[29895]), .B(p_input[19895]), .Z(n238) );
  AND U357 ( .A(p_input[9895]), .B(p_input[39895]), .Z(n237) );
  AND U358 ( .A(n239), .B(n240), .Z(o[9894]) );
  AND U359 ( .A(p_input[29894]), .B(p_input[19894]), .Z(n240) );
  AND U360 ( .A(p_input[9894]), .B(p_input[39894]), .Z(n239) );
  AND U361 ( .A(n241), .B(n242), .Z(o[9893]) );
  AND U362 ( .A(p_input[29893]), .B(p_input[19893]), .Z(n242) );
  AND U363 ( .A(p_input[9893]), .B(p_input[39893]), .Z(n241) );
  AND U364 ( .A(n243), .B(n244), .Z(o[9892]) );
  AND U365 ( .A(p_input[29892]), .B(p_input[19892]), .Z(n244) );
  AND U366 ( .A(p_input[9892]), .B(p_input[39892]), .Z(n243) );
  AND U367 ( .A(n245), .B(n246), .Z(o[9891]) );
  AND U368 ( .A(p_input[29891]), .B(p_input[19891]), .Z(n246) );
  AND U369 ( .A(p_input[9891]), .B(p_input[39891]), .Z(n245) );
  AND U370 ( .A(n247), .B(n248), .Z(o[9890]) );
  AND U371 ( .A(p_input[29890]), .B(p_input[19890]), .Z(n248) );
  AND U372 ( .A(p_input[9890]), .B(p_input[39890]), .Z(n247) );
  AND U373 ( .A(n249), .B(n250), .Z(o[988]) );
  AND U374 ( .A(p_input[20988]), .B(p_input[10988]), .Z(n250) );
  AND U375 ( .A(p_input[988]), .B(p_input[30988]), .Z(n249) );
  AND U376 ( .A(n251), .B(n252), .Z(o[9889]) );
  AND U377 ( .A(p_input[29889]), .B(p_input[19889]), .Z(n252) );
  AND U378 ( .A(p_input[9889]), .B(p_input[39889]), .Z(n251) );
  AND U379 ( .A(n253), .B(n254), .Z(o[9888]) );
  AND U380 ( .A(p_input[29888]), .B(p_input[19888]), .Z(n254) );
  AND U381 ( .A(p_input[9888]), .B(p_input[39888]), .Z(n253) );
  AND U382 ( .A(n255), .B(n256), .Z(o[9887]) );
  AND U383 ( .A(p_input[29887]), .B(p_input[19887]), .Z(n256) );
  AND U384 ( .A(p_input[9887]), .B(p_input[39887]), .Z(n255) );
  AND U385 ( .A(n257), .B(n258), .Z(o[9886]) );
  AND U386 ( .A(p_input[29886]), .B(p_input[19886]), .Z(n258) );
  AND U387 ( .A(p_input[9886]), .B(p_input[39886]), .Z(n257) );
  AND U388 ( .A(n259), .B(n260), .Z(o[9885]) );
  AND U389 ( .A(p_input[29885]), .B(p_input[19885]), .Z(n260) );
  AND U390 ( .A(p_input[9885]), .B(p_input[39885]), .Z(n259) );
  AND U391 ( .A(n261), .B(n262), .Z(o[9884]) );
  AND U392 ( .A(p_input[29884]), .B(p_input[19884]), .Z(n262) );
  AND U393 ( .A(p_input[9884]), .B(p_input[39884]), .Z(n261) );
  AND U394 ( .A(n263), .B(n264), .Z(o[9883]) );
  AND U395 ( .A(p_input[29883]), .B(p_input[19883]), .Z(n264) );
  AND U396 ( .A(p_input[9883]), .B(p_input[39883]), .Z(n263) );
  AND U397 ( .A(n265), .B(n266), .Z(o[9882]) );
  AND U398 ( .A(p_input[29882]), .B(p_input[19882]), .Z(n266) );
  AND U399 ( .A(p_input[9882]), .B(p_input[39882]), .Z(n265) );
  AND U400 ( .A(n267), .B(n268), .Z(o[9881]) );
  AND U401 ( .A(p_input[29881]), .B(p_input[19881]), .Z(n268) );
  AND U402 ( .A(p_input[9881]), .B(p_input[39881]), .Z(n267) );
  AND U403 ( .A(n269), .B(n270), .Z(o[9880]) );
  AND U404 ( .A(p_input[29880]), .B(p_input[19880]), .Z(n270) );
  AND U405 ( .A(p_input[9880]), .B(p_input[39880]), .Z(n269) );
  AND U406 ( .A(n271), .B(n272), .Z(o[987]) );
  AND U407 ( .A(p_input[20987]), .B(p_input[10987]), .Z(n272) );
  AND U408 ( .A(p_input[987]), .B(p_input[30987]), .Z(n271) );
  AND U409 ( .A(n273), .B(n274), .Z(o[9879]) );
  AND U410 ( .A(p_input[29879]), .B(p_input[19879]), .Z(n274) );
  AND U411 ( .A(p_input[9879]), .B(p_input[39879]), .Z(n273) );
  AND U412 ( .A(n275), .B(n276), .Z(o[9878]) );
  AND U413 ( .A(p_input[29878]), .B(p_input[19878]), .Z(n276) );
  AND U414 ( .A(p_input[9878]), .B(p_input[39878]), .Z(n275) );
  AND U415 ( .A(n277), .B(n278), .Z(o[9877]) );
  AND U416 ( .A(p_input[29877]), .B(p_input[19877]), .Z(n278) );
  AND U417 ( .A(p_input[9877]), .B(p_input[39877]), .Z(n277) );
  AND U418 ( .A(n279), .B(n280), .Z(o[9876]) );
  AND U419 ( .A(p_input[29876]), .B(p_input[19876]), .Z(n280) );
  AND U420 ( .A(p_input[9876]), .B(p_input[39876]), .Z(n279) );
  AND U421 ( .A(n281), .B(n282), .Z(o[9875]) );
  AND U422 ( .A(p_input[29875]), .B(p_input[19875]), .Z(n282) );
  AND U423 ( .A(p_input[9875]), .B(p_input[39875]), .Z(n281) );
  AND U424 ( .A(n283), .B(n284), .Z(o[9874]) );
  AND U425 ( .A(p_input[29874]), .B(p_input[19874]), .Z(n284) );
  AND U426 ( .A(p_input[9874]), .B(p_input[39874]), .Z(n283) );
  AND U427 ( .A(n285), .B(n286), .Z(o[9873]) );
  AND U428 ( .A(p_input[29873]), .B(p_input[19873]), .Z(n286) );
  AND U429 ( .A(p_input[9873]), .B(p_input[39873]), .Z(n285) );
  AND U430 ( .A(n287), .B(n288), .Z(o[9872]) );
  AND U431 ( .A(p_input[29872]), .B(p_input[19872]), .Z(n288) );
  AND U432 ( .A(p_input[9872]), .B(p_input[39872]), .Z(n287) );
  AND U433 ( .A(n289), .B(n290), .Z(o[9871]) );
  AND U434 ( .A(p_input[29871]), .B(p_input[19871]), .Z(n290) );
  AND U435 ( .A(p_input[9871]), .B(p_input[39871]), .Z(n289) );
  AND U436 ( .A(n291), .B(n292), .Z(o[9870]) );
  AND U437 ( .A(p_input[29870]), .B(p_input[19870]), .Z(n292) );
  AND U438 ( .A(p_input[9870]), .B(p_input[39870]), .Z(n291) );
  AND U439 ( .A(n293), .B(n294), .Z(o[986]) );
  AND U440 ( .A(p_input[20986]), .B(p_input[10986]), .Z(n294) );
  AND U441 ( .A(p_input[986]), .B(p_input[30986]), .Z(n293) );
  AND U442 ( .A(n295), .B(n296), .Z(o[9869]) );
  AND U443 ( .A(p_input[29869]), .B(p_input[19869]), .Z(n296) );
  AND U444 ( .A(p_input[9869]), .B(p_input[39869]), .Z(n295) );
  AND U445 ( .A(n297), .B(n298), .Z(o[9868]) );
  AND U446 ( .A(p_input[29868]), .B(p_input[19868]), .Z(n298) );
  AND U447 ( .A(p_input[9868]), .B(p_input[39868]), .Z(n297) );
  AND U448 ( .A(n299), .B(n300), .Z(o[9867]) );
  AND U449 ( .A(p_input[29867]), .B(p_input[19867]), .Z(n300) );
  AND U450 ( .A(p_input[9867]), .B(p_input[39867]), .Z(n299) );
  AND U451 ( .A(n301), .B(n302), .Z(o[9866]) );
  AND U452 ( .A(p_input[29866]), .B(p_input[19866]), .Z(n302) );
  AND U453 ( .A(p_input[9866]), .B(p_input[39866]), .Z(n301) );
  AND U454 ( .A(n303), .B(n304), .Z(o[9865]) );
  AND U455 ( .A(p_input[29865]), .B(p_input[19865]), .Z(n304) );
  AND U456 ( .A(p_input[9865]), .B(p_input[39865]), .Z(n303) );
  AND U457 ( .A(n305), .B(n306), .Z(o[9864]) );
  AND U458 ( .A(p_input[29864]), .B(p_input[19864]), .Z(n306) );
  AND U459 ( .A(p_input[9864]), .B(p_input[39864]), .Z(n305) );
  AND U460 ( .A(n307), .B(n308), .Z(o[9863]) );
  AND U461 ( .A(p_input[29863]), .B(p_input[19863]), .Z(n308) );
  AND U462 ( .A(p_input[9863]), .B(p_input[39863]), .Z(n307) );
  AND U463 ( .A(n309), .B(n310), .Z(o[9862]) );
  AND U464 ( .A(p_input[29862]), .B(p_input[19862]), .Z(n310) );
  AND U465 ( .A(p_input[9862]), .B(p_input[39862]), .Z(n309) );
  AND U466 ( .A(n311), .B(n312), .Z(o[9861]) );
  AND U467 ( .A(p_input[29861]), .B(p_input[19861]), .Z(n312) );
  AND U468 ( .A(p_input[9861]), .B(p_input[39861]), .Z(n311) );
  AND U469 ( .A(n313), .B(n314), .Z(o[9860]) );
  AND U470 ( .A(p_input[29860]), .B(p_input[19860]), .Z(n314) );
  AND U471 ( .A(p_input[9860]), .B(p_input[39860]), .Z(n313) );
  AND U472 ( .A(n315), .B(n316), .Z(o[985]) );
  AND U473 ( .A(p_input[20985]), .B(p_input[10985]), .Z(n316) );
  AND U474 ( .A(p_input[985]), .B(p_input[30985]), .Z(n315) );
  AND U475 ( .A(n317), .B(n318), .Z(o[9859]) );
  AND U476 ( .A(p_input[29859]), .B(p_input[19859]), .Z(n318) );
  AND U477 ( .A(p_input[9859]), .B(p_input[39859]), .Z(n317) );
  AND U478 ( .A(n319), .B(n320), .Z(o[9858]) );
  AND U479 ( .A(p_input[29858]), .B(p_input[19858]), .Z(n320) );
  AND U480 ( .A(p_input[9858]), .B(p_input[39858]), .Z(n319) );
  AND U481 ( .A(n321), .B(n322), .Z(o[9857]) );
  AND U482 ( .A(p_input[29857]), .B(p_input[19857]), .Z(n322) );
  AND U483 ( .A(p_input[9857]), .B(p_input[39857]), .Z(n321) );
  AND U484 ( .A(n323), .B(n324), .Z(o[9856]) );
  AND U485 ( .A(p_input[29856]), .B(p_input[19856]), .Z(n324) );
  AND U486 ( .A(p_input[9856]), .B(p_input[39856]), .Z(n323) );
  AND U487 ( .A(n325), .B(n326), .Z(o[9855]) );
  AND U488 ( .A(p_input[29855]), .B(p_input[19855]), .Z(n326) );
  AND U489 ( .A(p_input[9855]), .B(p_input[39855]), .Z(n325) );
  AND U490 ( .A(n327), .B(n328), .Z(o[9854]) );
  AND U491 ( .A(p_input[29854]), .B(p_input[19854]), .Z(n328) );
  AND U492 ( .A(p_input[9854]), .B(p_input[39854]), .Z(n327) );
  AND U493 ( .A(n329), .B(n330), .Z(o[9853]) );
  AND U494 ( .A(p_input[29853]), .B(p_input[19853]), .Z(n330) );
  AND U495 ( .A(p_input[9853]), .B(p_input[39853]), .Z(n329) );
  AND U496 ( .A(n331), .B(n332), .Z(o[9852]) );
  AND U497 ( .A(p_input[29852]), .B(p_input[19852]), .Z(n332) );
  AND U498 ( .A(p_input[9852]), .B(p_input[39852]), .Z(n331) );
  AND U499 ( .A(n333), .B(n334), .Z(o[9851]) );
  AND U500 ( .A(p_input[29851]), .B(p_input[19851]), .Z(n334) );
  AND U501 ( .A(p_input[9851]), .B(p_input[39851]), .Z(n333) );
  AND U502 ( .A(n335), .B(n336), .Z(o[9850]) );
  AND U503 ( .A(p_input[29850]), .B(p_input[19850]), .Z(n336) );
  AND U504 ( .A(p_input[9850]), .B(p_input[39850]), .Z(n335) );
  AND U505 ( .A(n337), .B(n338), .Z(o[984]) );
  AND U506 ( .A(p_input[20984]), .B(p_input[10984]), .Z(n338) );
  AND U507 ( .A(p_input[984]), .B(p_input[30984]), .Z(n337) );
  AND U508 ( .A(n339), .B(n340), .Z(o[9849]) );
  AND U509 ( .A(p_input[29849]), .B(p_input[19849]), .Z(n340) );
  AND U510 ( .A(p_input[9849]), .B(p_input[39849]), .Z(n339) );
  AND U511 ( .A(n341), .B(n342), .Z(o[9848]) );
  AND U512 ( .A(p_input[29848]), .B(p_input[19848]), .Z(n342) );
  AND U513 ( .A(p_input[9848]), .B(p_input[39848]), .Z(n341) );
  AND U514 ( .A(n343), .B(n344), .Z(o[9847]) );
  AND U515 ( .A(p_input[29847]), .B(p_input[19847]), .Z(n344) );
  AND U516 ( .A(p_input[9847]), .B(p_input[39847]), .Z(n343) );
  AND U517 ( .A(n345), .B(n346), .Z(o[9846]) );
  AND U518 ( .A(p_input[29846]), .B(p_input[19846]), .Z(n346) );
  AND U519 ( .A(p_input[9846]), .B(p_input[39846]), .Z(n345) );
  AND U520 ( .A(n347), .B(n348), .Z(o[9845]) );
  AND U521 ( .A(p_input[29845]), .B(p_input[19845]), .Z(n348) );
  AND U522 ( .A(p_input[9845]), .B(p_input[39845]), .Z(n347) );
  AND U523 ( .A(n349), .B(n350), .Z(o[9844]) );
  AND U524 ( .A(p_input[29844]), .B(p_input[19844]), .Z(n350) );
  AND U525 ( .A(p_input[9844]), .B(p_input[39844]), .Z(n349) );
  AND U526 ( .A(n351), .B(n352), .Z(o[9843]) );
  AND U527 ( .A(p_input[29843]), .B(p_input[19843]), .Z(n352) );
  AND U528 ( .A(p_input[9843]), .B(p_input[39843]), .Z(n351) );
  AND U529 ( .A(n353), .B(n354), .Z(o[9842]) );
  AND U530 ( .A(p_input[29842]), .B(p_input[19842]), .Z(n354) );
  AND U531 ( .A(p_input[9842]), .B(p_input[39842]), .Z(n353) );
  AND U532 ( .A(n355), .B(n356), .Z(o[9841]) );
  AND U533 ( .A(p_input[29841]), .B(p_input[19841]), .Z(n356) );
  AND U534 ( .A(p_input[9841]), .B(p_input[39841]), .Z(n355) );
  AND U535 ( .A(n357), .B(n358), .Z(o[9840]) );
  AND U536 ( .A(p_input[29840]), .B(p_input[19840]), .Z(n358) );
  AND U537 ( .A(p_input[9840]), .B(p_input[39840]), .Z(n357) );
  AND U538 ( .A(n359), .B(n360), .Z(o[983]) );
  AND U539 ( .A(p_input[20983]), .B(p_input[10983]), .Z(n360) );
  AND U540 ( .A(p_input[983]), .B(p_input[30983]), .Z(n359) );
  AND U541 ( .A(n361), .B(n362), .Z(o[9839]) );
  AND U542 ( .A(p_input[29839]), .B(p_input[19839]), .Z(n362) );
  AND U543 ( .A(p_input[9839]), .B(p_input[39839]), .Z(n361) );
  AND U544 ( .A(n363), .B(n364), .Z(o[9838]) );
  AND U545 ( .A(p_input[29838]), .B(p_input[19838]), .Z(n364) );
  AND U546 ( .A(p_input[9838]), .B(p_input[39838]), .Z(n363) );
  AND U547 ( .A(n365), .B(n366), .Z(o[9837]) );
  AND U548 ( .A(p_input[29837]), .B(p_input[19837]), .Z(n366) );
  AND U549 ( .A(p_input[9837]), .B(p_input[39837]), .Z(n365) );
  AND U550 ( .A(n367), .B(n368), .Z(o[9836]) );
  AND U551 ( .A(p_input[29836]), .B(p_input[19836]), .Z(n368) );
  AND U552 ( .A(p_input[9836]), .B(p_input[39836]), .Z(n367) );
  AND U553 ( .A(n369), .B(n370), .Z(o[9835]) );
  AND U554 ( .A(p_input[29835]), .B(p_input[19835]), .Z(n370) );
  AND U555 ( .A(p_input[9835]), .B(p_input[39835]), .Z(n369) );
  AND U556 ( .A(n371), .B(n372), .Z(o[9834]) );
  AND U557 ( .A(p_input[29834]), .B(p_input[19834]), .Z(n372) );
  AND U558 ( .A(p_input[9834]), .B(p_input[39834]), .Z(n371) );
  AND U559 ( .A(n373), .B(n374), .Z(o[9833]) );
  AND U560 ( .A(p_input[29833]), .B(p_input[19833]), .Z(n374) );
  AND U561 ( .A(p_input[9833]), .B(p_input[39833]), .Z(n373) );
  AND U562 ( .A(n375), .B(n376), .Z(o[9832]) );
  AND U563 ( .A(p_input[29832]), .B(p_input[19832]), .Z(n376) );
  AND U564 ( .A(p_input[9832]), .B(p_input[39832]), .Z(n375) );
  AND U565 ( .A(n377), .B(n378), .Z(o[9831]) );
  AND U566 ( .A(p_input[29831]), .B(p_input[19831]), .Z(n378) );
  AND U567 ( .A(p_input[9831]), .B(p_input[39831]), .Z(n377) );
  AND U568 ( .A(n379), .B(n380), .Z(o[9830]) );
  AND U569 ( .A(p_input[29830]), .B(p_input[19830]), .Z(n380) );
  AND U570 ( .A(p_input[9830]), .B(p_input[39830]), .Z(n379) );
  AND U571 ( .A(n381), .B(n382), .Z(o[982]) );
  AND U572 ( .A(p_input[20982]), .B(p_input[10982]), .Z(n382) );
  AND U573 ( .A(p_input[982]), .B(p_input[30982]), .Z(n381) );
  AND U574 ( .A(n383), .B(n384), .Z(o[9829]) );
  AND U575 ( .A(p_input[29829]), .B(p_input[19829]), .Z(n384) );
  AND U576 ( .A(p_input[9829]), .B(p_input[39829]), .Z(n383) );
  AND U577 ( .A(n385), .B(n386), .Z(o[9828]) );
  AND U578 ( .A(p_input[29828]), .B(p_input[19828]), .Z(n386) );
  AND U579 ( .A(p_input[9828]), .B(p_input[39828]), .Z(n385) );
  AND U580 ( .A(n387), .B(n388), .Z(o[9827]) );
  AND U581 ( .A(p_input[29827]), .B(p_input[19827]), .Z(n388) );
  AND U582 ( .A(p_input[9827]), .B(p_input[39827]), .Z(n387) );
  AND U583 ( .A(n389), .B(n390), .Z(o[9826]) );
  AND U584 ( .A(p_input[29826]), .B(p_input[19826]), .Z(n390) );
  AND U585 ( .A(p_input[9826]), .B(p_input[39826]), .Z(n389) );
  AND U586 ( .A(n391), .B(n392), .Z(o[9825]) );
  AND U587 ( .A(p_input[29825]), .B(p_input[19825]), .Z(n392) );
  AND U588 ( .A(p_input[9825]), .B(p_input[39825]), .Z(n391) );
  AND U589 ( .A(n393), .B(n394), .Z(o[9824]) );
  AND U590 ( .A(p_input[29824]), .B(p_input[19824]), .Z(n394) );
  AND U591 ( .A(p_input[9824]), .B(p_input[39824]), .Z(n393) );
  AND U592 ( .A(n395), .B(n396), .Z(o[9823]) );
  AND U593 ( .A(p_input[29823]), .B(p_input[19823]), .Z(n396) );
  AND U594 ( .A(p_input[9823]), .B(p_input[39823]), .Z(n395) );
  AND U595 ( .A(n397), .B(n398), .Z(o[9822]) );
  AND U596 ( .A(p_input[29822]), .B(p_input[19822]), .Z(n398) );
  AND U597 ( .A(p_input[9822]), .B(p_input[39822]), .Z(n397) );
  AND U598 ( .A(n399), .B(n400), .Z(o[9821]) );
  AND U599 ( .A(p_input[29821]), .B(p_input[19821]), .Z(n400) );
  AND U600 ( .A(p_input[9821]), .B(p_input[39821]), .Z(n399) );
  AND U601 ( .A(n401), .B(n402), .Z(o[9820]) );
  AND U602 ( .A(p_input[29820]), .B(p_input[19820]), .Z(n402) );
  AND U603 ( .A(p_input[9820]), .B(p_input[39820]), .Z(n401) );
  AND U604 ( .A(n403), .B(n404), .Z(o[981]) );
  AND U605 ( .A(p_input[20981]), .B(p_input[10981]), .Z(n404) );
  AND U606 ( .A(p_input[981]), .B(p_input[30981]), .Z(n403) );
  AND U607 ( .A(n405), .B(n406), .Z(o[9819]) );
  AND U608 ( .A(p_input[29819]), .B(p_input[19819]), .Z(n406) );
  AND U609 ( .A(p_input[9819]), .B(p_input[39819]), .Z(n405) );
  AND U610 ( .A(n407), .B(n408), .Z(o[9818]) );
  AND U611 ( .A(p_input[29818]), .B(p_input[19818]), .Z(n408) );
  AND U612 ( .A(p_input[9818]), .B(p_input[39818]), .Z(n407) );
  AND U613 ( .A(n409), .B(n410), .Z(o[9817]) );
  AND U614 ( .A(p_input[29817]), .B(p_input[19817]), .Z(n410) );
  AND U615 ( .A(p_input[9817]), .B(p_input[39817]), .Z(n409) );
  AND U616 ( .A(n411), .B(n412), .Z(o[9816]) );
  AND U617 ( .A(p_input[29816]), .B(p_input[19816]), .Z(n412) );
  AND U618 ( .A(p_input[9816]), .B(p_input[39816]), .Z(n411) );
  AND U619 ( .A(n413), .B(n414), .Z(o[9815]) );
  AND U620 ( .A(p_input[29815]), .B(p_input[19815]), .Z(n414) );
  AND U621 ( .A(p_input[9815]), .B(p_input[39815]), .Z(n413) );
  AND U622 ( .A(n415), .B(n416), .Z(o[9814]) );
  AND U623 ( .A(p_input[29814]), .B(p_input[19814]), .Z(n416) );
  AND U624 ( .A(p_input[9814]), .B(p_input[39814]), .Z(n415) );
  AND U625 ( .A(n417), .B(n418), .Z(o[9813]) );
  AND U626 ( .A(p_input[29813]), .B(p_input[19813]), .Z(n418) );
  AND U627 ( .A(p_input[9813]), .B(p_input[39813]), .Z(n417) );
  AND U628 ( .A(n419), .B(n420), .Z(o[9812]) );
  AND U629 ( .A(p_input[29812]), .B(p_input[19812]), .Z(n420) );
  AND U630 ( .A(p_input[9812]), .B(p_input[39812]), .Z(n419) );
  AND U631 ( .A(n421), .B(n422), .Z(o[9811]) );
  AND U632 ( .A(p_input[29811]), .B(p_input[19811]), .Z(n422) );
  AND U633 ( .A(p_input[9811]), .B(p_input[39811]), .Z(n421) );
  AND U634 ( .A(n423), .B(n424), .Z(o[9810]) );
  AND U635 ( .A(p_input[29810]), .B(p_input[19810]), .Z(n424) );
  AND U636 ( .A(p_input[9810]), .B(p_input[39810]), .Z(n423) );
  AND U637 ( .A(n425), .B(n426), .Z(o[980]) );
  AND U638 ( .A(p_input[20980]), .B(p_input[10980]), .Z(n426) );
  AND U639 ( .A(p_input[980]), .B(p_input[30980]), .Z(n425) );
  AND U640 ( .A(n427), .B(n428), .Z(o[9809]) );
  AND U641 ( .A(p_input[29809]), .B(p_input[19809]), .Z(n428) );
  AND U642 ( .A(p_input[9809]), .B(p_input[39809]), .Z(n427) );
  AND U643 ( .A(n429), .B(n430), .Z(o[9808]) );
  AND U644 ( .A(p_input[29808]), .B(p_input[19808]), .Z(n430) );
  AND U645 ( .A(p_input[9808]), .B(p_input[39808]), .Z(n429) );
  AND U646 ( .A(n431), .B(n432), .Z(o[9807]) );
  AND U647 ( .A(p_input[29807]), .B(p_input[19807]), .Z(n432) );
  AND U648 ( .A(p_input[9807]), .B(p_input[39807]), .Z(n431) );
  AND U649 ( .A(n433), .B(n434), .Z(o[9806]) );
  AND U650 ( .A(p_input[29806]), .B(p_input[19806]), .Z(n434) );
  AND U651 ( .A(p_input[9806]), .B(p_input[39806]), .Z(n433) );
  AND U652 ( .A(n435), .B(n436), .Z(o[9805]) );
  AND U653 ( .A(p_input[29805]), .B(p_input[19805]), .Z(n436) );
  AND U654 ( .A(p_input[9805]), .B(p_input[39805]), .Z(n435) );
  AND U655 ( .A(n437), .B(n438), .Z(o[9804]) );
  AND U656 ( .A(p_input[29804]), .B(p_input[19804]), .Z(n438) );
  AND U657 ( .A(p_input[9804]), .B(p_input[39804]), .Z(n437) );
  AND U658 ( .A(n439), .B(n440), .Z(o[9803]) );
  AND U659 ( .A(p_input[29803]), .B(p_input[19803]), .Z(n440) );
  AND U660 ( .A(p_input[9803]), .B(p_input[39803]), .Z(n439) );
  AND U661 ( .A(n441), .B(n442), .Z(o[9802]) );
  AND U662 ( .A(p_input[29802]), .B(p_input[19802]), .Z(n442) );
  AND U663 ( .A(p_input[9802]), .B(p_input[39802]), .Z(n441) );
  AND U664 ( .A(n443), .B(n444), .Z(o[9801]) );
  AND U665 ( .A(p_input[29801]), .B(p_input[19801]), .Z(n444) );
  AND U666 ( .A(p_input[9801]), .B(p_input[39801]), .Z(n443) );
  AND U667 ( .A(n445), .B(n446), .Z(o[9800]) );
  AND U668 ( .A(p_input[29800]), .B(p_input[19800]), .Z(n446) );
  AND U669 ( .A(p_input[9800]), .B(p_input[39800]), .Z(n445) );
  AND U670 ( .A(n447), .B(n448), .Z(o[97]) );
  AND U671 ( .A(p_input[20097]), .B(p_input[10097]), .Z(n448) );
  AND U672 ( .A(p_input[97]), .B(p_input[30097]), .Z(n447) );
  AND U673 ( .A(n449), .B(n450), .Z(o[979]) );
  AND U674 ( .A(p_input[20979]), .B(p_input[10979]), .Z(n450) );
  AND U675 ( .A(p_input[979]), .B(p_input[30979]), .Z(n449) );
  AND U676 ( .A(n451), .B(n452), .Z(o[9799]) );
  AND U677 ( .A(p_input[29799]), .B(p_input[19799]), .Z(n452) );
  AND U678 ( .A(p_input[9799]), .B(p_input[39799]), .Z(n451) );
  AND U679 ( .A(n453), .B(n454), .Z(o[9798]) );
  AND U680 ( .A(p_input[29798]), .B(p_input[19798]), .Z(n454) );
  AND U681 ( .A(p_input[9798]), .B(p_input[39798]), .Z(n453) );
  AND U682 ( .A(n455), .B(n456), .Z(o[9797]) );
  AND U683 ( .A(p_input[29797]), .B(p_input[19797]), .Z(n456) );
  AND U684 ( .A(p_input[9797]), .B(p_input[39797]), .Z(n455) );
  AND U685 ( .A(n457), .B(n458), .Z(o[9796]) );
  AND U686 ( .A(p_input[29796]), .B(p_input[19796]), .Z(n458) );
  AND U687 ( .A(p_input[9796]), .B(p_input[39796]), .Z(n457) );
  AND U688 ( .A(n459), .B(n460), .Z(o[9795]) );
  AND U689 ( .A(p_input[29795]), .B(p_input[19795]), .Z(n460) );
  AND U690 ( .A(p_input[9795]), .B(p_input[39795]), .Z(n459) );
  AND U691 ( .A(n461), .B(n462), .Z(o[9794]) );
  AND U692 ( .A(p_input[29794]), .B(p_input[19794]), .Z(n462) );
  AND U693 ( .A(p_input[9794]), .B(p_input[39794]), .Z(n461) );
  AND U694 ( .A(n463), .B(n464), .Z(o[9793]) );
  AND U695 ( .A(p_input[29793]), .B(p_input[19793]), .Z(n464) );
  AND U696 ( .A(p_input[9793]), .B(p_input[39793]), .Z(n463) );
  AND U697 ( .A(n465), .B(n466), .Z(o[9792]) );
  AND U698 ( .A(p_input[29792]), .B(p_input[19792]), .Z(n466) );
  AND U699 ( .A(p_input[9792]), .B(p_input[39792]), .Z(n465) );
  AND U700 ( .A(n467), .B(n468), .Z(o[9791]) );
  AND U701 ( .A(p_input[29791]), .B(p_input[19791]), .Z(n468) );
  AND U702 ( .A(p_input[9791]), .B(p_input[39791]), .Z(n467) );
  AND U703 ( .A(n469), .B(n470), .Z(o[9790]) );
  AND U704 ( .A(p_input[29790]), .B(p_input[19790]), .Z(n470) );
  AND U705 ( .A(p_input[9790]), .B(p_input[39790]), .Z(n469) );
  AND U706 ( .A(n471), .B(n472), .Z(o[978]) );
  AND U707 ( .A(p_input[20978]), .B(p_input[10978]), .Z(n472) );
  AND U708 ( .A(p_input[978]), .B(p_input[30978]), .Z(n471) );
  AND U709 ( .A(n473), .B(n474), .Z(o[9789]) );
  AND U710 ( .A(p_input[29789]), .B(p_input[19789]), .Z(n474) );
  AND U711 ( .A(p_input[9789]), .B(p_input[39789]), .Z(n473) );
  AND U712 ( .A(n475), .B(n476), .Z(o[9788]) );
  AND U713 ( .A(p_input[29788]), .B(p_input[19788]), .Z(n476) );
  AND U714 ( .A(p_input[9788]), .B(p_input[39788]), .Z(n475) );
  AND U715 ( .A(n477), .B(n478), .Z(o[9787]) );
  AND U716 ( .A(p_input[29787]), .B(p_input[19787]), .Z(n478) );
  AND U717 ( .A(p_input[9787]), .B(p_input[39787]), .Z(n477) );
  AND U718 ( .A(n479), .B(n480), .Z(o[9786]) );
  AND U719 ( .A(p_input[29786]), .B(p_input[19786]), .Z(n480) );
  AND U720 ( .A(p_input[9786]), .B(p_input[39786]), .Z(n479) );
  AND U721 ( .A(n481), .B(n482), .Z(o[9785]) );
  AND U722 ( .A(p_input[29785]), .B(p_input[19785]), .Z(n482) );
  AND U723 ( .A(p_input[9785]), .B(p_input[39785]), .Z(n481) );
  AND U724 ( .A(n483), .B(n484), .Z(o[9784]) );
  AND U725 ( .A(p_input[29784]), .B(p_input[19784]), .Z(n484) );
  AND U726 ( .A(p_input[9784]), .B(p_input[39784]), .Z(n483) );
  AND U727 ( .A(n485), .B(n486), .Z(o[9783]) );
  AND U728 ( .A(p_input[29783]), .B(p_input[19783]), .Z(n486) );
  AND U729 ( .A(p_input[9783]), .B(p_input[39783]), .Z(n485) );
  AND U730 ( .A(n487), .B(n488), .Z(o[9782]) );
  AND U731 ( .A(p_input[29782]), .B(p_input[19782]), .Z(n488) );
  AND U732 ( .A(p_input[9782]), .B(p_input[39782]), .Z(n487) );
  AND U733 ( .A(n489), .B(n490), .Z(o[9781]) );
  AND U734 ( .A(p_input[29781]), .B(p_input[19781]), .Z(n490) );
  AND U735 ( .A(p_input[9781]), .B(p_input[39781]), .Z(n489) );
  AND U736 ( .A(n491), .B(n492), .Z(o[9780]) );
  AND U737 ( .A(p_input[29780]), .B(p_input[19780]), .Z(n492) );
  AND U738 ( .A(p_input[9780]), .B(p_input[39780]), .Z(n491) );
  AND U739 ( .A(n493), .B(n494), .Z(o[977]) );
  AND U740 ( .A(p_input[20977]), .B(p_input[10977]), .Z(n494) );
  AND U741 ( .A(p_input[977]), .B(p_input[30977]), .Z(n493) );
  AND U742 ( .A(n495), .B(n496), .Z(o[9779]) );
  AND U743 ( .A(p_input[29779]), .B(p_input[19779]), .Z(n496) );
  AND U744 ( .A(p_input[9779]), .B(p_input[39779]), .Z(n495) );
  AND U745 ( .A(n497), .B(n498), .Z(o[9778]) );
  AND U746 ( .A(p_input[29778]), .B(p_input[19778]), .Z(n498) );
  AND U747 ( .A(p_input[9778]), .B(p_input[39778]), .Z(n497) );
  AND U748 ( .A(n499), .B(n500), .Z(o[9777]) );
  AND U749 ( .A(p_input[29777]), .B(p_input[19777]), .Z(n500) );
  AND U750 ( .A(p_input[9777]), .B(p_input[39777]), .Z(n499) );
  AND U751 ( .A(n501), .B(n502), .Z(o[9776]) );
  AND U752 ( .A(p_input[29776]), .B(p_input[19776]), .Z(n502) );
  AND U753 ( .A(p_input[9776]), .B(p_input[39776]), .Z(n501) );
  AND U754 ( .A(n503), .B(n504), .Z(o[9775]) );
  AND U755 ( .A(p_input[29775]), .B(p_input[19775]), .Z(n504) );
  AND U756 ( .A(p_input[9775]), .B(p_input[39775]), .Z(n503) );
  AND U757 ( .A(n505), .B(n506), .Z(o[9774]) );
  AND U758 ( .A(p_input[29774]), .B(p_input[19774]), .Z(n506) );
  AND U759 ( .A(p_input[9774]), .B(p_input[39774]), .Z(n505) );
  AND U760 ( .A(n507), .B(n508), .Z(o[9773]) );
  AND U761 ( .A(p_input[29773]), .B(p_input[19773]), .Z(n508) );
  AND U762 ( .A(p_input[9773]), .B(p_input[39773]), .Z(n507) );
  AND U763 ( .A(n509), .B(n510), .Z(o[9772]) );
  AND U764 ( .A(p_input[29772]), .B(p_input[19772]), .Z(n510) );
  AND U765 ( .A(p_input[9772]), .B(p_input[39772]), .Z(n509) );
  AND U766 ( .A(n511), .B(n512), .Z(o[9771]) );
  AND U767 ( .A(p_input[29771]), .B(p_input[19771]), .Z(n512) );
  AND U768 ( .A(p_input[9771]), .B(p_input[39771]), .Z(n511) );
  AND U769 ( .A(n513), .B(n514), .Z(o[9770]) );
  AND U770 ( .A(p_input[29770]), .B(p_input[19770]), .Z(n514) );
  AND U771 ( .A(p_input[9770]), .B(p_input[39770]), .Z(n513) );
  AND U772 ( .A(n515), .B(n516), .Z(o[976]) );
  AND U773 ( .A(p_input[20976]), .B(p_input[10976]), .Z(n516) );
  AND U774 ( .A(p_input[976]), .B(p_input[30976]), .Z(n515) );
  AND U775 ( .A(n517), .B(n518), .Z(o[9769]) );
  AND U776 ( .A(p_input[29769]), .B(p_input[19769]), .Z(n518) );
  AND U777 ( .A(p_input[9769]), .B(p_input[39769]), .Z(n517) );
  AND U778 ( .A(n519), .B(n520), .Z(o[9768]) );
  AND U779 ( .A(p_input[29768]), .B(p_input[19768]), .Z(n520) );
  AND U780 ( .A(p_input[9768]), .B(p_input[39768]), .Z(n519) );
  AND U781 ( .A(n521), .B(n522), .Z(o[9767]) );
  AND U782 ( .A(p_input[29767]), .B(p_input[19767]), .Z(n522) );
  AND U783 ( .A(p_input[9767]), .B(p_input[39767]), .Z(n521) );
  AND U784 ( .A(n523), .B(n524), .Z(o[9766]) );
  AND U785 ( .A(p_input[29766]), .B(p_input[19766]), .Z(n524) );
  AND U786 ( .A(p_input[9766]), .B(p_input[39766]), .Z(n523) );
  AND U787 ( .A(n525), .B(n526), .Z(o[9765]) );
  AND U788 ( .A(p_input[29765]), .B(p_input[19765]), .Z(n526) );
  AND U789 ( .A(p_input[9765]), .B(p_input[39765]), .Z(n525) );
  AND U790 ( .A(n527), .B(n528), .Z(o[9764]) );
  AND U791 ( .A(p_input[29764]), .B(p_input[19764]), .Z(n528) );
  AND U792 ( .A(p_input[9764]), .B(p_input[39764]), .Z(n527) );
  AND U793 ( .A(n529), .B(n530), .Z(o[9763]) );
  AND U794 ( .A(p_input[29763]), .B(p_input[19763]), .Z(n530) );
  AND U795 ( .A(p_input[9763]), .B(p_input[39763]), .Z(n529) );
  AND U796 ( .A(n531), .B(n532), .Z(o[9762]) );
  AND U797 ( .A(p_input[29762]), .B(p_input[19762]), .Z(n532) );
  AND U798 ( .A(p_input[9762]), .B(p_input[39762]), .Z(n531) );
  AND U799 ( .A(n533), .B(n534), .Z(o[9761]) );
  AND U800 ( .A(p_input[29761]), .B(p_input[19761]), .Z(n534) );
  AND U801 ( .A(p_input[9761]), .B(p_input[39761]), .Z(n533) );
  AND U802 ( .A(n535), .B(n536), .Z(o[9760]) );
  AND U803 ( .A(p_input[29760]), .B(p_input[19760]), .Z(n536) );
  AND U804 ( .A(p_input[9760]), .B(p_input[39760]), .Z(n535) );
  AND U805 ( .A(n537), .B(n538), .Z(o[975]) );
  AND U806 ( .A(p_input[20975]), .B(p_input[10975]), .Z(n538) );
  AND U807 ( .A(p_input[975]), .B(p_input[30975]), .Z(n537) );
  AND U808 ( .A(n539), .B(n540), .Z(o[9759]) );
  AND U809 ( .A(p_input[29759]), .B(p_input[19759]), .Z(n540) );
  AND U810 ( .A(p_input[9759]), .B(p_input[39759]), .Z(n539) );
  AND U811 ( .A(n541), .B(n542), .Z(o[9758]) );
  AND U812 ( .A(p_input[29758]), .B(p_input[19758]), .Z(n542) );
  AND U813 ( .A(p_input[9758]), .B(p_input[39758]), .Z(n541) );
  AND U814 ( .A(n543), .B(n544), .Z(o[9757]) );
  AND U815 ( .A(p_input[29757]), .B(p_input[19757]), .Z(n544) );
  AND U816 ( .A(p_input[9757]), .B(p_input[39757]), .Z(n543) );
  AND U817 ( .A(n545), .B(n546), .Z(o[9756]) );
  AND U818 ( .A(p_input[29756]), .B(p_input[19756]), .Z(n546) );
  AND U819 ( .A(p_input[9756]), .B(p_input[39756]), .Z(n545) );
  AND U820 ( .A(n547), .B(n548), .Z(o[9755]) );
  AND U821 ( .A(p_input[29755]), .B(p_input[19755]), .Z(n548) );
  AND U822 ( .A(p_input[9755]), .B(p_input[39755]), .Z(n547) );
  AND U823 ( .A(n549), .B(n550), .Z(o[9754]) );
  AND U824 ( .A(p_input[29754]), .B(p_input[19754]), .Z(n550) );
  AND U825 ( .A(p_input[9754]), .B(p_input[39754]), .Z(n549) );
  AND U826 ( .A(n551), .B(n552), .Z(o[9753]) );
  AND U827 ( .A(p_input[29753]), .B(p_input[19753]), .Z(n552) );
  AND U828 ( .A(p_input[9753]), .B(p_input[39753]), .Z(n551) );
  AND U829 ( .A(n553), .B(n554), .Z(o[9752]) );
  AND U830 ( .A(p_input[29752]), .B(p_input[19752]), .Z(n554) );
  AND U831 ( .A(p_input[9752]), .B(p_input[39752]), .Z(n553) );
  AND U832 ( .A(n555), .B(n556), .Z(o[9751]) );
  AND U833 ( .A(p_input[29751]), .B(p_input[19751]), .Z(n556) );
  AND U834 ( .A(p_input[9751]), .B(p_input[39751]), .Z(n555) );
  AND U835 ( .A(n557), .B(n558), .Z(o[9750]) );
  AND U836 ( .A(p_input[29750]), .B(p_input[19750]), .Z(n558) );
  AND U837 ( .A(p_input[9750]), .B(p_input[39750]), .Z(n557) );
  AND U838 ( .A(n559), .B(n560), .Z(o[974]) );
  AND U839 ( .A(p_input[20974]), .B(p_input[10974]), .Z(n560) );
  AND U840 ( .A(p_input[974]), .B(p_input[30974]), .Z(n559) );
  AND U841 ( .A(n561), .B(n562), .Z(o[9749]) );
  AND U842 ( .A(p_input[29749]), .B(p_input[19749]), .Z(n562) );
  AND U843 ( .A(p_input[9749]), .B(p_input[39749]), .Z(n561) );
  AND U844 ( .A(n563), .B(n564), .Z(o[9748]) );
  AND U845 ( .A(p_input[29748]), .B(p_input[19748]), .Z(n564) );
  AND U846 ( .A(p_input[9748]), .B(p_input[39748]), .Z(n563) );
  AND U847 ( .A(n565), .B(n566), .Z(o[9747]) );
  AND U848 ( .A(p_input[29747]), .B(p_input[19747]), .Z(n566) );
  AND U849 ( .A(p_input[9747]), .B(p_input[39747]), .Z(n565) );
  AND U850 ( .A(n567), .B(n568), .Z(o[9746]) );
  AND U851 ( .A(p_input[29746]), .B(p_input[19746]), .Z(n568) );
  AND U852 ( .A(p_input[9746]), .B(p_input[39746]), .Z(n567) );
  AND U853 ( .A(n569), .B(n570), .Z(o[9745]) );
  AND U854 ( .A(p_input[29745]), .B(p_input[19745]), .Z(n570) );
  AND U855 ( .A(p_input[9745]), .B(p_input[39745]), .Z(n569) );
  AND U856 ( .A(n571), .B(n572), .Z(o[9744]) );
  AND U857 ( .A(p_input[29744]), .B(p_input[19744]), .Z(n572) );
  AND U858 ( .A(p_input[9744]), .B(p_input[39744]), .Z(n571) );
  AND U859 ( .A(n573), .B(n574), .Z(o[9743]) );
  AND U860 ( .A(p_input[29743]), .B(p_input[19743]), .Z(n574) );
  AND U861 ( .A(p_input[9743]), .B(p_input[39743]), .Z(n573) );
  AND U862 ( .A(n575), .B(n576), .Z(o[9742]) );
  AND U863 ( .A(p_input[29742]), .B(p_input[19742]), .Z(n576) );
  AND U864 ( .A(p_input[9742]), .B(p_input[39742]), .Z(n575) );
  AND U865 ( .A(n577), .B(n578), .Z(o[9741]) );
  AND U866 ( .A(p_input[29741]), .B(p_input[19741]), .Z(n578) );
  AND U867 ( .A(p_input[9741]), .B(p_input[39741]), .Z(n577) );
  AND U868 ( .A(n579), .B(n580), .Z(o[9740]) );
  AND U869 ( .A(p_input[29740]), .B(p_input[19740]), .Z(n580) );
  AND U870 ( .A(p_input[9740]), .B(p_input[39740]), .Z(n579) );
  AND U871 ( .A(n581), .B(n582), .Z(o[973]) );
  AND U872 ( .A(p_input[20973]), .B(p_input[10973]), .Z(n582) );
  AND U873 ( .A(p_input[973]), .B(p_input[30973]), .Z(n581) );
  AND U874 ( .A(n583), .B(n584), .Z(o[9739]) );
  AND U875 ( .A(p_input[29739]), .B(p_input[19739]), .Z(n584) );
  AND U876 ( .A(p_input[9739]), .B(p_input[39739]), .Z(n583) );
  AND U877 ( .A(n585), .B(n586), .Z(o[9738]) );
  AND U878 ( .A(p_input[29738]), .B(p_input[19738]), .Z(n586) );
  AND U879 ( .A(p_input[9738]), .B(p_input[39738]), .Z(n585) );
  AND U880 ( .A(n587), .B(n588), .Z(o[9737]) );
  AND U881 ( .A(p_input[29737]), .B(p_input[19737]), .Z(n588) );
  AND U882 ( .A(p_input[9737]), .B(p_input[39737]), .Z(n587) );
  AND U883 ( .A(n589), .B(n590), .Z(o[9736]) );
  AND U884 ( .A(p_input[29736]), .B(p_input[19736]), .Z(n590) );
  AND U885 ( .A(p_input[9736]), .B(p_input[39736]), .Z(n589) );
  AND U886 ( .A(n591), .B(n592), .Z(o[9735]) );
  AND U887 ( .A(p_input[29735]), .B(p_input[19735]), .Z(n592) );
  AND U888 ( .A(p_input[9735]), .B(p_input[39735]), .Z(n591) );
  AND U889 ( .A(n593), .B(n594), .Z(o[9734]) );
  AND U890 ( .A(p_input[29734]), .B(p_input[19734]), .Z(n594) );
  AND U891 ( .A(p_input[9734]), .B(p_input[39734]), .Z(n593) );
  AND U892 ( .A(n595), .B(n596), .Z(o[9733]) );
  AND U893 ( .A(p_input[29733]), .B(p_input[19733]), .Z(n596) );
  AND U894 ( .A(p_input[9733]), .B(p_input[39733]), .Z(n595) );
  AND U895 ( .A(n597), .B(n598), .Z(o[9732]) );
  AND U896 ( .A(p_input[29732]), .B(p_input[19732]), .Z(n598) );
  AND U897 ( .A(p_input[9732]), .B(p_input[39732]), .Z(n597) );
  AND U898 ( .A(n599), .B(n600), .Z(o[9731]) );
  AND U899 ( .A(p_input[29731]), .B(p_input[19731]), .Z(n600) );
  AND U900 ( .A(p_input[9731]), .B(p_input[39731]), .Z(n599) );
  AND U901 ( .A(n601), .B(n602), .Z(o[9730]) );
  AND U902 ( .A(p_input[29730]), .B(p_input[19730]), .Z(n602) );
  AND U903 ( .A(p_input[9730]), .B(p_input[39730]), .Z(n601) );
  AND U904 ( .A(n603), .B(n604), .Z(o[972]) );
  AND U905 ( .A(p_input[20972]), .B(p_input[10972]), .Z(n604) );
  AND U906 ( .A(p_input[972]), .B(p_input[30972]), .Z(n603) );
  AND U907 ( .A(n605), .B(n606), .Z(o[9729]) );
  AND U908 ( .A(p_input[29729]), .B(p_input[19729]), .Z(n606) );
  AND U909 ( .A(p_input[9729]), .B(p_input[39729]), .Z(n605) );
  AND U910 ( .A(n607), .B(n608), .Z(o[9728]) );
  AND U911 ( .A(p_input[29728]), .B(p_input[19728]), .Z(n608) );
  AND U912 ( .A(p_input[9728]), .B(p_input[39728]), .Z(n607) );
  AND U913 ( .A(n609), .B(n610), .Z(o[9727]) );
  AND U914 ( .A(p_input[29727]), .B(p_input[19727]), .Z(n610) );
  AND U915 ( .A(p_input[9727]), .B(p_input[39727]), .Z(n609) );
  AND U916 ( .A(n611), .B(n612), .Z(o[9726]) );
  AND U917 ( .A(p_input[29726]), .B(p_input[19726]), .Z(n612) );
  AND U918 ( .A(p_input[9726]), .B(p_input[39726]), .Z(n611) );
  AND U919 ( .A(n613), .B(n614), .Z(o[9725]) );
  AND U920 ( .A(p_input[29725]), .B(p_input[19725]), .Z(n614) );
  AND U921 ( .A(p_input[9725]), .B(p_input[39725]), .Z(n613) );
  AND U922 ( .A(n615), .B(n616), .Z(o[9724]) );
  AND U923 ( .A(p_input[29724]), .B(p_input[19724]), .Z(n616) );
  AND U924 ( .A(p_input[9724]), .B(p_input[39724]), .Z(n615) );
  AND U925 ( .A(n617), .B(n618), .Z(o[9723]) );
  AND U926 ( .A(p_input[29723]), .B(p_input[19723]), .Z(n618) );
  AND U927 ( .A(p_input[9723]), .B(p_input[39723]), .Z(n617) );
  AND U928 ( .A(n619), .B(n620), .Z(o[9722]) );
  AND U929 ( .A(p_input[29722]), .B(p_input[19722]), .Z(n620) );
  AND U930 ( .A(p_input[9722]), .B(p_input[39722]), .Z(n619) );
  AND U931 ( .A(n621), .B(n622), .Z(o[9721]) );
  AND U932 ( .A(p_input[29721]), .B(p_input[19721]), .Z(n622) );
  AND U933 ( .A(p_input[9721]), .B(p_input[39721]), .Z(n621) );
  AND U934 ( .A(n623), .B(n624), .Z(o[9720]) );
  AND U935 ( .A(p_input[29720]), .B(p_input[19720]), .Z(n624) );
  AND U936 ( .A(p_input[9720]), .B(p_input[39720]), .Z(n623) );
  AND U937 ( .A(n625), .B(n626), .Z(o[971]) );
  AND U938 ( .A(p_input[20971]), .B(p_input[10971]), .Z(n626) );
  AND U939 ( .A(p_input[971]), .B(p_input[30971]), .Z(n625) );
  AND U940 ( .A(n627), .B(n628), .Z(o[9719]) );
  AND U941 ( .A(p_input[29719]), .B(p_input[19719]), .Z(n628) );
  AND U942 ( .A(p_input[9719]), .B(p_input[39719]), .Z(n627) );
  AND U943 ( .A(n629), .B(n630), .Z(o[9718]) );
  AND U944 ( .A(p_input[29718]), .B(p_input[19718]), .Z(n630) );
  AND U945 ( .A(p_input[9718]), .B(p_input[39718]), .Z(n629) );
  AND U946 ( .A(n631), .B(n632), .Z(o[9717]) );
  AND U947 ( .A(p_input[29717]), .B(p_input[19717]), .Z(n632) );
  AND U948 ( .A(p_input[9717]), .B(p_input[39717]), .Z(n631) );
  AND U949 ( .A(n633), .B(n634), .Z(o[9716]) );
  AND U950 ( .A(p_input[29716]), .B(p_input[19716]), .Z(n634) );
  AND U951 ( .A(p_input[9716]), .B(p_input[39716]), .Z(n633) );
  AND U952 ( .A(n635), .B(n636), .Z(o[9715]) );
  AND U953 ( .A(p_input[29715]), .B(p_input[19715]), .Z(n636) );
  AND U954 ( .A(p_input[9715]), .B(p_input[39715]), .Z(n635) );
  AND U955 ( .A(n637), .B(n638), .Z(o[9714]) );
  AND U956 ( .A(p_input[29714]), .B(p_input[19714]), .Z(n638) );
  AND U957 ( .A(p_input[9714]), .B(p_input[39714]), .Z(n637) );
  AND U958 ( .A(n639), .B(n640), .Z(o[9713]) );
  AND U959 ( .A(p_input[29713]), .B(p_input[19713]), .Z(n640) );
  AND U960 ( .A(p_input[9713]), .B(p_input[39713]), .Z(n639) );
  AND U961 ( .A(n641), .B(n642), .Z(o[9712]) );
  AND U962 ( .A(p_input[29712]), .B(p_input[19712]), .Z(n642) );
  AND U963 ( .A(p_input[9712]), .B(p_input[39712]), .Z(n641) );
  AND U964 ( .A(n643), .B(n644), .Z(o[9711]) );
  AND U965 ( .A(p_input[29711]), .B(p_input[19711]), .Z(n644) );
  AND U966 ( .A(p_input[9711]), .B(p_input[39711]), .Z(n643) );
  AND U967 ( .A(n645), .B(n646), .Z(o[9710]) );
  AND U968 ( .A(p_input[29710]), .B(p_input[19710]), .Z(n646) );
  AND U969 ( .A(p_input[9710]), .B(p_input[39710]), .Z(n645) );
  AND U970 ( .A(n647), .B(n648), .Z(o[970]) );
  AND U971 ( .A(p_input[20970]), .B(p_input[10970]), .Z(n648) );
  AND U972 ( .A(p_input[970]), .B(p_input[30970]), .Z(n647) );
  AND U973 ( .A(n649), .B(n650), .Z(o[9709]) );
  AND U974 ( .A(p_input[29709]), .B(p_input[19709]), .Z(n650) );
  AND U975 ( .A(p_input[9709]), .B(p_input[39709]), .Z(n649) );
  AND U976 ( .A(n651), .B(n652), .Z(o[9708]) );
  AND U977 ( .A(p_input[29708]), .B(p_input[19708]), .Z(n652) );
  AND U978 ( .A(p_input[9708]), .B(p_input[39708]), .Z(n651) );
  AND U979 ( .A(n653), .B(n654), .Z(o[9707]) );
  AND U980 ( .A(p_input[29707]), .B(p_input[19707]), .Z(n654) );
  AND U981 ( .A(p_input[9707]), .B(p_input[39707]), .Z(n653) );
  AND U982 ( .A(n655), .B(n656), .Z(o[9706]) );
  AND U983 ( .A(p_input[29706]), .B(p_input[19706]), .Z(n656) );
  AND U984 ( .A(p_input[9706]), .B(p_input[39706]), .Z(n655) );
  AND U985 ( .A(n657), .B(n658), .Z(o[9705]) );
  AND U986 ( .A(p_input[29705]), .B(p_input[19705]), .Z(n658) );
  AND U987 ( .A(p_input[9705]), .B(p_input[39705]), .Z(n657) );
  AND U988 ( .A(n659), .B(n660), .Z(o[9704]) );
  AND U989 ( .A(p_input[29704]), .B(p_input[19704]), .Z(n660) );
  AND U990 ( .A(p_input[9704]), .B(p_input[39704]), .Z(n659) );
  AND U991 ( .A(n661), .B(n662), .Z(o[9703]) );
  AND U992 ( .A(p_input[29703]), .B(p_input[19703]), .Z(n662) );
  AND U993 ( .A(p_input[9703]), .B(p_input[39703]), .Z(n661) );
  AND U994 ( .A(n663), .B(n664), .Z(o[9702]) );
  AND U995 ( .A(p_input[29702]), .B(p_input[19702]), .Z(n664) );
  AND U996 ( .A(p_input[9702]), .B(p_input[39702]), .Z(n663) );
  AND U997 ( .A(n665), .B(n666), .Z(o[9701]) );
  AND U998 ( .A(p_input[29701]), .B(p_input[19701]), .Z(n666) );
  AND U999 ( .A(p_input[9701]), .B(p_input[39701]), .Z(n665) );
  AND U1000 ( .A(n667), .B(n668), .Z(o[9700]) );
  AND U1001 ( .A(p_input[29700]), .B(p_input[19700]), .Z(n668) );
  AND U1002 ( .A(p_input[9700]), .B(p_input[39700]), .Z(n667) );
  AND U1003 ( .A(n669), .B(n670), .Z(o[96]) );
  AND U1004 ( .A(p_input[20096]), .B(p_input[10096]), .Z(n670) );
  AND U1005 ( .A(p_input[96]), .B(p_input[30096]), .Z(n669) );
  AND U1006 ( .A(n671), .B(n672), .Z(o[969]) );
  AND U1007 ( .A(p_input[20969]), .B(p_input[10969]), .Z(n672) );
  AND U1008 ( .A(p_input[969]), .B(p_input[30969]), .Z(n671) );
  AND U1009 ( .A(n673), .B(n674), .Z(o[9699]) );
  AND U1010 ( .A(p_input[29699]), .B(p_input[19699]), .Z(n674) );
  AND U1011 ( .A(p_input[9699]), .B(p_input[39699]), .Z(n673) );
  AND U1012 ( .A(n675), .B(n676), .Z(o[9698]) );
  AND U1013 ( .A(p_input[29698]), .B(p_input[19698]), .Z(n676) );
  AND U1014 ( .A(p_input[9698]), .B(p_input[39698]), .Z(n675) );
  AND U1015 ( .A(n677), .B(n678), .Z(o[9697]) );
  AND U1016 ( .A(p_input[29697]), .B(p_input[19697]), .Z(n678) );
  AND U1017 ( .A(p_input[9697]), .B(p_input[39697]), .Z(n677) );
  AND U1018 ( .A(n679), .B(n680), .Z(o[9696]) );
  AND U1019 ( .A(p_input[29696]), .B(p_input[19696]), .Z(n680) );
  AND U1020 ( .A(p_input[9696]), .B(p_input[39696]), .Z(n679) );
  AND U1021 ( .A(n681), .B(n682), .Z(o[9695]) );
  AND U1022 ( .A(p_input[29695]), .B(p_input[19695]), .Z(n682) );
  AND U1023 ( .A(p_input[9695]), .B(p_input[39695]), .Z(n681) );
  AND U1024 ( .A(n683), .B(n684), .Z(o[9694]) );
  AND U1025 ( .A(p_input[29694]), .B(p_input[19694]), .Z(n684) );
  AND U1026 ( .A(p_input[9694]), .B(p_input[39694]), .Z(n683) );
  AND U1027 ( .A(n685), .B(n686), .Z(o[9693]) );
  AND U1028 ( .A(p_input[29693]), .B(p_input[19693]), .Z(n686) );
  AND U1029 ( .A(p_input[9693]), .B(p_input[39693]), .Z(n685) );
  AND U1030 ( .A(n687), .B(n688), .Z(o[9692]) );
  AND U1031 ( .A(p_input[29692]), .B(p_input[19692]), .Z(n688) );
  AND U1032 ( .A(p_input[9692]), .B(p_input[39692]), .Z(n687) );
  AND U1033 ( .A(n689), .B(n690), .Z(o[9691]) );
  AND U1034 ( .A(p_input[29691]), .B(p_input[19691]), .Z(n690) );
  AND U1035 ( .A(p_input[9691]), .B(p_input[39691]), .Z(n689) );
  AND U1036 ( .A(n691), .B(n692), .Z(o[9690]) );
  AND U1037 ( .A(p_input[29690]), .B(p_input[19690]), .Z(n692) );
  AND U1038 ( .A(p_input[9690]), .B(p_input[39690]), .Z(n691) );
  AND U1039 ( .A(n693), .B(n694), .Z(o[968]) );
  AND U1040 ( .A(p_input[20968]), .B(p_input[10968]), .Z(n694) );
  AND U1041 ( .A(p_input[968]), .B(p_input[30968]), .Z(n693) );
  AND U1042 ( .A(n695), .B(n696), .Z(o[9689]) );
  AND U1043 ( .A(p_input[29689]), .B(p_input[19689]), .Z(n696) );
  AND U1044 ( .A(p_input[9689]), .B(p_input[39689]), .Z(n695) );
  AND U1045 ( .A(n697), .B(n698), .Z(o[9688]) );
  AND U1046 ( .A(p_input[29688]), .B(p_input[19688]), .Z(n698) );
  AND U1047 ( .A(p_input[9688]), .B(p_input[39688]), .Z(n697) );
  AND U1048 ( .A(n699), .B(n700), .Z(o[9687]) );
  AND U1049 ( .A(p_input[29687]), .B(p_input[19687]), .Z(n700) );
  AND U1050 ( .A(p_input[9687]), .B(p_input[39687]), .Z(n699) );
  AND U1051 ( .A(n701), .B(n702), .Z(o[9686]) );
  AND U1052 ( .A(p_input[29686]), .B(p_input[19686]), .Z(n702) );
  AND U1053 ( .A(p_input[9686]), .B(p_input[39686]), .Z(n701) );
  AND U1054 ( .A(n703), .B(n704), .Z(o[9685]) );
  AND U1055 ( .A(p_input[29685]), .B(p_input[19685]), .Z(n704) );
  AND U1056 ( .A(p_input[9685]), .B(p_input[39685]), .Z(n703) );
  AND U1057 ( .A(n705), .B(n706), .Z(o[9684]) );
  AND U1058 ( .A(p_input[29684]), .B(p_input[19684]), .Z(n706) );
  AND U1059 ( .A(p_input[9684]), .B(p_input[39684]), .Z(n705) );
  AND U1060 ( .A(n707), .B(n708), .Z(o[9683]) );
  AND U1061 ( .A(p_input[29683]), .B(p_input[19683]), .Z(n708) );
  AND U1062 ( .A(p_input[9683]), .B(p_input[39683]), .Z(n707) );
  AND U1063 ( .A(n709), .B(n710), .Z(o[9682]) );
  AND U1064 ( .A(p_input[29682]), .B(p_input[19682]), .Z(n710) );
  AND U1065 ( .A(p_input[9682]), .B(p_input[39682]), .Z(n709) );
  AND U1066 ( .A(n711), .B(n712), .Z(o[9681]) );
  AND U1067 ( .A(p_input[29681]), .B(p_input[19681]), .Z(n712) );
  AND U1068 ( .A(p_input[9681]), .B(p_input[39681]), .Z(n711) );
  AND U1069 ( .A(n713), .B(n714), .Z(o[9680]) );
  AND U1070 ( .A(p_input[29680]), .B(p_input[19680]), .Z(n714) );
  AND U1071 ( .A(p_input[9680]), .B(p_input[39680]), .Z(n713) );
  AND U1072 ( .A(n715), .B(n716), .Z(o[967]) );
  AND U1073 ( .A(p_input[20967]), .B(p_input[10967]), .Z(n716) );
  AND U1074 ( .A(p_input[967]), .B(p_input[30967]), .Z(n715) );
  AND U1075 ( .A(n717), .B(n718), .Z(o[9679]) );
  AND U1076 ( .A(p_input[29679]), .B(p_input[19679]), .Z(n718) );
  AND U1077 ( .A(p_input[9679]), .B(p_input[39679]), .Z(n717) );
  AND U1078 ( .A(n719), .B(n720), .Z(o[9678]) );
  AND U1079 ( .A(p_input[29678]), .B(p_input[19678]), .Z(n720) );
  AND U1080 ( .A(p_input[9678]), .B(p_input[39678]), .Z(n719) );
  AND U1081 ( .A(n721), .B(n722), .Z(o[9677]) );
  AND U1082 ( .A(p_input[29677]), .B(p_input[19677]), .Z(n722) );
  AND U1083 ( .A(p_input[9677]), .B(p_input[39677]), .Z(n721) );
  AND U1084 ( .A(n723), .B(n724), .Z(o[9676]) );
  AND U1085 ( .A(p_input[29676]), .B(p_input[19676]), .Z(n724) );
  AND U1086 ( .A(p_input[9676]), .B(p_input[39676]), .Z(n723) );
  AND U1087 ( .A(n725), .B(n726), .Z(o[9675]) );
  AND U1088 ( .A(p_input[29675]), .B(p_input[19675]), .Z(n726) );
  AND U1089 ( .A(p_input[9675]), .B(p_input[39675]), .Z(n725) );
  AND U1090 ( .A(n727), .B(n728), .Z(o[9674]) );
  AND U1091 ( .A(p_input[29674]), .B(p_input[19674]), .Z(n728) );
  AND U1092 ( .A(p_input[9674]), .B(p_input[39674]), .Z(n727) );
  AND U1093 ( .A(n729), .B(n730), .Z(o[9673]) );
  AND U1094 ( .A(p_input[29673]), .B(p_input[19673]), .Z(n730) );
  AND U1095 ( .A(p_input[9673]), .B(p_input[39673]), .Z(n729) );
  AND U1096 ( .A(n731), .B(n732), .Z(o[9672]) );
  AND U1097 ( .A(p_input[29672]), .B(p_input[19672]), .Z(n732) );
  AND U1098 ( .A(p_input[9672]), .B(p_input[39672]), .Z(n731) );
  AND U1099 ( .A(n733), .B(n734), .Z(o[9671]) );
  AND U1100 ( .A(p_input[29671]), .B(p_input[19671]), .Z(n734) );
  AND U1101 ( .A(p_input[9671]), .B(p_input[39671]), .Z(n733) );
  AND U1102 ( .A(n735), .B(n736), .Z(o[9670]) );
  AND U1103 ( .A(p_input[29670]), .B(p_input[19670]), .Z(n736) );
  AND U1104 ( .A(p_input[9670]), .B(p_input[39670]), .Z(n735) );
  AND U1105 ( .A(n737), .B(n738), .Z(o[966]) );
  AND U1106 ( .A(p_input[20966]), .B(p_input[10966]), .Z(n738) );
  AND U1107 ( .A(p_input[966]), .B(p_input[30966]), .Z(n737) );
  AND U1108 ( .A(n739), .B(n740), .Z(o[9669]) );
  AND U1109 ( .A(p_input[29669]), .B(p_input[19669]), .Z(n740) );
  AND U1110 ( .A(p_input[9669]), .B(p_input[39669]), .Z(n739) );
  AND U1111 ( .A(n741), .B(n742), .Z(o[9668]) );
  AND U1112 ( .A(p_input[29668]), .B(p_input[19668]), .Z(n742) );
  AND U1113 ( .A(p_input[9668]), .B(p_input[39668]), .Z(n741) );
  AND U1114 ( .A(n743), .B(n744), .Z(o[9667]) );
  AND U1115 ( .A(p_input[29667]), .B(p_input[19667]), .Z(n744) );
  AND U1116 ( .A(p_input[9667]), .B(p_input[39667]), .Z(n743) );
  AND U1117 ( .A(n745), .B(n746), .Z(o[9666]) );
  AND U1118 ( .A(p_input[29666]), .B(p_input[19666]), .Z(n746) );
  AND U1119 ( .A(p_input[9666]), .B(p_input[39666]), .Z(n745) );
  AND U1120 ( .A(n747), .B(n748), .Z(o[9665]) );
  AND U1121 ( .A(p_input[29665]), .B(p_input[19665]), .Z(n748) );
  AND U1122 ( .A(p_input[9665]), .B(p_input[39665]), .Z(n747) );
  AND U1123 ( .A(n749), .B(n750), .Z(o[9664]) );
  AND U1124 ( .A(p_input[29664]), .B(p_input[19664]), .Z(n750) );
  AND U1125 ( .A(p_input[9664]), .B(p_input[39664]), .Z(n749) );
  AND U1126 ( .A(n751), .B(n752), .Z(o[9663]) );
  AND U1127 ( .A(p_input[29663]), .B(p_input[19663]), .Z(n752) );
  AND U1128 ( .A(p_input[9663]), .B(p_input[39663]), .Z(n751) );
  AND U1129 ( .A(n753), .B(n754), .Z(o[9662]) );
  AND U1130 ( .A(p_input[29662]), .B(p_input[19662]), .Z(n754) );
  AND U1131 ( .A(p_input[9662]), .B(p_input[39662]), .Z(n753) );
  AND U1132 ( .A(n755), .B(n756), .Z(o[9661]) );
  AND U1133 ( .A(p_input[29661]), .B(p_input[19661]), .Z(n756) );
  AND U1134 ( .A(p_input[9661]), .B(p_input[39661]), .Z(n755) );
  AND U1135 ( .A(n757), .B(n758), .Z(o[9660]) );
  AND U1136 ( .A(p_input[29660]), .B(p_input[19660]), .Z(n758) );
  AND U1137 ( .A(p_input[9660]), .B(p_input[39660]), .Z(n757) );
  AND U1138 ( .A(n759), .B(n760), .Z(o[965]) );
  AND U1139 ( .A(p_input[20965]), .B(p_input[10965]), .Z(n760) );
  AND U1140 ( .A(p_input[965]), .B(p_input[30965]), .Z(n759) );
  AND U1141 ( .A(n761), .B(n762), .Z(o[9659]) );
  AND U1142 ( .A(p_input[29659]), .B(p_input[19659]), .Z(n762) );
  AND U1143 ( .A(p_input[9659]), .B(p_input[39659]), .Z(n761) );
  AND U1144 ( .A(n763), .B(n764), .Z(o[9658]) );
  AND U1145 ( .A(p_input[29658]), .B(p_input[19658]), .Z(n764) );
  AND U1146 ( .A(p_input[9658]), .B(p_input[39658]), .Z(n763) );
  AND U1147 ( .A(n765), .B(n766), .Z(o[9657]) );
  AND U1148 ( .A(p_input[29657]), .B(p_input[19657]), .Z(n766) );
  AND U1149 ( .A(p_input[9657]), .B(p_input[39657]), .Z(n765) );
  AND U1150 ( .A(n767), .B(n768), .Z(o[9656]) );
  AND U1151 ( .A(p_input[29656]), .B(p_input[19656]), .Z(n768) );
  AND U1152 ( .A(p_input[9656]), .B(p_input[39656]), .Z(n767) );
  AND U1153 ( .A(n769), .B(n770), .Z(o[9655]) );
  AND U1154 ( .A(p_input[29655]), .B(p_input[19655]), .Z(n770) );
  AND U1155 ( .A(p_input[9655]), .B(p_input[39655]), .Z(n769) );
  AND U1156 ( .A(n771), .B(n772), .Z(o[9654]) );
  AND U1157 ( .A(p_input[29654]), .B(p_input[19654]), .Z(n772) );
  AND U1158 ( .A(p_input[9654]), .B(p_input[39654]), .Z(n771) );
  AND U1159 ( .A(n773), .B(n774), .Z(o[9653]) );
  AND U1160 ( .A(p_input[29653]), .B(p_input[19653]), .Z(n774) );
  AND U1161 ( .A(p_input[9653]), .B(p_input[39653]), .Z(n773) );
  AND U1162 ( .A(n775), .B(n776), .Z(o[9652]) );
  AND U1163 ( .A(p_input[29652]), .B(p_input[19652]), .Z(n776) );
  AND U1164 ( .A(p_input[9652]), .B(p_input[39652]), .Z(n775) );
  AND U1165 ( .A(n777), .B(n778), .Z(o[9651]) );
  AND U1166 ( .A(p_input[29651]), .B(p_input[19651]), .Z(n778) );
  AND U1167 ( .A(p_input[9651]), .B(p_input[39651]), .Z(n777) );
  AND U1168 ( .A(n779), .B(n780), .Z(o[9650]) );
  AND U1169 ( .A(p_input[29650]), .B(p_input[19650]), .Z(n780) );
  AND U1170 ( .A(p_input[9650]), .B(p_input[39650]), .Z(n779) );
  AND U1171 ( .A(n781), .B(n782), .Z(o[964]) );
  AND U1172 ( .A(p_input[20964]), .B(p_input[10964]), .Z(n782) );
  AND U1173 ( .A(p_input[964]), .B(p_input[30964]), .Z(n781) );
  AND U1174 ( .A(n783), .B(n784), .Z(o[9649]) );
  AND U1175 ( .A(p_input[29649]), .B(p_input[19649]), .Z(n784) );
  AND U1176 ( .A(p_input[9649]), .B(p_input[39649]), .Z(n783) );
  AND U1177 ( .A(n785), .B(n786), .Z(o[9648]) );
  AND U1178 ( .A(p_input[29648]), .B(p_input[19648]), .Z(n786) );
  AND U1179 ( .A(p_input[9648]), .B(p_input[39648]), .Z(n785) );
  AND U1180 ( .A(n787), .B(n788), .Z(o[9647]) );
  AND U1181 ( .A(p_input[29647]), .B(p_input[19647]), .Z(n788) );
  AND U1182 ( .A(p_input[9647]), .B(p_input[39647]), .Z(n787) );
  AND U1183 ( .A(n789), .B(n790), .Z(o[9646]) );
  AND U1184 ( .A(p_input[29646]), .B(p_input[19646]), .Z(n790) );
  AND U1185 ( .A(p_input[9646]), .B(p_input[39646]), .Z(n789) );
  AND U1186 ( .A(n791), .B(n792), .Z(o[9645]) );
  AND U1187 ( .A(p_input[29645]), .B(p_input[19645]), .Z(n792) );
  AND U1188 ( .A(p_input[9645]), .B(p_input[39645]), .Z(n791) );
  AND U1189 ( .A(n793), .B(n794), .Z(o[9644]) );
  AND U1190 ( .A(p_input[29644]), .B(p_input[19644]), .Z(n794) );
  AND U1191 ( .A(p_input[9644]), .B(p_input[39644]), .Z(n793) );
  AND U1192 ( .A(n795), .B(n796), .Z(o[9643]) );
  AND U1193 ( .A(p_input[29643]), .B(p_input[19643]), .Z(n796) );
  AND U1194 ( .A(p_input[9643]), .B(p_input[39643]), .Z(n795) );
  AND U1195 ( .A(n797), .B(n798), .Z(o[9642]) );
  AND U1196 ( .A(p_input[29642]), .B(p_input[19642]), .Z(n798) );
  AND U1197 ( .A(p_input[9642]), .B(p_input[39642]), .Z(n797) );
  AND U1198 ( .A(n799), .B(n800), .Z(o[9641]) );
  AND U1199 ( .A(p_input[29641]), .B(p_input[19641]), .Z(n800) );
  AND U1200 ( .A(p_input[9641]), .B(p_input[39641]), .Z(n799) );
  AND U1201 ( .A(n801), .B(n802), .Z(o[9640]) );
  AND U1202 ( .A(p_input[29640]), .B(p_input[19640]), .Z(n802) );
  AND U1203 ( .A(p_input[9640]), .B(p_input[39640]), .Z(n801) );
  AND U1204 ( .A(n803), .B(n804), .Z(o[963]) );
  AND U1205 ( .A(p_input[20963]), .B(p_input[10963]), .Z(n804) );
  AND U1206 ( .A(p_input[963]), .B(p_input[30963]), .Z(n803) );
  AND U1207 ( .A(n805), .B(n806), .Z(o[9639]) );
  AND U1208 ( .A(p_input[29639]), .B(p_input[19639]), .Z(n806) );
  AND U1209 ( .A(p_input[9639]), .B(p_input[39639]), .Z(n805) );
  AND U1210 ( .A(n807), .B(n808), .Z(o[9638]) );
  AND U1211 ( .A(p_input[29638]), .B(p_input[19638]), .Z(n808) );
  AND U1212 ( .A(p_input[9638]), .B(p_input[39638]), .Z(n807) );
  AND U1213 ( .A(n809), .B(n810), .Z(o[9637]) );
  AND U1214 ( .A(p_input[29637]), .B(p_input[19637]), .Z(n810) );
  AND U1215 ( .A(p_input[9637]), .B(p_input[39637]), .Z(n809) );
  AND U1216 ( .A(n811), .B(n812), .Z(o[9636]) );
  AND U1217 ( .A(p_input[29636]), .B(p_input[19636]), .Z(n812) );
  AND U1218 ( .A(p_input[9636]), .B(p_input[39636]), .Z(n811) );
  AND U1219 ( .A(n813), .B(n814), .Z(o[9635]) );
  AND U1220 ( .A(p_input[29635]), .B(p_input[19635]), .Z(n814) );
  AND U1221 ( .A(p_input[9635]), .B(p_input[39635]), .Z(n813) );
  AND U1222 ( .A(n815), .B(n816), .Z(o[9634]) );
  AND U1223 ( .A(p_input[29634]), .B(p_input[19634]), .Z(n816) );
  AND U1224 ( .A(p_input[9634]), .B(p_input[39634]), .Z(n815) );
  AND U1225 ( .A(n817), .B(n818), .Z(o[9633]) );
  AND U1226 ( .A(p_input[29633]), .B(p_input[19633]), .Z(n818) );
  AND U1227 ( .A(p_input[9633]), .B(p_input[39633]), .Z(n817) );
  AND U1228 ( .A(n819), .B(n820), .Z(o[9632]) );
  AND U1229 ( .A(p_input[29632]), .B(p_input[19632]), .Z(n820) );
  AND U1230 ( .A(p_input[9632]), .B(p_input[39632]), .Z(n819) );
  AND U1231 ( .A(n821), .B(n822), .Z(o[9631]) );
  AND U1232 ( .A(p_input[29631]), .B(p_input[19631]), .Z(n822) );
  AND U1233 ( .A(p_input[9631]), .B(p_input[39631]), .Z(n821) );
  AND U1234 ( .A(n823), .B(n824), .Z(o[9630]) );
  AND U1235 ( .A(p_input[29630]), .B(p_input[19630]), .Z(n824) );
  AND U1236 ( .A(p_input[9630]), .B(p_input[39630]), .Z(n823) );
  AND U1237 ( .A(n825), .B(n826), .Z(o[962]) );
  AND U1238 ( .A(p_input[20962]), .B(p_input[10962]), .Z(n826) );
  AND U1239 ( .A(p_input[962]), .B(p_input[30962]), .Z(n825) );
  AND U1240 ( .A(n827), .B(n828), .Z(o[9629]) );
  AND U1241 ( .A(p_input[29629]), .B(p_input[19629]), .Z(n828) );
  AND U1242 ( .A(p_input[9629]), .B(p_input[39629]), .Z(n827) );
  AND U1243 ( .A(n829), .B(n830), .Z(o[9628]) );
  AND U1244 ( .A(p_input[29628]), .B(p_input[19628]), .Z(n830) );
  AND U1245 ( .A(p_input[9628]), .B(p_input[39628]), .Z(n829) );
  AND U1246 ( .A(n831), .B(n832), .Z(o[9627]) );
  AND U1247 ( .A(p_input[29627]), .B(p_input[19627]), .Z(n832) );
  AND U1248 ( .A(p_input[9627]), .B(p_input[39627]), .Z(n831) );
  AND U1249 ( .A(n833), .B(n834), .Z(o[9626]) );
  AND U1250 ( .A(p_input[29626]), .B(p_input[19626]), .Z(n834) );
  AND U1251 ( .A(p_input[9626]), .B(p_input[39626]), .Z(n833) );
  AND U1252 ( .A(n835), .B(n836), .Z(o[9625]) );
  AND U1253 ( .A(p_input[29625]), .B(p_input[19625]), .Z(n836) );
  AND U1254 ( .A(p_input[9625]), .B(p_input[39625]), .Z(n835) );
  AND U1255 ( .A(n837), .B(n838), .Z(o[9624]) );
  AND U1256 ( .A(p_input[29624]), .B(p_input[19624]), .Z(n838) );
  AND U1257 ( .A(p_input[9624]), .B(p_input[39624]), .Z(n837) );
  AND U1258 ( .A(n839), .B(n840), .Z(o[9623]) );
  AND U1259 ( .A(p_input[29623]), .B(p_input[19623]), .Z(n840) );
  AND U1260 ( .A(p_input[9623]), .B(p_input[39623]), .Z(n839) );
  AND U1261 ( .A(n841), .B(n842), .Z(o[9622]) );
  AND U1262 ( .A(p_input[29622]), .B(p_input[19622]), .Z(n842) );
  AND U1263 ( .A(p_input[9622]), .B(p_input[39622]), .Z(n841) );
  AND U1264 ( .A(n843), .B(n844), .Z(o[9621]) );
  AND U1265 ( .A(p_input[29621]), .B(p_input[19621]), .Z(n844) );
  AND U1266 ( .A(p_input[9621]), .B(p_input[39621]), .Z(n843) );
  AND U1267 ( .A(n845), .B(n846), .Z(o[9620]) );
  AND U1268 ( .A(p_input[29620]), .B(p_input[19620]), .Z(n846) );
  AND U1269 ( .A(p_input[9620]), .B(p_input[39620]), .Z(n845) );
  AND U1270 ( .A(n847), .B(n848), .Z(o[961]) );
  AND U1271 ( .A(p_input[20961]), .B(p_input[10961]), .Z(n848) );
  AND U1272 ( .A(p_input[961]), .B(p_input[30961]), .Z(n847) );
  AND U1273 ( .A(n849), .B(n850), .Z(o[9619]) );
  AND U1274 ( .A(p_input[29619]), .B(p_input[19619]), .Z(n850) );
  AND U1275 ( .A(p_input[9619]), .B(p_input[39619]), .Z(n849) );
  AND U1276 ( .A(n851), .B(n852), .Z(o[9618]) );
  AND U1277 ( .A(p_input[29618]), .B(p_input[19618]), .Z(n852) );
  AND U1278 ( .A(p_input[9618]), .B(p_input[39618]), .Z(n851) );
  AND U1279 ( .A(n853), .B(n854), .Z(o[9617]) );
  AND U1280 ( .A(p_input[29617]), .B(p_input[19617]), .Z(n854) );
  AND U1281 ( .A(p_input[9617]), .B(p_input[39617]), .Z(n853) );
  AND U1282 ( .A(n855), .B(n856), .Z(o[9616]) );
  AND U1283 ( .A(p_input[29616]), .B(p_input[19616]), .Z(n856) );
  AND U1284 ( .A(p_input[9616]), .B(p_input[39616]), .Z(n855) );
  AND U1285 ( .A(n857), .B(n858), .Z(o[9615]) );
  AND U1286 ( .A(p_input[29615]), .B(p_input[19615]), .Z(n858) );
  AND U1287 ( .A(p_input[9615]), .B(p_input[39615]), .Z(n857) );
  AND U1288 ( .A(n859), .B(n860), .Z(o[9614]) );
  AND U1289 ( .A(p_input[29614]), .B(p_input[19614]), .Z(n860) );
  AND U1290 ( .A(p_input[9614]), .B(p_input[39614]), .Z(n859) );
  AND U1291 ( .A(n861), .B(n862), .Z(o[9613]) );
  AND U1292 ( .A(p_input[29613]), .B(p_input[19613]), .Z(n862) );
  AND U1293 ( .A(p_input[9613]), .B(p_input[39613]), .Z(n861) );
  AND U1294 ( .A(n863), .B(n864), .Z(o[9612]) );
  AND U1295 ( .A(p_input[29612]), .B(p_input[19612]), .Z(n864) );
  AND U1296 ( .A(p_input[9612]), .B(p_input[39612]), .Z(n863) );
  AND U1297 ( .A(n865), .B(n866), .Z(o[9611]) );
  AND U1298 ( .A(p_input[29611]), .B(p_input[19611]), .Z(n866) );
  AND U1299 ( .A(p_input[9611]), .B(p_input[39611]), .Z(n865) );
  AND U1300 ( .A(n867), .B(n868), .Z(o[9610]) );
  AND U1301 ( .A(p_input[29610]), .B(p_input[19610]), .Z(n868) );
  AND U1302 ( .A(p_input[9610]), .B(p_input[39610]), .Z(n867) );
  AND U1303 ( .A(n869), .B(n870), .Z(o[960]) );
  AND U1304 ( .A(p_input[20960]), .B(p_input[10960]), .Z(n870) );
  AND U1305 ( .A(p_input[960]), .B(p_input[30960]), .Z(n869) );
  AND U1306 ( .A(n871), .B(n872), .Z(o[9609]) );
  AND U1307 ( .A(p_input[29609]), .B(p_input[19609]), .Z(n872) );
  AND U1308 ( .A(p_input[9609]), .B(p_input[39609]), .Z(n871) );
  AND U1309 ( .A(n873), .B(n874), .Z(o[9608]) );
  AND U1310 ( .A(p_input[29608]), .B(p_input[19608]), .Z(n874) );
  AND U1311 ( .A(p_input[9608]), .B(p_input[39608]), .Z(n873) );
  AND U1312 ( .A(n875), .B(n876), .Z(o[9607]) );
  AND U1313 ( .A(p_input[29607]), .B(p_input[19607]), .Z(n876) );
  AND U1314 ( .A(p_input[9607]), .B(p_input[39607]), .Z(n875) );
  AND U1315 ( .A(n877), .B(n878), .Z(o[9606]) );
  AND U1316 ( .A(p_input[29606]), .B(p_input[19606]), .Z(n878) );
  AND U1317 ( .A(p_input[9606]), .B(p_input[39606]), .Z(n877) );
  AND U1318 ( .A(n879), .B(n880), .Z(o[9605]) );
  AND U1319 ( .A(p_input[29605]), .B(p_input[19605]), .Z(n880) );
  AND U1320 ( .A(p_input[9605]), .B(p_input[39605]), .Z(n879) );
  AND U1321 ( .A(n881), .B(n882), .Z(o[9604]) );
  AND U1322 ( .A(p_input[29604]), .B(p_input[19604]), .Z(n882) );
  AND U1323 ( .A(p_input[9604]), .B(p_input[39604]), .Z(n881) );
  AND U1324 ( .A(n883), .B(n884), .Z(o[9603]) );
  AND U1325 ( .A(p_input[29603]), .B(p_input[19603]), .Z(n884) );
  AND U1326 ( .A(p_input[9603]), .B(p_input[39603]), .Z(n883) );
  AND U1327 ( .A(n885), .B(n886), .Z(o[9602]) );
  AND U1328 ( .A(p_input[29602]), .B(p_input[19602]), .Z(n886) );
  AND U1329 ( .A(p_input[9602]), .B(p_input[39602]), .Z(n885) );
  AND U1330 ( .A(n887), .B(n888), .Z(o[9601]) );
  AND U1331 ( .A(p_input[29601]), .B(p_input[19601]), .Z(n888) );
  AND U1332 ( .A(p_input[9601]), .B(p_input[39601]), .Z(n887) );
  AND U1333 ( .A(n889), .B(n890), .Z(o[9600]) );
  AND U1334 ( .A(p_input[29600]), .B(p_input[19600]), .Z(n890) );
  AND U1335 ( .A(p_input[9600]), .B(p_input[39600]), .Z(n889) );
  AND U1336 ( .A(n891), .B(n892), .Z(o[95]) );
  AND U1337 ( .A(p_input[20095]), .B(p_input[10095]), .Z(n892) );
  AND U1338 ( .A(p_input[95]), .B(p_input[30095]), .Z(n891) );
  AND U1339 ( .A(n893), .B(n894), .Z(o[959]) );
  AND U1340 ( .A(p_input[20959]), .B(p_input[10959]), .Z(n894) );
  AND U1341 ( .A(p_input[959]), .B(p_input[30959]), .Z(n893) );
  AND U1342 ( .A(n895), .B(n896), .Z(o[9599]) );
  AND U1343 ( .A(p_input[29599]), .B(p_input[19599]), .Z(n896) );
  AND U1344 ( .A(p_input[9599]), .B(p_input[39599]), .Z(n895) );
  AND U1345 ( .A(n897), .B(n898), .Z(o[9598]) );
  AND U1346 ( .A(p_input[29598]), .B(p_input[19598]), .Z(n898) );
  AND U1347 ( .A(p_input[9598]), .B(p_input[39598]), .Z(n897) );
  AND U1348 ( .A(n899), .B(n900), .Z(o[9597]) );
  AND U1349 ( .A(p_input[29597]), .B(p_input[19597]), .Z(n900) );
  AND U1350 ( .A(p_input[9597]), .B(p_input[39597]), .Z(n899) );
  AND U1351 ( .A(n901), .B(n902), .Z(o[9596]) );
  AND U1352 ( .A(p_input[29596]), .B(p_input[19596]), .Z(n902) );
  AND U1353 ( .A(p_input[9596]), .B(p_input[39596]), .Z(n901) );
  AND U1354 ( .A(n903), .B(n904), .Z(o[9595]) );
  AND U1355 ( .A(p_input[29595]), .B(p_input[19595]), .Z(n904) );
  AND U1356 ( .A(p_input[9595]), .B(p_input[39595]), .Z(n903) );
  AND U1357 ( .A(n905), .B(n906), .Z(o[9594]) );
  AND U1358 ( .A(p_input[29594]), .B(p_input[19594]), .Z(n906) );
  AND U1359 ( .A(p_input[9594]), .B(p_input[39594]), .Z(n905) );
  AND U1360 ( .A(n907), .B(n908), .Z(o[9593]) );
  AND U1361 ( .A(p_input[29593]), .B(p_input[19593]), .Z(n908) );
  AND U1362 ( .A(p_input[9593]), .B(p_input[39593]), .Z(n907) );
  AND U1363 ( .A(n909), .B(n910), .Z(o[9592]) );
  AND U1364 ( .A(p_input[29592]), .B(p_input[19592]), .Z(n910) );
  AND U1365 ( .A(p_input[9592]), .B(p_input[39592]), .Z(n909) );
  AND U1366 ( .A(n911), .B(n912), .Z(o[9591]) );
  AND U1367 ( .A(p_input[29591]), .B(p_input[19591]), .Z(n912) );
  AND U1368 ( .A(p_input[9591]), .B(p_input[39591]), .Z(n911) );
  AND U1369 ( .A(n913), .B(n914), .Z(o[9590]) );
  AND U1370 ( .A(p_input[29590]), .B(p_input[19590]), .Z(n914) );
  AND U1371 ( .A(p_input[9590]), .B(p_input[39590]), .Z(n913) );
  AND U1372 ( .A(n915), .B(n916), .Z(o[958]) );
  AND U1373 ( .A(p_input[20958]), .B(p_input[10958]), .Z(n916) );
  AND U1374 ( .A(p_input[958]), .B(p_input[30958]), .Z(n915) );
  AND U1375 ( .A(n917), .B(n918), .Z(o[9589]) );
  AND U1376 ( .A(p_input[29589]), .B(p_input[19589]), .Z(n918) );
  AND U1377 ( .A(p_input[9589]), .B(p_input[39589]), .Z(n917) );
  AND U1378 ( .A(n919), .B(n920), .Z(o[9588]) );
  AND U1379 ( .A(p_input[29588]), .B(p_input[19588]), .Z(n920) );
  AND U1380 ( .A(p_input[9588]), .B(p_input[39588]), .Z(n919) );
  AND U1381 ( .A(n921), .B(n922), .Z(o[9587]) );
  AND U1382 ( .A(p_input[29587]), .B(p_input[19587]), .Z(n922) );
  AND U1383 ( .A(p_input[9587]), .B(p_input[39587]), .Z(n921) );
  AND U1384 ( .A(n923), .B(n924), .Z(o[9586]) );
  AND U1385 ( .A(p_input[29586]), .B(p_input[19586]), .Z(n924) );
  AND U1386 ( .A(p_input[9586]), .B(p_input[39586]), .Z(n923) );
  AND U1387 ( .A(n925), .B(n926), .Z(o[9585]) );
  AND U1388 ( .A(p_input[29585]), .B(p_input[19585]), .Z(n926) );
  AND U1389 ( .A(p_input[9585]), .B(p_input[39585]), .Z(n925) );
  AND U1390 ( .A(n927), .B(n928), .Z(o[9584]) );
  AND U1391 ( .A(p_input[29584]), .B(p_input[19584]), .Z(n928) );
  AND U1392 ( .A(p_input[9584]), .B(p_input[39584]), .Z(n927) );
  AND U1393 ( .A(n929), .B(n930), .Z(o[9583]) );
  AND U1394 ( .A(p_input[29583]), .B(p_input[19583]), .Z(n930) );
  AND U1395 ( .A(p_input[9583]), .B(p_input[39583]), .Z(n929) );
  AND U1396 ( .A(n931), .B(n932), .Z(o[9582]) );
  AND U1397 ( .A(p_input[29582]), .B(p_input[19582]), .Z(n932) );
  AND U1398 ( .A(p_input[9582]), .B(p_input[39582]), .Z(n931) );
  AND U1399 ( .A(n933), .B(n934), .Z(o[9581]) );
  AND U1400 ( .A(p_input[29581]), .B(p_input[19581]), .Z(n934) );
  AND U1401 ( .A(p_input[9581]), .B(p_input[39581]), .Z(n933) );
  AND U1402 ( .A(n935), .B(n936), .Z(o[9580]) );
  AND U1403 ( .A(p_input[29580]), .B(p_input[19580]), .Z(n936) );
  AND U1404 ( .A(p_input[9580]), .B(p_input[39580]), .Z(n935) );
  AND U1405 ( .A(n937), .B(n938), .Z(o[957]) );
  AND U1406 ( .A(p_input[20957]), .B(p_input[10957]), .Z(n938) );
  AND U1407 ( .A(p_input[957]), .B(p_input[30957]), .Z(n937) );
  AND U1408 ( .A(n939), .B(n940), .Z(o[9579]) );
  AND U1409 ( .A(p_input[29579]), .B(p_input[19579]), .Z(n940) );
  AND U1410 ( .A(p_input[9579]), .B(p_input[39579]), .Z(n939) );
  AND U1411 ( .A(n941), .B(n942), .Z(o[9578]) );
  AND U1412 ( .A(p_input[29578]), .B(p_input[19578]), .Z(n942) );
  AND U1413 ( .A(p_input[9578]), .B(p_input[39578]), .Z(n941) );
  AND U1414 ( .A(n943), .B(n944), .Z(o[9577]) );
  AND U1415 ( .A(p_input[29577]), .B(p_input[19577]), .Z(n944) );
  AND U1416 ( .A(p_input[9577]), .B(p_input[39577]), .Z(n943) );
  AND U1417 ( .A(n945), .B(n946), .Z(o[9576]) );
  AND U1418 ( .A(p_input[29576]), .B(p_input[19576]), .Z(n946) );
  AND U1419 ( .A(p_input[9576]), .B(p_input[39576]), .Z(n945) );
  AND U1420 ( .A(n947), .B(n948), .Z(o[9575]) );
  AND U1421 ( .A(p_input[29575]), .B(p_input[19575]), .Z(n948) );
  AND U1422 ( .A(p_input[9575]), .B(p_input[39575]), .Z(n947) );
  AND U1423 ( .A(n949), .B(n950), .Z(o[9574]) );
  AND U1424 ( .A(p_input[29574]), .B(p_input[19574]), .Z(n950) );
  AND U1425 ( .A(p_input[9574]), .B(p_input[39574]), .Z(n949) );
  AND U1426 ( .A(n951), .B(n952), .Z(o[9573]) );
  AND U1427 ( .A(p_input[29573]), .B(p_input[19573]), .Z(n952) );
  AND U1428 ( .A(p_input[9573]), .B(p_input[39573]), .Z(n951) );
  AND U1429 ( .A(n953), .B(n954), .Z(o[9572]) );
  AND U1430 ( .A(p_input[29572]), .B(p_input[19572]), .Z(n954) );
  AND U1431 ( .A(p_input[9572]), .B(p_input[39572]), .Z(n953) );
  AND U1432 ( .A(n955), .B(n956), .Z(o[9571]) );
  AND U1433 ( .A(p_input[29571]), .B(p_input[19571]), .Z(n956) );
  AND U1434 ( .A(p_input[9571]), .B(p_input[39571]), .Z(n955) );
  AND U1435 ( .A(n957), .B(n958), .Z(o[9570]) );
  AND U1436 ( .A(p_input[29570]), .B(p_input[19570]), .Z(n958) );
  AND U1437 ( .A(p_input[9570]), .B(p_input[39570]), .Z(n957) );
  AND U1438 ( .A(n959), .B(n960), .Z(o[956]) );
  AND U1439 ( .A(p_input[20956]), .B(p_input[10956]), .Z(n960) );
  AND U1440 ( .A(p_input[956]), .B(p_input[30956]), .Z(n959) );
  AND U1441 ( .A(n961), .B(n962), .Z(o[9569]) );
  AND U1442 ( .A(p_input[29569]), .B(p_input[19569]), .Z(n962) );
  AND U1443 ( .A(p_input[9569]), .B(p_input[39569]), .Z(n961) );
  AND U1444 ( .A(n963), .B(n964), .Z(o[9568]) );
  AND U1445 ( .A(p_input[29568]), .B(p_input[19568]), .Z(n964) );
  AND U1446 ( .A(p_input[9568]), .B(p_input[39568]), .Z(n963) );
  AND U1447 ( .A(n965), .B(n966), .Z(o[9567]) );
  AND U1448 ( .A(p_input[29567]), .B(p_input[19567]), .Z(n966) );
  AND U1449 ( .A(p_input[9567]), .B(p_input[39567]), .Z(n965) );
  AND U1450 ( .A(n967), .B(n968), .Z(o[9566]) );
  AND U1451 ( .A(p_input[29566]), .B(p_input[19566]), .Z(n968) );
  AND U1452 ( .A(p_input[9566]), .B(p_input[39566]), .Z(n967) );
  AND U1453 ( .A(n969), .B(n970), .Z(o[9565]) );
  AND U1454 ( .A(p_input[29565]), .B(p_input[19565]), .Z(n970) );
  AND U1455 ( .A(p_input[9565]), .B(p_input[39565]), .Z(n969) );
  AND U1456 ( .A(n971), .B(n972), .Z(o[9564]) );
  AND U1457 ( .A(p_input[29564]), .B(p_input[19564]), .Z(n972) );
  AND U1458 ( .A(p_input[9564]), .B(p_input[39564]), .Z(n971) );
  AND U1459 ( .A(n973), .B(n974), .Z(o[9563]) );
  AND U1460 ( .A(p_input[29563]), .B(p_input[19563]), .Z(n974) );
  AND U1461 ( .A(p_input[9563]), .B(p_input[39563]), .Z(n973) );
  AND U1462 ( .A(n975), .B(n976), .Z(o[9562]) );
  AND U1463 ( .A(p_input[29562]), .B(p_input[19562]), .Z(n976) );
  AND U1464 ( .A(p_input[9562]), .B(p_input[39562]), .Z(n975) );
  AND U1465 ( .A(n977), .B(n978), .Z(o[9561]) );
  AND U1466 ( .A(p_input[29561]), .B(p_input[19561]), .Z(n978) );
  AND U1467 ( .A(p_input[9561]), .B(p_input[39561]), .Z(n977) );
  AND U1468 ( .A(n979), .B(n980), .Z(o[9560]) );
  AND U1469 ( .A(p_input[29560]), .B(p_input[19560]), .Z(n980) );
  AND U1470 ( .A(p_input[9560]), .B(p_input[39560]), .Z(n979) );
  AND U1471 ( .A(n981), .B(n982), .Z(o[955]) );
  AND U1472 ( .A(p_input[20955]), .B(p_input[10955]), .Z(n982) );
  AND U1473 ( .A(p_input[955]), .B(p_input[30955]), .Z(n981) );
  AND U1474 ( .A(n983), .B(n984), .Z(o[9559]) );
  AND U1475 ( .A(p_input[29559]), .B(p_input[19559]), .Z(n984) );
  AND U1476 ( .A(p_input[9559]), .B(p_input[39559]), .Z(n983) );
  AND U1477 ( .A(n985), .B(n986), .Z(o[9558]) );
  AND U1478 ( .A(p_input[29558]), .B(p_input[19558]), .Z(n986) );
  AND U1479 ( .A(p_input[9558]), .B(p_input[39558]), .Z(n985) );
  AND U1480 ( .A(n987), .B(n988), .Z(o[9557]) );
  AND U1481 ( .A(p_input[29557]), .B(p_input[19557]), .Z(n988) );
  AND U1482 ( .A(p_input[9557]), .B(p_input[39557]), .Z(n987) );
  AND U1483 ( .A(n989), .B(n990), .Z(o[9556]) );
  AND U1484 ( .A(p_input[29556]), .B(p_input[19556]), .Z(n990) );
  AND U1485 ( .A(p_input[9556]), .B(p_input[39556]), .Z(n989) );
  AND U1486 ( .A(n991), .B(n992), .Z(o[9555]) );
  AND U1487 ( .A(p_input[29555]), .B(p_input[19555]), .Z(n992) );
  AND U1488 ( .A(p_input[9555]), .B(p_input[39555]), .Z(n991) );
  AND U1489 ( .A(n993), .B(n994), .Z(o[9554]) );
  AND U1490 ( .A(p_input[29554]), .B(p_input[19554]), .Z(n994) );
  AND U1491 ( .A(p_input[9554]), .B(p_input[39554]), .Z(n993) );
  AND U1492 ( .A(n995), .B(n996), .Z(o[9553]) );
  AND U1493 ( .A(p_input[29553]), .B(p_input[19553]), .Z(n996) );
  AND U1494 ( .A(p_input[9553]), .B(p_input[39553]), .Z(n995) );
  AND U1495 ( .A(n997), .B(n998), .Z(o[9552]) );
  AND U1496 ( .A(p_input[29552]), .B(p_input[19552]), .Z(n998) );
  AND U1497 ( .A(p_input[9552]), .B(p_input[39552]), .Z(n997) );
  AND U1498 ( .A(n999), .B(n1000), .Z(o[9551]) );
  AND U1499 ( .A(p_input[29551]), .B(p_input[19551]), .Z(n1000) );
  AND U1500 ( .A(p_input[9551]), .B(p_input[39551]), .Z(n999) );
  AND U1501 ( .A(n1001), .B(n1002), .Z(o[9550]) );
  AND U1502 ( .A(p_input[29550]), .B(p_input[19550]), .Z(n1002) );
  AND U1503 ( .A(p_input[9550]), .B(p_input[39550]), .Z(n1001) );
  AND U1504 ( .A(n1003), .B(n1004), .Z(o[954]) );
  AND U1505 ( .A(p_input[20954]), .B(p_input[10954]), .Z(n1004) );
  AND U1506 ( .A(p_input[954]), .B(p_input[30954]), .Z(n1003) );
  AND U1507 ( .A(n1005), .B(n1006), .Z(o[9549]) );
  AND U1508 ( .A(p_input[29549]), .B(p_input[19549]), .Z(n1006) );
  AND U1509 ( .A(p_input[9549]), .B(p_input[39549]), .Z(n1005) );
  AND U1510 ( .A(n1007), .B(n1008), .Z(o[9548]) );
  AND U1511 ( .A(p_input[29548]), .B(p_input[19548]), .Z(n1008) );
  AND U1512 ( .A(p_input[9548]), .B(p_input[39548]), .Z(n1007) );
  AND U1513 ( .A(n1009), .B(n1010), .Z(o[9547]) );
  AND U1514 ( .A(p_input[29547]), .B(p_input[19547]), .Z(n1010) );
  AND U1515 ( .A(p_input[9547]), .B(p_input[39547]), .Z(n1009) );
  AND U1516 ( .A(n1011), .B(n1012), .Z(o[9546]) );
  AND U1517 ( .A(p_input[29546]), .B(p_input[19546]), .Z(n1012) );
  AND U1518 ( .A(p_input[9546]), .B(p_input[39546]), .Z(n1011) );
  AND U1519 ( .A(n1013), .B(n1014), .Z(o[9545]) );
  AND U1520 ( .A(p_input[29545]), .B(p_input[19545]), .Z(n1014) );
  AND U1521 ( .A(p_input[9545]), .B(p_input[39545]), .Z(n1013) );
  AND U1522 ( .A(n1015), .B(n1016), .Z(o[9544]) );
  AND U1523 ( .A(p_input[29544]), .B(p_input[19544]), .Z(n1016) );
  AND U1524 ( .A(p_input[9544]), .B(p_input[39544]), .Z(n1015) );
  AND U1525 ( .A(n1017), .B(n1018), .Z(o[9543]) );
  AND U1526 ( .A(p_input[29543]), .B(p_input[19543]), .Z(n1018) );
  AND U1527 ( .A(p_input[9543]), .B(p_input[39543]), .Z(n1017) );
  AND U1528 ( .A(n1019), .B(n1020), .Z(o[9542]) );
  AND U1529 ( .A(p_input[29542]), .B(p_input[19542]), .Z(n1020) );
  AND U1530 ( .A(p_input[9542]), .B(p_input[39542]), .Z(n1019) );
  AND U1531 ( .A(n1021), .B(n1022), .Z(o[9541]) );
  AND U1532 ( .A(p_input[29541]), .B(p_input[19541]), .Z(n1022) );
  AND U1533 ( .A(p_input[9541]), .B(p_input[39541]), .Z(n1021) );
  AND U1534 ( .A(n1023), .B(n1024), .Z(o[9540]) );
  AND U1535 ( .A(p_input[29540]), .B(p_input[19540]), .Z(n1024) );
  AND U1536 ( .A(p_input[9540]), .B(p_input[39540]), .Z(n1023) );
  AND U1537 ( .A(n1025), .B(n1026), .Z(o[953]) );
  AND U1538 ( .A(p_input[20953]), .B(p_input[10953]), .Z(n1026) );
  AND U1539 ( .A(p_input[953]), .B(p_input[30953]), .Z(n1025) );
  AND U1540 ( .A(n1027), .B(n1028), .Z(o[9539]) );
  AND U1541 ( .A(p_input[29539]), .B(p_input[19539]), .Z(n1028) );
  AND U1542 ( .A(p_input[9539]), .B(p_input[39539]), .Z(n1027) );
  AND U1543 ( .A(n1029), .B(n1030), .Z(o[9538]) );
  AND U1544 ( .A(p_input[29538]), .B(p_input[19538]), .Z(n1030) );
  AND U1545 ( .A(p_input[9538]), .B(p_input[39538]), .Z(n1029) );
  AND U1546 ( .A(n1031), .B(n1032), .Z(o[9537]) );
  AND U1547 ( .A(p_input[29537]), .B(p_input[19537]), .Z(n1032) );
  AND U1548 ( .A(p_input[9537]), .B(p_input[39537]), .Z(n1031) );
  AND U1549 ( .A(n1033), .B(n1034), .Z(o[9536]) );
  AND U1550 ( .A(p_input[29536]), .B(p_input[19536]), .Z(n1034) );
  AND U1551 ( .A(p_input[9536]), .B(p_input[39536]), .Z(n1033) );
  AND U1552 ( .A(n1035), .B(n1036), .Z(o[9535]) );
  AND U1553 ( .A(p_input[29535]), .B(p_input[19535]), .Z(n1036) );
  AND U1554 ( .A(p_input[9535]), .B(p_input[39535]), .Z(n1035) );
  AND U1555 ( .A(n1037), .B(n1038), .Z(o[9534]) );
  AND U1556 ( .A(p_input[29534]), .B(p_input[19534]), .Z(n1038) );
  AND U1557 ( .A(p_input[9534]), .B(p_input[39534]), .Z(n1037) );
  AND U1558 ( .A(n1039), .B(n1040), .Z(o[9533]) );
  AND U1559 ( .A(p_input[29533]), .B(p_input[19533]), .Z(n1040) );
  AND U1560 ( .A(p_input[9533]), .B(p_input[39533]), .Z(n1039) );
  AND U1561 ( .A(n1041), .B(n1042), .Z(o[9532]) );
  AND U1562 ( .A(p_input[29532]), .B(p_input[19532]), .Z(n1042) );
  AND U1563 ( .A(p_input[9532]), .B(p_input[39532]), .Z(n1041) );
  AND U1564 ( .A(n1043), .B(n1044), .Z(o[9531]) );
  AND U1565 ( .A(p_input[29531]), .B(p_input[19531]), .Z(n1044) );
  AND U1566 ( .A(p_input[9531]), .B(p_input[39531]), .Z(n1043) );
  AND U1567 ( .A(n1045), .B(n1046), .Z(o[9530]) );
  AND U1568 ( .A(p_input[29530]), .B(p_input[19530]), .Z(n1046) );
  AND U1569 ( .A(p_input[9530]), .B(p_input[39530]), .Z(n1045) );
  AND U1570 ( .A(n1047), .B(n1048), .Z(o[952]) );
  AND U1571 ( .A(p_input[20952]), .B(p_input[10952]), .Z(n1048) );
  AND U1572 ( .A(p_input[952]), .B(p_input[30952]), .Z(n1047) );
  AND U1573 ( .A(n1049), .B(n1050), .Z(o[9529]) );
  AND U1574 ( .A(p_input[29529]), .B(p_input[19529]), .Z(n1050) );
  AND U1575 ( .A(p_input[9529]), .B(p_input[39529]), .Z(n1049) );
  AND U1576 ( .A(n1051), .B(n1052), .Z(o[9528]) );
  AND U1577 ( .A(p_input[29528]), .B(p_input[19528]), .Z(n1052) );
  AND U1578 ( .A(p_input[9528]), .B(p_input[39528]), .Z(n1051) );
  AND U1579 ( .A(n1053), .B(n1054), .Z(o[9527]) );
  AND U1580 ( .A(p_input[29527]), .B(p_input[19527]), .Z(n1054) );
  AND U1581 ( .A(p_input[9527]), .B(p_input[39527]), .Z(n1053) );
  AND U1582 ( .A(n1055), .B(n1056), .Z(o[9526]) );
  AND U1583 ( .A(p_input[29526]), .B(p_input[19526]), .Z(n1056) );
  AND U1584 ( .A(p_input[9526]), .B(p_input[39526]), .Z(n1055) );
  AND U1585 ( .A(n1057), .B(n1058), .Z(o[9525]) );
  AND U1586 ( .A(p_input[29525]), .B(p_input[19525]), .Z(n1058) );
  AND U1587 ( .A(p_input[9525]), .B(p_input[39525]), .Z(n1057) );
  AND U1588 ( .A(n1059), .B(n1060), .Z(o[9524]) );
  AND U1589 ( .A(p_input[29524]), .B(p_input[19524]), .Z(n1060) );
  AND U1590 ( .A(p_input[9524]), .B(p_input[39524]), .Z(n1059) );
  AND U1591 ( .A(n1061), .B(n1062), .Z(o[9523]) );
  AND U1592 ( .A(p_input[29523]), .B(p_input[19523]), .Z(n1062) );
  AND U1593 ( .A(p_input[9523]), .B(p_input[39523]), .Z(n1061) );
  AND U1594 ( .A(n1063), .B(n1064), .Z(o[9522]) );
  AND U1595 ( .A(p_input[29522]), .B(p_input[19522]), .Z(n1064) );
  AND U1596 ( .A(p_input[9522]), .B(p_input[39522]), .Z(n1063) );
  AND U1597 ( .A(n1065), .B(n1066), .Z(o[9521]) );
  AND U1598 ( .A(p_input[29521]), .B(p_input[19521]), .Z(n1066) );
  AND U1599 ( .A(p_input[9521]), .B(p_input[39521]), .Z(n1065) );
  AND U1600 ( .A(n1067), .B(n1068), .Z(o[9520]) );
  AND U1601 ( .A(p_input[29520]), .B(p_input[19520]), .Z(n1068) );
  AND U1602 ( .A(p_input[9520]), .B(p_input[39520]), .Z(n1067) );
  AND U1603 ( .A(n1069), .B(n1070), .Z(o[951]) );
  AND U1604 ( .A(p_input[20951]), .B(p_input[10951]), .Z(n1070) );
  AND U1605 ( .A(p_input[951]), .B(p_input[30951]), .Z(n1069) );
  AND U1606 ( .A(n1071), .B(n1072), .Z(o[9519]) );
  AND U1607 ( .A(p_input[29519]), .B(p_input[19519]), .Z(n1072) );
  AND U1608 ( .A(p_input[9519]), .B(p_input[39519]), .Z(n1071) );
  AND U1609 ( .A(n1073), .B(n1074), .Z(o[9518]) );
  AND U1610 ( .A(p_input[29518]), .B(p_input[19518]), .Z(n1074) );
  AND U1611 ( .A(p_input[9518]), .B(p_input[39518]), .Z(n1073) );
  AND U1612 ( .A(n1075), .B(n1076), .Z(o[9517]) );
  AND U1613 ( .A(p_input[29517]), .B(p_input[19517]), .Z(n1076) );
  AND U1614 ( .A(p_input[9517]), .B(p_input[39517]), .Z(n1075) );
  AND U1615 ( .A(n1077), .B(n1078), .Z(o[9516]) );
  AND U1616 ( .A(p_input[29516]), .B(p_input[19516]), .Z(n1078) );
  AND U1617 ( .A(p_input[9516]), .B(p_input[39516]), .Z(n1077) );
  AND U1618 ( .A(n1079), .B(n1080), .Z(o[9515]) );
  AND U1619 ( .A(p_input[29515]), .B(p_input[19515]), .Z(n1080) );
  AND U1620 ( .A(p_input[9515]), .B(p_input[39515]), .Z(n1079) );
  AND U1621 ( .A(n1081), .B(n1082), .Z(o[9514]) );
  AND U1622 ( .A(p_input[29514]), .B(p_input[19514]), .Z(n1082) );
  AND U1623 ( .A(p_input[9514]), .B(p_input[39514]), .Z(n1081) );
  AND U1624 ( .A(n1083), .B(n1084), .Z(o[9513]) );
  AND U1625 ( .A(p_input[29513]), .B(p_input[19513]), .Z(n1084) );
  AND U1626 ( .A(p_input[9513]), .B(p_input[39513]), .Z(n1083) );
  AND U1627 ( .A(n1085), .B(n1086), .Z(o[9512]) );
  AND U1628 ( .A(p_input[29512]), .B(p_input[19512]), .Z(n1086) );
  AND U1629 ( .A(p_input[9512]), .B(p_input[39512]), .Z(n1085) );
  AND U1630 ( .A(n1087), .B(n1088), .Z(o[9511]) );
  AND U1631 ( .A(p_input[29511]), .B(p_input[19511]), .Z(n1088) );
  AND U1632 ( .A(p_input[9511]), .B(p_input[39511]), .Z(n1087) );
  AND U1633 ( .A(n1089), .B(n1090), .Z(o[9510]) );
  AND U1634 ( .A(p_input[29510]), .B(p_input[19510]), .Z(n1090) );
  AND U1635 ( .A(p_input[9510]), .B(p_input[39510]), .Z(n1089) );
  AND U1636 ( .A(n1091), .B(n1092), .Z(o[950]) );
  AND U1637 ( .A(p_input[20950]), .B(p_input[10950]), .Z(n1092) );
  AND U1638 ( .A(p_input[950]), .B(p_input[30950]), .Z(n1091) );
  AND U1639 ( .A(n1093), .B(n1094), .Z(o[9509]) );
  AND U1640 ( .A(p_input[29509]), .B(p_input[19509]), .Z(n1094) );
  AND U1641 ( .A(p_input[9509]), .B(p_input[39509]), .Z(n1093) );
  AND U1642 ( .A(n1095), .B(n1096), .Z(o[9508]) );
  AND U1643 ( .A(p_input[29508]), .B(p_input[19508]), .Z(n1096) );
  AND U1644 ( .A(p_input[9508]), .B(p_input[39508]), .Z(n1095) );
  AND U1645 ( .A(n1097), .B(n1098), .Z(o[9507]) );
  AND U1646 ( .A(p_input[29507]), .B(p_input[19507]), .Z(n1098) );
  AND U1647 ( .A(p_input[9507]), .B(p_input[39507]), .Z(n1097) );
  AND U1648 ( .A(n1099), .B(n1100), .Z(o[9506]) );
  AND U1649 ( .A(p_input[29506]), .B(p_input[19506]), .Z(n1100) );
  AND U1650 ( .A(p_input[9506]), .B(p_input[39506]), .Z(n1099) );
  AND U1651 ( .A(n1101), .B(n1102), .Z(o[9505]) );
  AND U1652 ( .A(p_input[29505]), .B(p_input[19505]), .Z(n1102) );
  AND U1653 ( .A(p_input[9505]), .B(p_input[39505]), .Z(n1101) );
  AND U1654 ( .A(n1103), .B(n1104), .Z(o[9504]) );
  AND U1655 ( .A(p_input[29504]), .B(p_input[19504]), .Z(n1104) );
  AND U1656 ( .A(p_input[9504]), .B(p_input[39504]), .Z(n1103) );
  AND U1657 ( .A(n1105), .B(n1106), .Z(o[9503]) );
  AND U1658 ( .A(p_input[29503]), .B(p_input[19503]), .Z(n1106) );
  AND U1659 ( .A(p_input[9503]), .B(p_input[39503]), .Z(n1105) );
  AND U1660 ( .A(n1107), .B(n1108), .Z(o[9502]) );
  AND U1661 ( .A(p_input[29502]), .B(p_input[19502]), .Z(n1108) );
  AND U1662 ( .A(p_input[9502]), .B(p_input[39502]), .Z(n1107) );
  AND U1663 ( .A(n1109), .B(n1110), .Z(o[9501]) );
  AND U1664 ( .A(p_input[29501]), .B(p_input[19501]), .Z(n1110) );
  AND U1665 ( .A(p_input[9501]), .B(p_input[39501]), .Z(n1109) );
  AND U1666 ( .A(n1111), .B(n1112), .Z(o[9500]) );
  AND U1667 ( .A(p_input[29500]), .B(p_input[19500]), .Z(n1112) );
  AND U1668 ( .A(p_input[9500]), .B(p_input[39500]), .Z(n1111) );
  AND U1669 ( .A(n1113), .B(n1114), .Z(o[94]) );
  AND U1670 ( .A(p_input[20094]), .B(p_input[10094]), .Z(n1114) );
  AND U1671 ( .A(p_input[94]), .B(p_input[30094]), .Z(n1113) );
  AND U1672 ( .A(n1115), .B(n1116), .Z(o[949]) );
  AND U1673 ( .A(p_input[20949]), .B(p_input[10949]), .Z(n1116) );
  AND U1674 ( .A(p_input[949]), .B(p_input[30949]), .Z(n1115) );
  AND U1675 ( .A(n1117), .B(n1118), .Z(o[9499]) );
  AND U1676 ( .A(p_input[29499]), .B(p_input[19499]), .Z(n1118) );
  AND U1677 ( .A(p_input[9499]), .B(p_input[39499]), .Z(n1117) );
  AND U1678 ( .A(n1119), .B(n1120), .Z(o[9498]) );
  AND U1679 ( .A(p_input[29498]), .B(p_input[19498]), .Z(n1120) );
  AND U1680 ( .A(p_input[9498]), .B(p_input[39498]), .Z(n1119) );
  AND U1681 ( .A(n1121), .B(n1122), .Z(o[9497]) );
  AND U1682 ( .A(p_input[29497]), .B(p_input[19497]), .Z(n1122) );
  AND U1683 ( .A(p_input[9497]), .B(p_input[39497]), .Z(n1121) );
  AND U1684 ( .A(n1123), .B(n1124), .Z(o[9496]) );
  AND U1685 ( .A(p_input[29496]), .B(p_input[19496]), .Z(n1124) );
  AND U1686 ( .A(p_input[9496]), .B(p_input[39496]), .Z(n1123) );
  AND U1687 ( .A(n1125), .B(n1126), .Z(o[9495]) );
  AND U1688 ( .A(p_input[29495]), .B(p_input[19495]), .Z(n1126) );
  AND U1689 ( .A(p_input[9495]), .B(p_input[39495]), .Z(n1125) );
  AND U1690 ( .A(n1127), .B(n1128), .Z(o[9494]) );
  AND U1691 ( .A(p_input[29494]), .B(p_input[19494]), .Z(n1128) );
  AND U1692 ( .A(p_input[9494]), .B(p_input[39494]), .Z(n1127) );
  AND U1693 ( .A(n1129), .B(n1130), .Z(o[9493]) );
  AND U1694 ( .A(p_input[29493]), .B(p_input[19493]), .Z(n1130) );
  AND U1695 ( .A(p_input[9493]), .B(p_input[39493]), .Z(n1129) );
  AND U1696 ( .A(n1131), .B(n1132), .Z(o[9492]) );
  AND U1697 ( .A(p_input[29492]), .B(p_input[19492]), .Z(n1132) );
  AND U1698 ( .A(p_input[9492]), .B(p_input[39492]), .Z(n1131) );
  AND U1699 ( .A(n1133), .B(n1134), .Z(o[9491]) );
  AND U1700 ( .A(p_input[29491]), .B(p_input[19491]), .Z(n1134) );
  AND U1701 ( .A(p_input[9491]), .B(p_input[39491]), .Z(n1133) );
  AND U1702 ( .A(n1135), .B(n1136), .Z(o[9490]) );
  AND U1703 ( .A(p_input[29490]), .B(p_input[19490]), .Z(n1136) );
  AND U1704 ( .A(p_input[9490]), .B(p_input[39490]), .Z(n1135) );
  AND U1705 ( .A(n1137), .B(n1138), .Z(o[948]) );
  AND U1706 ( .A(p_input[20948]), .B(p_input[10948]), .Z(n1138) );
  AND U1707 ( .A(p_input[948]), .B(p_input[30948]), .Z(n1137) );
  AND U1708 ( .A(n1139), .B(n1140), .Z(o[9489]) );
  AND U1709 ( .A(p_input[29489]), .B(p_input[19489]), .Z(n1140) );
  AND U1710 ( .A(p_input[9489]), .B(p_input[39489]), .Z(n1139) );
  AND U1711 ( .A(n1141), .B(n1142), .Z(o[9488]) );
  AND U1712 ( .A(p_input[29488]), .B(p_input[19488]), .Z(n1142) );
  AND U1713 ( .A(p_input[9488]), .B(p_input[39488]), .Z(n1141) );
  AND U1714 ( .A(n1143), .B(n1144), .Z(o[9487]) );
  AND U1715 ( .A(p_input[29487]), .B(p_input[19487]), .Z(n1144) );
  AND U1716 ( .A(p_input[9487]), .B(p_input[39487]), .Z(n1143) );
  AND U1717 ( .A(n1145), .B(n1146), .Z(o[9486]) );
  AND U1718 ( .A(p_input[29486]), .B(p_input[19486]), .Z(n1146) );
  AND U1719 ( .A(p_input[9486]), .B(p_input[39486]), .Z(n1145) );
  AND U1720 ( .A(n1147), .B(n1148), .Z(o[9485]) );
  AND U1721 ( .A(p_input[29485]), .B(p_input[19485]), .Z(n1148) );
  AND U1722 ( .A(p_input[9485]), .B(p_input[39485]), .Z(n1147) );
  AND U1723 ( .A(n1149), .B(n1150), .Z(o[9484]) );
  AND U1724 ( .A(p_input[29484]), .B(p_input[19484]), .Z(n1150) );
  AND U1725 ( .A(p_input[9484]), .B(p_input[39484]), .Z(n1149) );
  AND U1726 ( .A(n1151), .B(n1152), .Z(o[9483]) );
  AND U1727 ( .A(p_input[29483]), .B(p_input[19483]), .Z(n1152) );
  AND U1728 ( .A(p_input[9483]), .B(p_input[39483]), .Z(n1151) );
  AND U1729 ( .A(n1153), .B(n1154), .Z(o[9482]) );
  AND U1730 ( .A(p_input[29482]), .B(p_input[19482]), .Z(n1154) );
  AND U1731 ( .A(p_input[9482]), .B(p_input[39482]), .Z(n1153) );
  AND U1732 ( .A(n1155), .B(n1156), .Z(o[9481]) );
  AND U1733 ( .A(p_input[29481]), .B(p_input[19481]), .Z(n1156) );
  AND U1734 ( .A(p_input[9481]), .B(p_input[39481]), .Z(n1155) );
  AND U1735 ( .A(n1157), .B(n1158), .Z(o[9480]) );
  AND U1736 ( .A(p_input[29480]), .B(p_input[19480]), .Z(n1158) );
  AND U1737 ( .A(p_input[9480]), .B(p_input[39480]), .Z(n1157) );
  AND U1738 ( .A(n1159), .B(n1160), .Z(o[947]) );
  AND U1739 ( .A(p_input[20947]), .B(p_input[10947]), .Z(n1160) );
  AND U1740 ( .A(p_input[947]), .B(p_input[30947]), .Z(n1159) );
  AND U1741 ( .A(n1161), .B(n1162), .Z(o[9479]) );
  AND U1742 ( .A(p_input[29479]), .B(p_input[19479]), .Z(n1162) );
  AND U1743 ( .A(p_input[9479]), .B(p_input[39479]), .Z(n1161) );
  AND U1744 ( .A(n1163), .B(n1164), .Z(o[9478]) );
  AND U1745 ( .A(p_input[29478]), .B(p_input[19478]), .Z(n1164) );
  AND U1746 ( .A(p_input[9478]), .B(p_input[39478]), .Z(n1163) );
  AND U1747 ( .A(n1165), .B(n1166), .Z(o[9477]) );
  AND U1748 ( .A(p_input[29477]), .B(p_input[19477]), .Z(n1166) );
  AND U1749 ( .A(p_input[9477]), .B(p_input[39477]), .Z(n1165) );
  AND U1750 ( .A(n1167), .B(n1168), .Z(o[9476]) );
  AND U1751 ( .A(p_input[29476]), .B(p_input[19476]), .Z(n1168) );
  AND U1752 ( .A(p_input[9476]), .B(p_input[39476]), .Z(n1167) );
  AND U1753 ( .A(n1169), .B(n1170), .Z(o[9475]) );
  AND U1754 ( .A(p_input[29475]), .B(p_input[19475]), .Z(n1170) );
  AND U1755 ( .A(p_input[9475]), .B(p_input[39475]), .Z(n1169) );
  AND U1756 ( .A(n1171), .B(n1172), .Z(o[9474]) );
  AND U1757 ( .A(p_input[29474]), .B(p_input[19474]), .Z(n1172) );
  AND U1758 ( .A(p_input[9474]), .B(p_input[39474]), .Z(n1171) );
  AND U1759 ( .A(n1173), .B(n1174), .Z(o[9473]) );
  AND U1760 ( .A(p_input[29473]), .B(p_input[19473]), .Z(n1174) );
  AND U1761 ( .A(p_input[9473]), .B(p_input[39473]), .Z(n1173) );
  AND U1762 ( .A(n1175), .B(n1176), .Z(o[9472]) );
  AND U1763 ( .A(p_input[29472]), .B(p_input[19472]), .Z(n1176) );
  AND U1764 ( .A(p_input[9472]), .B(p_input[39472]), .Z(n1175) );
  AND U1765 ( .A(n1177), .B(n1178), .Z(o[9471]) );
  AND U1766 ( .A(p_input[29471]), .B(p_input[19471]), .Z(n1178) );
  AND U1767 ( .A(p_input[9471]), .B(p_input[39471]), .Z(n1177) );
  AND U1768 ( .A(n1179), .B(n1180), .Z(o[9470]) );
  AND U1769 ( .A(p_input[29470]), .B(p_input[19470]), .Z(n1180) );
  AND U1770 ( .A(p_input[9470]), .B(p_input[39470]), .Z(n1179) );
  AND U1771 ( .A(n1181), .B(n1182), .Z(o[946]) );
  AND U1772 ( .A(p_input[20946]), .B(p_input[10946]), .Z(n1182) );
  AND U1773 ( .A(p_input[946]), .B(p_input[30946]), .Z(n1181) );
  AND U1774 ( .A(n1183), .B(n1184), .Z(o[9469]) );
  AND U1775 ( .A(p_input[29469]), .B(p_input[19469]), .Z(n1184) );
  AND U1776 ( .A(p_input[9469]), .B(p_input[39469]), .Z(n1183) );
  AND U1777 ( .A(n1185), .B(n1186), .Z(o[9468]) );
  AND U1778 ( .A(p_input[29468]), .B(p_input[19468]), .Z(n1186) );
  AND U1779 ( .A(p_input[9468]), .B(p_input[39468]), .Z(n1185) );
  AND U1780 ( .A(n1187), .B(n1188), .Z(o[9467]) );
  AND U1781 ( .A(p_input[29467]), .B(p_input[19467]), .Z(n1188) );
  AND U1782 ( .A(p_input[9467]), .B(p_input[39467]), .Z(n1187) );
  AND U1783 ( .A(n1189), .B(n1190), .Z(o[9466]) );
  AND U1784 ( .A(p_input[29466]), .B(p_input[19466]), .Z(n1190) );
  AND U1785 ( .A(p_input[9466]), .B(p_input[39466]), .Z(n1189) );
  AND U1786 ( .A(n1191), .B(n1192), .Z(o[9465]) );
  AND U1787 ( .A(p_input[29465]), .B(p_input[19465]), .Z(n1192) );
  AND U1788 ( .A(p_input[9465]), .B(p_input[39465]), .Z(n1191) );
  AND U1789 ( .A(n1193), .B(n1194), .Z(o[9464]) );
  AND U1790 ( .A(p_input[29464]), .B(p_input[19464]), .Z(n1194) );
  AND U1791 ( .A(p_input[9464]), .B(p_input[39464]), .Z(n1193) );
  AND U1792 ( .A(n1195), .B(n1196), .Z(o[9463]) );
  AND U1793 ( .A(p_input[29463]), .B(p_input[19463]), .Z(n1196) );
  AND U1794 ( .A(p_input[9463]), .B(p_input[39463]), .Z(n1195) );
  AND U1795 ( .A(n1197), .B(n1198), .Z(o[9462]) );
  AND U1796 ( .A(p_input[29462]), .B(p_input[19462]), .Z(n1198) );
  AND U1797 ( .A(p_input[9462]), .B(p_input[39462]), .Z(n1197) );
  AND U1798 ( .A(n1199), .B(n1200), .Z(o[9461]) );
  AND U1799 ( .A(p_input[29461]), .B(p_input[19461]), .Z(n1200) );
  AND U1800 ( .A(p_input[9461]), .B(p_input[39461]), .Z(n1199) );
  AND U1801 ( .A(n1201), .B(n1202), .Z(o[9460]) );
  AND U1802 ( .A(p_input[29460]), .B(p_input[19460]), .Z(n1202) );
  AND U1803 ( .A(p_input[9460]), .B(p_input[39460]), .Z(n1201) );
  AND U1804 ( .A(n1203), .B(n1204), .Z(o[945]) );
  AND U1805 ( .A(p_input[20945]), .B(p_input[10945]), .Z(n1204) );
  AND U1806 ( .A(p_input[945]), .B(p_input[30945]), .Z(n1203) );
  AND U1807 ( .A(n1205), .B(n1206), .Z(o[9459]) );
  AND U1808 ( .A(p_input[29459]), .B(p_input[19459]), .Z(n1206) );
  AND U1809 ( .A(p_input[9459]), .B(p_input[39459]), .Z(n1205) );
  AND U1810 ( .A(n1207), .B(n1208), .Z(o[9458]) );
  AND U1811 ( .A(p_input[29458]), .B(p_input[19458]), .Z(n1208) );
  AND U1812 ( .A(p_input[9458]), .B(p_input[39458]), .Z(n1207) );
  AND U1813 ( .A(n1209), .B(n1210), .Z(o[9457]) );
  AND U1814 ( .A(p_input[29457]), .B(p_input[19457]), .Z(n1210) );
  AND U1815 ( .A(p_input[9457]), .B(p_input[39457]), .Z(n1209) );
  AND U1816 ( .A(n1211), .B(n1212), .Z(o[9456]) );
  AND U1817 ( .A(p_input[29456]), .B(p_input[19456]), .Z(n1212) );
  AND U1818 ( .A(p_input[9456]), .B(p_input[39456]), .Z(n1211) );
  AND U1819 ( .A(n1213), .B(n1214), .Z(o[9455]) );
  AND U1820 ( .A(p_input[29455]), .B(p_input[19455]), .Z(n1214) );
  AND U1821 ( .A(p_input[9455]), .B(p_input[39455]), .Z(n1213) );
  AND U1822 ( .A(n1215), .B(n1216), .Z(o[9454]) );
  AND U1823 ( .A(p_input[29454]), .B(p_input[19454]), .Z(n1216) );
  AND U1824 ( .A(p_input[9454]), .B(p_input[39454]), .Z(n1215) );
  AND U1825 ( .A(n1217), .B(n1218), .Z(o[9453]) );
  AND U1826 ( .A(p_input[29453]), .B(p_input[19453]), .Z(n1218) );
  AND U1827 ( .A(p_input[9453]), .B(p_input[39453]), .Z(n1217) );
  AND U1828 ( .A(n1219), .B(n1220), .Z(o[9452]) );
  AND U1829 ( .A(p_input[29452]), .B(p_input[19452]), .Z(n1220) );
  AND U1830 ( .A(p_input[9452]), .B(p_input[39452]), .Z(n1219) );
  AND U1831 ( .A(n1221), .B(n1222), .Z(o[9451]) );
  AND U1832 ( .A(p_input[29451]), .B(p_input[19451]), .Z(n1222) );
  AND U1833 ( .A(p_input[9451]), .B(p_input[39451]), .Z(n1221) );
  AND U1834 ( .A(n1223), .B(n1224), .Z(o[9450]) );
  AND U1835 ( .A(p_input[29450]), .B(p_input[19450]), .Z(n1224) );
  AND U1836 ( .A(p_input[9450]), .B(p_input[39450]), .Z(n1223) );
  AND U1837 ( .A(n1225), .B(n1226), .Z(o[944]) );
  AND U1838 ( .A(p_input[20944]), .B(p_input[10944]), .Z(n1226) );
  AND U1839 ( .A(p_input[944]), .B(p_input[30944]), .Z(n1225) );
  AND U1840 ( .A(n1227), .B(n1228), .Z(o[9449]) );
  AND U1841 ( .A(p_input[29449]), .B(p_input[19449]), .Z(n1228) );
  AND U1842 ( .A(p_input[9449]), .B(p_input[39449]), .Z(n1227) );
  AND U1843 ( .A(n1229), .B(n1230), .Z(o[9448]) );
  AND U1844 ( .A(p_input[29448]), .B(p_input[19448]), .Z(n1230) );
  AND U1845 ( .A(p_input[9448]), .B(p_input[39448]), .Z(n1229) );
  AND U1846 ( .A(n1231), .B(n1232), .Z(o[9447]) );
  AND U1847 ( .A(p_input[29447]), .B(p_input[19447]), .Z(n1232) );
  AND U1848 ( .A(p_input[9447]), .B(p_input[39447]), .Z(n1231) );
  AND U1849 ( .A(n1233), .B(n1234), .Z(o[9446]) );
  AND U1850 ( .A(p_input[29446]), .B(p_input[19446]), .Z(n1234) );
  AND U1851 ( .A(p_input[9446]), .B(p_input[39446]), .Z(n1233) );
  AND U1852 ( .A(n1235), .B(n1236), .Z(o[9445]) );
  AND U1853 ( .A(p_input[29445]), .B(p_input[19445]), .Z(n1236) );
  AND U1854 ( .A(p_input[9445]), .B(p_input[39445]), .Z(n1235) );
  AND U1855 ( .A(n1237), .B(n1238), .Z(o[9444]) );
  AND U1856 ( .A(p_input[29444]), .B(p_input[19444]), .Z(n1238) );
  AND U1857 ( .A(p_input[9444]), .B(p_input[39444]), .Z(n1237) );
  AND U1858 ( .A(n1239), .B(n1240), .Z(o[9443]) );
  AND U1859 ( .A(p_input[29443]), .B(p_input[19443]), .Z(n1240) );
  AND U1860 ( .A(p_input[9443]), .B(p_input[39443]), .Z(n1239) );
  AND U1861 ( .A(n1241), .B(n1242), .Z(o[9442]) );
  AND U1862 ( .A(p_input[29442]), .B(p_input[19442]), .Z(n1242) );
  AND U1863 ( .A(p_input[9442]), .B(p_input[39442]), .Z(n1241) );
  AND U1864 ( .A(n1243), .B(n1244), .Z(o[9441]) );
  AND U1865 ( .A(p_input[29441]), .B(p_input[19441]), .Z(n1244) );
  AND U1866 ( .A(p_input[9441]), .B(p_input[39441]), .Z(n1243) );
  AND U1867 ( .A(n1245), .B(n1246), .Z(o[9440]) );
  AND U1868 ( .A(p_input[29440]), .B(p_input[19440]), .Z(n1246) );
  AND U1869 ( .A(p_input[9440]), .B(p_input[39440]), .Z(n1245) );
  AND U1870 ( .A(n1247), .B(n1248), .Z(o[943]) );
  AND U1871 ( .A(p_input[20943]), .B(p_input[10943]), .Z(n1248) );
  AND U1872 ( .A(p_input[943]), .B(p_input[30943]), .Z(n1247) );
  AND U1873 ( .A(n1249), .B(n1250), .Z(o[9439]) );
  AND U1874 ( .A(p_input[29439]), .B(p_input[19439]), .Z(n1250) );
  AND U1875 ( .A(p_input[9439]), .B(p_input[39439]), .Z(n1249) );
  AND U1876 ( .A(n1251), .B(n1252), .Z(o[9438]) );
  AND U1877 ( .A(p_input[29438]), .B(p_input[19438]), .Z(n1252) );
  AND U1878 ( .A(p_input[9438]), .B(p_input[39438]), .Z(n1251) );
  AND U1879 ( .A(n1253), .B(n1254), .Z(o[9437]) );
  AND U1880 ( .A(p_input[29437]), .B(p_input[19437]), .Z(n1254) );
  AND U1881 ( .A(p_input[9437]), .B(p_input[39437]), .Z(n1253) );
  AND U1882 ( .A(n1255), .B(n1256), .Z(o[9436]) );
  AND U1883 ( .A(p_input[29436]), .B(p_input[19436]), .Z(n1256) );
  AND U1884 ( .A(p_input[9436]), .B(p_input[39436]), .Z(n1255) );
  AND U1885 ( .A(n1257), .B(n1258), .Z(o[9435]) );
  AND U1886 ( .A(p_input[29435]), .B(p_input[19435]), .Z(n1258) );
  AND U1887 ( .A(p_input[9435]), .B(p_input[39435]), .Z(n1257) );
  AND U1888 ( .A(n1259), .B(n1260), .Z(o[9434]) );
  AND U1889 ( .A(p_input[29434]), .B(p_input[19434]), .Z(n1260) );
  AND U1890 ( .A(p_input[9434]), .B(p_input[39434]), .Z(n1259) );
  AND U1891 ( .A(n1261), .B(n1262), .Z(o[9433]) );
  AND U1892 ( .A(p_input[29433]), .B(p_input[19433]), .Z(n1262) );
  AND U1893 ( .A(p_input[9433]), .B(p_input[39433]), .Z(n1261) );
  AND U1894 ( .A(n1263), .B(n1264), .Z(o[9432]) );
  AND U1895 ( .A(p_input[29432]), .B(p_input[19432]), .Z(n1264) );
  AND U1896 ( .A(p_input[9432]), .B(p_input[39432]), .Z(n1263) );
  AND U1897 ( .A(n1265), .B(n1266), .Z(o[9431]) );
  AND U1898 ( .A(p_input[29431]), .B(p_input[19431]), .Z(n1266) );
  AND U1899 ( .A(p_input[9431]), .B(p_input[39431]), .Z(n1265) );
  AND U1900 ( .A(n1267), .B(n1268), .Z(o[9430]) );
  AND U1901 ( .A(p_input[29430]), .B(p_input[19430]), .Z(n1268) );
  AND U1902 ( .A(p_input[9430]), .B(p_input[39430]), .Z(n1267) );
  AND U1903 ( .A(n1269), .B(n1270), .Z(o[942]) );
  AND U1904 ( .A(p_input[20942]), .B(p_input[10942]), .Z(n1270) );
  AND U1905 ( .A(p_input[942]), .B(p_input[30942]), .Z(n1269) );
  AND U1906 ( .A(n1271), .B(n1272), .Z(o[9429]) );
  AND U1907 ( .A(p_input[29429]), .B(p_input[19429]), .Z(n1272) );
  AND U1908 ( .A(p_input[9429]), .B(p_input[39429]), .Z(n1271) );
  AND U1909 ( .A(n1273), .B(n1274), .Z(o[9428]) );
  AND U1910 ( .A(p_input[29428]), .B(p_input[19428]), .Z(n1274) );
  AND U1911 ( .A(p_input[9428]), .B(p_input[39428]), .Z(n1273) );
  AND U1912 ( .A(n1275), .B(n1276), .Z(o[9427]) );
  AND U1913 ( .A(p_input[29427]), .B(p_input[19427]), .Z(n1276) );
  AND U1914 ( .A(p_input[9427]), .B(p_input[39427]), .Z(n1275) );
  AND U1915 ( .A(n1277), .B(n1278), .Z(o[9426]) );
  AND U1916 ( .A(p_input[29426]), .B(p_input[19426]), .Z(n1278) );
  AND U1917 ( .A(p_input[9426]), .B(p_input[39426]), .Z(n1277) );
  AND U1918 ( .A(n1279), .B(n1280), .Z(o[9425]) );
  AND U1919 ( .A(p_input[29425]), .B(p_input[19425]), .Z(n1280) );
  AND U1920 ( .A(p_input[9425]), .B(p_input[39425]), .Z(n1279) );
  AND U1921 ( .A(n1281), .B(n1282), .Z(o[9424]) );
  AND U1922 ( .A(p_input[29424]), .B(p_input[19424]), .Z(n1282) );
  AND U1923 ( .A(p_input[9424]), .B(p_input[39424]), .Z(n1281) );
  AND U1924 ( .A(n1283), .B(n1284), .Z(o[9423]) );
  AND U1925 ( .A(p_input[29423]), .B(p_input[19423]), .Z(n1284) );
  AND U1926 ( .A(p_input[9423]), .B(p_input[39423]), .Z(n1283) );
  AND U1927 ( .A(n1285), .B(n1286), .Z(o[9422]) );
  AND U1928 ( .A(p_input[29422]), .B(p_input[19422]), .Z(n1286) );
  AND U1929 ( .A(p_input[9422]), .B(p_input[39422]), .Z(n1285) );
  AND U1930 ( .A(n1287), .B(n1288), .Z(o[9421]) );
  AND U1931 ( .A(p_input[29421]), .B(p_input[19421]), .Z(n1288) );
  AND U1932 ( .A(p_input[9421]), .B(p_input[39421]), .Z(n1287) );
  AND U1933 ( .A(n1289), .B(n1290), .Z(o[9420]) );
  AND U1934 ( .A(p_input[29420]), .B(p_input[19420]), .Z(n1290) );
  AND U1935 ( .A(p_input[9420]), .B(p_input[39420]), .Z(n1289) );
  AND U1936 ( .A(n1291), .B(n1292), .Z(o[941]) );
  AND U1937 ( .A(p_input[20941]), .B(p_input[10941]), .Z(n1292) );
  AND U1938 ( .A(p_input[941]), .B(p_input[30941]), .Z(n1291) );
  AND U1939 ( .A(n1293), .B(n1294), .Z(o[9419]) );
  AND U1940 ( .A(p_input[29419]), .B(p_input[19419]), .Z(n1294) );
  AND U1941 ( .A(p_input[9419]), .B(p_input[39419]), .Z(n1293) );
  AND U1942 ( .A(n1295), .B(n1296), .Z(o[9418]) );
  AND U1943 ( .A(p_input[29418]), .B(p_input[19418]), .Z(n1296) );
  AND U1944 ( .A(p_input[9418]), .B(p_input[39418]), .Z(n1295) );
  AND U1945 ( .A(n1297), .B(n1298), .Z(o[9417]) );
  AND U1946 ( .A(p_input[29417]), .B(p_input[19417]), .Z(n1298) );
  AND U1947 ( .A(p_input[9417]), .B(p_input[39417]), .Z(n1297) );
  AND U1948 ( .A(n1299), .B(n1300), .Z(o[9416]) );
  AND U1949 ( .A(p_input[29416]), .B(p_input[19416]), .Z(n1300) );
  AND U1950 ( .A(p_input[9416]), .B(p_input[39416]), .Z(n1299) );
  AND U1951 ( .A(n1301), .B(n1302), .Z(o[9415]) );
  AND U1952 ( .A(p_input[29415]), .B(p_input[19415]), .Z(n1302) );
  AND U1953 ( .A(p_input[9415]), .B(p_input[39415]), .Z(n1301) );
  AND U1954 ( .A(n1303), .B(n1304), .Z(o[9414]) );
  AND U1955 ( .A(p_input[29414]), .B(p_input[19414]), .Z(n1304) );
  AND U1956 ( .A(p_input[9414]), .B(p_input[39414]), .Z(n1303) );
  AND U1957 ( .A(n1305), .B(n1306), .Z(o[9413]) );
  AND U1958 ( .A(p_input[29413]), .B(p_input[19413]), .Z(n1306) );
  AND U1959 ( .A(p_input[9413]), .B(p_input[39413]), .Z(n1305) );
  AND U1960 ( .A(n1307), .B(n1308), .Z(o[9412]) );
  AND U1961 ( .A(p_input[29412]), .B(p_input[19412]), .Z(n1308) );
  AND U1962 ( .A(p_input[9412]), .B(p_input[39412]), .Z(n1307) );
  AND U1963 ( .A(n1309), .B(n1310), .Z(o[9411]) );
  AND U1964 ( .A(p_input[29411]), .B(p_input[19411]), .Z(n1310) );
  AND U1965 ( .A(p_input[9411]), .B(p_input[39411]), .Z(n1309) );
  AND U1966 ( .A(n1311), .B(n1312), .Z(o[9410]) );
  AND U1967 ( .A(p_input[29410]), .B(p_input[19410]), .Z(n1312) );
  AND U1968 ( .A(p_input[9410]), .B(p_input[39410]), .Z(n1311) );
  AND U1969 ( .A(n1313), .B(n1314), .Z(o[940]) );
  AND U1970 ( .A(p_input[20940]), .B(p_input[10940]), .Z(n1314) );
  AND U1971 ( .A(p_input[940]), .B(p_input[30940]), .Z(n1313) );
  AND U1972 ( .A(n1315), .B(n1316), .Z(o[9409]) );
  AND U1973 ( .A(p_input[29409]), .B(p_input[19409]), .Z(n1316) );
  AND U1974 ( .A(p_input[9409]), .B(p_input[39409]), .Z(n1315) );
  AND U1975 ( .A(n1317), .B(n1318), .Z(o[9408]) );
  AND U1976 ( .A(p_input[29408]), .B(p_input[19408]), .Z(n1318) );
  AND U1977 ( .A(p_input[9408]), .B(p_input[39408]), .Z(n1317) );
  AND U1978 ( .A(n1319), .B(n1320), .Z(o[9407]) );
  AND U1979 ( .A(p_input[29407]), .B(p_input[19407]), .Z(n1320) );
  AND U1980 ( .A(p_input[9407]), .B(p_input[39407]), .Z(n1319) );
  AND U1981 ( .A(n1321), .B(n1322), .Z(o[9406]) );
  AND U1982 ( .A(p_input[29406]), .B(p_input[19406]), .Z(n1322) );
  AND U1983 ( .A(p_input[9406]), .B(p_input[39406]), .Z(n1321) );
  AND U1984 ( .A(n1323), .B(n1324), .Z(o[9405]) );
  AND U1985 ( .A(p_input[29405]), .B(p_input[19405]), .Z(n1324) );
  AND U1986 ( .A(p_input[9405]), .B(p_input[39405]), .Z(n1323) );
  AND U1987 ( .A(n1325), .B(n1326), .Z(o[9404]) );
  AND U1988 ( .A(p_input[29404]), .B(p_input[19404]), .Z(n1326) );
  AND U1989 ( .A(p_input[9404]), .B(p_input[39404]), .Z(n1325) );
  AND U1990 ( .A(n1327), .B(n1328), .Z(o[9403]) );
  AND U1991 ( .A(p_input[29403]), .B(p_input[19403]), .Z(n1328) );
  AND U1992 ( .A(p_input[9403]), .B(p_input[39403]), .Z(n1327) );
  AND U1993 ( .A(n1329), .B(n1330), .Z(o[9402]) );
  AND U1994 ( .A(p_input[29402]), .B(p_input[19402]), .Z(n1330) );
  AND U1995 ( .A(p_input[9402]), .B(p_input[39402]), .Z(n1329) );
  AND U1996 ( .A(n1331), .B(n1332), .Z(o[9401]) );
  AND U1997 ( .A(p_input[29401]), .B(p_input[19401]), .Z(n1332) );
  AND U1998 ( .A(p_input[9401]), .B(p_input[39401]), .Z(n1331) );
  AND U1999 ( .A(n1333), .B(n1334), .Z(o[9400]) );
  AND U2000 ( .A(p_input[29400]), .B(p_input[19400]), .Z(n1334) );
  AND U2001 ( .A(p_input[9400]), .B(p_input[39400]), .Z(n1333) );
  AND U2002 ( .A(n1335), .B(n1336), .Z(o[93]) );
  AND U2003 ( .A(p_input[20093]), .B(p_input[10093]), .Z(n1336) );
  AND U2004 ( .A(p_input[93]), .B(p_input[30093]), .Z(n1335) );
  AND U2005 ( .A(n1337), .B(n1338), .Z(o[939]) );
  AND U2006 ( .A(p_input[20939]), .B(p_input[10939]), .Z(n1338) );
  AND U2007 ( .A(p_input[939]), .B(p_input[30939]), .Z(n1337) );
  AND U2008 ( .A(n1339), .B(n1340), .Z(o[9399]) );
  AND U2009 ( .A(p_input[29399]), .B(p_input[19399]), .Z(n1340) );
  AND U2010 ( .A(p_input[9399]), .B(p_input[39399]), .Z(n1339) );
  AND U2011 ( .A(n1341), .B(n1342), .Z(o[9398]) );
  AND U2012 ( .A(p_input[29398]), .B(p_input[19398]), .Z(n1342) );
  AND U2013 ( .A(p_input[9398]), .B(p_input[39398]), .Z(n1341) );
  AND U2014 ( .A(n1343), .B(n1344), .Z(o[9397]) );
  AND U2015 ( .A(p_input[29397]), .B(p_input[19397]), .Z(n1344) );
  AND U2016 ( .A(p_input[9397]), .B(p_input[39397]), .Z(n1343) );
  AND U2017 ( .A(n1345), .B(n1346), .Z(o[9396]) );
  AND U2018 ( .A(p_input[29396]), .B(p_input[19396]), .Z(n1346) );
  AND U2019 ( .A(p_input[9396]), .B(p_input[39396]), .Z(n1345) );
  AND U2020 ( .A(n1347), .B(n1348), .Z(o[9395]) );
  AND U2021 ( .A(p_input[29395]), .B(p_input[19395]), .Z(n1348) );
  AND U2022 ( .A(p_input[9395]), .B(p_input[39395]), .Z(n1347) );
  AND U2023 ( .A(n1349), .B(n1350), .Z(o[9394]) );
  AND U2024 ( .A(p_input[29394]), .B(p_input[19394]), .Z(n1350) );
  AND U2025 ( .A(p_input[9394]), .B(p_input[39394]), .Z(n1349) );
  AND U2026 ( .A(n1351), .B(n1352), .Z(o[9393]) );
  AND U2027 ( .A(p_input[29393]), .B(p_input[19393]), .Z(n1352) );
  AND U2028 ( .A(p_input[9393]), .B(p_input[39393]), .Z(n1351) );
  AND U2029 ( .A(n1353), .B(n1354), .Z(o[9392]) );
  AND U2030 ( .A(p_input[29392]), .B(p_input[19392]), .Z(n1354) );
  AND U2031 ( .A(p_input[9392]), .B(p_input[39392]), .Z(n1353) );
  AND U2032 ( .A(n1355), .B(n1356), .Z(o[9391]) );
  AND U2033 ( .A(p_input[29391]), .B(p_input[19391]), .Z(n1356) );
  AND U2034 ( .A(p_input[9391]), .B(p_input[39391]), .Z(n1355) );
  AND U2035 ( .A(n1357), .B(n1358), .Z(o[9390]) );
  AND U2036 ( .A(p_input[29390]), .B(p_input[19390]), .Z(n1358) );
  AND U2037 ( .A(p_input[9390]), .B(p_input[39390]), .Z(n1357) );
  AND U2038 ( .A(n1359), .B(n1360), .Z(o[938]) );
  AND U2039 ( .A(p_input[20938]), .B(p_input[10938]), .Z(n1360) );
  AND U2040 ( .A(p_input[938]), .B(p_input[30938]), .Z(n1359) );
  AND U2041 ( .A(n1361), .B(n1362), .Z(o[9389]) );
  AND U2042 ( .A(p_input[29389]), .B(p_input[19389]), .Z(n1362) );
  AND U2043 ( .A(p_input[9389]), .B(p_input[39389]), .Z(n1361) );
  AND U2044 ( .A(n1363), .B(n1364), .Z(o[9388]) );
  AND U2045 ( .A(p_input[29388]), .B(p_input[19388]), .Z(n1364) );
  AND U2046 ( .A(p_input[9388]), .B(p_input[39388]), .Z(n1363) );
  AND U2047 ( .A(n1365), .B(n1366), .Z(o[9387]) );
  AND U2048 ( .A(p_input[29387]), .B(p_input[19387]), .Z(n1366) );
  AND U2049 ( .A(p_input[9387]), .B(p_input[39387]), .Z(n1365) );
  AND U2050 ( .A(n1367), .B(n1368), .Z(o[9386]) );
  AND U2051 ( .A(p_input[29386]), .B(p_input[19386]), .Z(n1368) );
  AND U2052 ( .A(p_input[9386]), .B(p_input[39386]), .Z(n1367) );
  AND U2053 ( .A(n1369), .B(n1370), .Z(o[9385]) );
  AND U2054 ( .A(p_input[29385]), .B(p_input[19385]), .Z(n1370) );
  AND U2055 ( .A(p_input[9385]), .B(p_input[39385]), .Z(n1369) );
  AND U2056 ( .A(n1371), .B(n1372), .Z(o[9384]) );
  AND U2057 ( .A(p_input[29384]), .B(p_input[19384]), .Z(n1372) );
  AND U2058 ( .A(p_input[9384]), .B(p_input[39384]), .Z(n1371) );
  AND U2059 ( .A(n1373), .B(n1374), .Z(o[9383]) );
  AND U2060 ( .A(p_input[29383]), .B(p_input[19383]), .Z(n1374) );
  AND U2061 ( .A(p_input[9383]), .B(p_input[39383]), .Z(n1373) );
  AND U2062 ( .A(n1375), .B(n1376), .Z(o[9382]) );
  AND U2063 ( .A(p_input[29382]), .B(p_input[19382]), .Z(n1376) );
  AND U2064 ( .A(p_input[9382]), .B(p_input[39382]), .Z(n1375) );
  AND U2065 ( .A(n1377), .B(n1378), .Z(o[9381]) );
  AND U2066 ( .A(p_input[29381]), .B(p_input[19381]), .Z(n1378) );
  AND U2067 ( .A(p_input[9381]), .B(p_input[39381]), .Z(n1377) );
  AND U2068 ( .A(n1379), .B(n1380), .Z(o[9380]) );
  AND U2069 ( .A(p_input[29380]), .B(p_input[19380]), .Z(n1380) );
  AND U2070 ( .A(p_input[9380]), .B(p_input[39380]), .Z(n1379) );
  AND U2071 ( .A(n1381), .B(n1382), .Z(o[937]) );
  AND U2072 ( .A(p_input[20937]), .B(p_input[10937]), .Z(n1382) );
  AND U2073 ( .A(p_input[937]), .B(p_input[30937]), .Z(n1381) );
  AND U2074 ( .A(n1383), .B(n1384), .Z(o[9379]) );
  AND U2075 ( .A(p_input[29379]), .B(p_input[19379]), .Z(n1384) );
  AND U2076 ( .A(p_input[9379]), .B(p_input[39379]), .Z(n1383) );
  AND U2077 ( .A(n1385), .B(n1386), .Z(o[9378]) );
  AND U2078 ( .A(p_input[29378]), .B(p_input[19378]), .Z(n1386) );
  AND U2079 ( .A(p_input[9378]), .B(p_input[39378]), .Z(n1385) );
  AND U2080 ( .A(n1387), .B(n1388), .Z(o[9377]) );
  AND U2081 ( .A(p_input[29377]), .B(p_input[19377]), .Z(n1388) );
  AND U2082 ( .A(p_input[9377]), .B(p_input[39377]), .Z(n1387) );
  AND U2083 ( .A(n1389), .B(n1390), .Z(o[9376]) );
  AND U2084 ( .A(p_input[29376]), .B(p_input[19376]), .Z(n1390) );
  AND U2085 ( .A(p_input[9376]), .B(p_input[39376]), .Z(n1389) );
  AND U2086 ( .A(n1391), .B(n1392), .Z(o[9375]) );
  AND U2087 ( .A(p_input[29375]), .B(p_input[19375]), .Z(n1392) );
  AND U2088 ( .A(p_input[9375]), .B(p_input[39375]), .Z(n1391) );
  AND U2089 ( .A(n1393), .B(n1394), .Z(o[9374]) );
  AND U2090 ( .A(p_input[29374]), .B(p_input[19374]), .Z(n1394) );
  AND U2091 ( .A(p_input[9374]), .B(p_input[39374]), .Z(n1393) );
  AND U2092 ( .A(n1395), .B(n1396), .Z(o[9373]) );
  AND U2093 ( .A(p_input[29373]), .B(p_input[19373]), .Z(n1396) );
  AND U2094 ( .A(p_input[9373]), .B(p_input[39373]), .Z(n1395) );
  AND U2095 ( .A(n1397), .B(n1398), .Z(o[9372]) );
  AND U2096 ( .A(p_input[29372]), .B(p_input[19372]), .Z(n1398) );
  AND U2097 ( .A(p_input[9372]), .B(p_input[39372]), .Z(n1397) );
  AND U2098 ( .A(n1399), .B(n1400), .Z(o[9371]) );
  AND U2099 ( .A(p_input[29371]), .B(p_input[19371]), .Z(n1400) );
  AND U2100 ( .A(p_input[9371]), .B(p_input[39371]), .Z(n1399) );
  AND U2101 ( .A(n1401), .B(n1402), .Z(o[9370]) );
  AND U2102 ( .A(p_input[29370]), .B(p_input[19370]), .Z(n1402) );
  AND U2103 ( .A(p_input[9370]), .B(p_input[39370]), .Z(n1401) );
  AND U2104 ( .A(n1403), .B(n1404), .Z(o[936]) );
  AND U2105 ( .A(p_input[20936]), .B(p_input[10936]), .Z(n1404) );
  AND U2106 ( .A(p_input[936]), .B(p_input[30936]), .Z(n1403) );
  AND U2107 ( .A(n1405), .B(n1406), .Z(o[9369]) );
  AND U2108 ( .A(p_input[29369]), .B(p_input[19369]), .Z(n1406) );
  AND U2109 ( .A(p_input[9369]), .B(p_input[39369]), .Z(n1405) );
  AND U2110 ( .A(n1407), .B(n1408), .Z(o[9368]) );
  AND U2111 ( .A(p_input[29368]), .B(p_input[19368]), .Z(n1408) );
  AND U2112 ( .A(p_input[9368]), .B(p_input[39368]), .Z(n1407) );
  AND U2113 ( .A(n1409), .B(n1410), .Z(o[9367]) );
  AND U2114 ( .A(p_input[29367]), .B(p_input[19367]), .Z(n1410) );
  AND U2115 ( .A(p_input[9367]), .B(p_input[39367]), .Z(n1409) );
  AND U2116 ( .A(n1411), .B(n1412), .Z(o[9366]) );
  AND U2117 ( .A(p_input[29366]), .B(p_input[19366]), .Z(n1412) );
  AND U2118 ( .A(p_input[9366]), .B(p_input[39366]), .Z(n1411) );
  AND U2119 ( .A(n1413), .B(n1414), .Z(o[9365]) );
  AND U2120 ( .A(p_input[29365]), .B(p_input[19365]), .Z(n1414) );
  AND U2121 ( .A(p_input[9365]), .B(p_input[39365]), .Z(n1413) );
  AND U2122 ( .A(n1415), .B(n1416), .Z(o[9364]) );
  AND U2123 ( .A(p_input[29364]), .B(p_input[19364]), .Z(n1416) );
  AND U2124 ( .A(p_input[9364]), .B(p_input[39364]), .Z(n1415) );
  AND U2125 ( .A(n1417), .B(n1418), .Z(o[9363]) );
  AND U2126 ( .A(p_input[29363]), .B(p_input[19363]), .Z(n1418) );
  AND U2127 ( .A(p_input[9363]), .B(p_input[39363]), .Z(n1417) );
  AND U2128 ( .A(n1419), .B(n1420), .Z(o[9362]) );
  AND U2129 ( .A(p_input[29362]), .B(p_input[19362]), .Z(n1420) );
  AND U2130 ( .A(p_input[9362]), .B(p_input[39362]), .Z(n1419) );
  AND U2131 ( .A(n1421), .B(n1422), .Z(o[9361]) );
  AND U2132 ( .A(p_input[29361]), .B(p_input[19361]), .Z(n1422) );
  AND U2133 ( .A(p_input[9361]), .B(p_input[39361]), .Z(n1421) );
  AND U2134 ( .A(n1423), .B(n1424), .Z(o[9360]) );
  AND U2135 ( .A(p_input[29360]), .B(p_input[19360]), .Z(n1424) );
  AND U2136 ( .A(p_input[9360]), .B(p_input[39360]), .Z(n1423) );
  AND U2137 ( .A(n1425), .B(n1426), .Z(o[935]) );
  AND U2138 ( .A(p_input[20935]), .B(p_input[10935]), .Z(n1426) );
  AND U2139 ( .A(p_input[935]), .B(p_input[30935]), .Z(n1425) );
  AND U2140 ( .A(n1427), .B(n1428), .Z(o[9359]) );
  AND U2141 ( .A(p_input[29359]), .B(p_input[19359]), .Z(n1428) );
  AND U2142 ( .A(p_input[9359]), .B(p_input[39359]), .Z(n1427) );
  AND U2143 ( .A(n1429), .B(n1430), .Z(o[9358]) );
  AND U2144 ( .A(p_input[29358]), .B(p_input[19358]), .Z(n1430) );
  AND U2145 ( .A(p_input[9358]), .B(p_input[39358]), .Z(n1429) );
  AND U2146 ( .A(n1431), .B(n1432), .Z(o[9357]) );
  AND U2147 ( .A(p_input[29357]), .B(p_input[19357]), .Z(n1432) );
  AND U2148 ( .A(p_input[9357]), .B(p_input[39357]), .Z(n1431) );
  AND U2149 ( .A(n1433), .B(n1434), .Z(o[9356]) );
  AND U2150 ( .A(p_input[29356]), .B(p_input[19356]), .Z(n1434) );
  AND U2151 ( .A(p_input[9356]), .B(p_input[39356]), .Z(n1433) );
  AND U2152 ( .A(n1435), .B(n1436), .Z(o[9355]) );
  AND U2153 ( .A(p_input[29355]), .B(p_input[19355]), .Z(n1436) );
  AND U2154 ( .A(p_input[9355]), .B(p_input[39355]), .Z(n1435) );
  AND U2155 ( .A(n1437), .B(n1438), .Z(o[9354]) );
  AND U2156 ( .A(p_input[29354]), .B(p_input[19354]), .Z(n1438) );
  AND U2157 ( .A(p_input[9354]), .B(p_input[39354]), .Z(n1437) );
  AND U2158 ( .A(n1439), .B(n1440), .Z(o[9353]) );
  AND U2159 ( .A(p_input[29353]), .B(p_input[19353]), .Z(n1440) );
  AND U2160 ( .A(p_input[9353]), .B(p_input[39353]), .Z(n1439) );
  AND U2161 ( .A(n1441), .B(n1442), .Z(o[9352]) );
  AND U2162 ( .A(p_input[29352]), .B(p_input[19352]), .Z(n1442) );
  AND U2163 ( .A(p_input[9352]), .B(p_input[39352]), .Z(n1441) );
  AND U2164 ( .A(n1443), .B(n1444), .Z(o[9351]) );
  AND U2165 ( .A(p_input[29351]), .B(p_input[19351]), .Z(n1444) );
  AND U2166 ( .A(p_input[9351]), .B(p_input[39351]), .Z(n1443) );
  AND U2167 ( .A(n1445), .B(n1446), .Z(o[9350]) );
  AND U2168 ( .A(p_input[29350]), .B(p_input[19350]), .Z(n1446) );
  AND U2169 ( .A(p_input[9350]), .B(p_input[39350]), .Z(n1445) );
  AND U2170 ( .A(n1447), .B(n1448), .Z(o[934]) );
  AND U2171 ( .A(p_input[20934]), .B(p_input[10934]), .Z(n1448) );
  AND U2172 ( .A(p_input[934]), .B(p_input[30934]), .Z(n1447) );
  AND U2173 ( .A(n1449), .B(n1450), .Z(o[9349]) );
  AND U2174 ( .A(p_input[29349]), .B(p_input[19349]), .Z(n1450) );
  AND U2175 ( .A(p_input[9349]), .B(p_input[39349]), .Z(n1449) );
  AND U2176 ( .A(n1451), .B(n1452), .Z(o[9348]) );
  AND U2177 ( .A(p_input[29348]), .B(p_input[19348]), .Z(n1452) );
  AND U2178 ( .A(p_input[9348]), .B(p_input[39348]), .Z(n1451) );
  AND U2179 ( .A(n1453), .B(n1454), .Z(o[9347]) );
  AND U2180 ( .A(p_input[29347]), .B(p_input[19347]), .Z(n1454) );
  AND U2181 ( .A(p_input[9347]), .B(p_input[39347]), .Z(n1453) );
  AND U2182 ( .A(n1455), .B(n1456), .Z(o[9346]) );
  AND U2183 ( .A(p_input[29346]), .B(p_input[19346]), .Z(n1456) );
  AND U2184 ( .A(p_input[9346]), .B(p_input[39346]), .Z(n1455) );
  AND U2185 ( .A(n1457), .B(n1458), .Z(o[9345]) );
  AND U2186 ( .A(p_input[29345]), .B(p_input[19345]), .Z(n1458) );
  AND U2187 ( .A(p_input[9345]), .B(p_input[39345]), .Z(n1457) );
  AND U2188 ( .A(n1459), .B(n1460), .Z(o[9344]) );
  AND U2189 ( .A(p_input[29344]), .B(p_input[19344]), .Z(n1460) );
  AND U2190 ( .A(p_input[9344]), .B(p_input[39344]), .Z(n1459) );
  AND U2191 ( .A(n1461), .B(n1462), .Z(o[9343]) );
  AND U2192 ( .A(p_input[29343]), .B(p_input[19343]), .Z(n1462) );
  AND U2193 ( .A(p_input[9343]), .B(p_input[39343]), .Z(n1461) );
  AND U2194 ( .A(n1463), .B(n1464), .Z(o[9342]) );
  AND U2195 ( .A(p_input[29342]), .B(p_input[19342]), .Z(n1464) );
  AND U2196 ( .A(p_input[9342]), .B(p_input[39342]), .Z(n1463) );
  AND U2197 ( .A(n1465), .B(n1466), .Z(o[9341]) );
  AND U2198 ( .A(p_input[29341]), .B(p_input[19341]), .Z(n1466) );
  AND U2199 ( .A(p_input[9341]), .B(p_input[39341]), .Z(n1465) );
  AND U2200 ( .A(n1467), .B(n1468), .Z(o[9340]) );
  AND U2201 ( .A(p_input[29340]), .B(p_input[19340]), .Z(n1468) );
  AND U2202 ( .A(p_input[9340]), .B(p_input[39340]), .Z(n1467) );
  AND U2203 ( .A(n1469), .B(n1470), .Z(o[933]) );
  AND U2204 ( .A(p_input[20933]), .B(p_input[10933]), .Z(n1470) );
  AND U2205 ( .A(p_input[933]), .B(p_input[30933]), .Z(n1469) );
  AND U2206 ( .A(n1471), .B(n1472), .Z(o[9339]) );
  AND U2207 ( .A(p_input[29339]), .B(p_input[19339]), .Z(n1472) );
  AND U2208 ( .A(p_input[9339]), .B(p_input[39339]), .Z(n1471) );
  AND U2209 ( .A(n1473), .B(n1474), .Z(o[9338]) );
  AND U2210 ( .A(p_input[29338]), .B(p_input[19338]), .Z(n1474) );
  AND U2211 ( .A(p_input[9338]), .B(p_input[39338]), .Z(n1473) );
  AND U2212 ( .A(n1475), .B(n1476), .Z(o[9337]) );
  AND U2213 ( .A(p_input[29337]), .B(p_input[19337]), .Z(n1476) );
  AND U2214 ( .A(p_input[9337]), .B(p_input[39337]), .Z(n1475) );
  AND U2215 ( .A(n1477), .B(n1478), .Z(o[9336]) );
  AND U2216 ( .A(p_input[29336]), .B(p_input[19336]), .Z(n1478) );
  AND U2217 ( .A(p_input[9336]), .B(p_input[39336]), .Z(n1477) );
  AND U2218 ( .A(n1479), .B(n1480), .Z(o[9335]) );
  AND U2219 ( .A(p_input[29335]), .B(p_input[19335]), .Z(n1480) );
  AND U2220 ( .A(p_input[9335]), .B(p_input[39335]), .Z(n1479) );
  AND U2221 ( .A(n1481), .B(n1482), .Z(o[9334]) );
  AND U2222 ( .A(p_input[29334]), .B(p_input[19334]), .Z(n1482) );
  AND U2223 ( .A(p_input[9334]), .B(p_input[39334]), .Z(n1481) );
  AND U2224 ( .A(n1483), .B(n1484), .Z(o[9333]) );
  AND U2225 ( .A(p_input[29333]), .B(p_input[19333]), .Z(n1484) );
  AND U2226 ( .A(p_input[9333]), .B(p_input[39333]), .Z(n1483) );
  AND U2227 ( .A(n1485), .B(n1486), .Z(o[9332]) );
  AND U2228 ( .A(p_input[29332]), .B(p_input[19332]), .Z(n1486) );
  AND U2229 ( .A(p_input[9332]), .B(p_input[39332]), .Z(n1485) );
  AND U2230 ( .A(n1487), .B(n1488), .Z(o[9331]) );
  AND U2231 ( .A(p_input[29331]), .B(p_input[19331]), .Z(n1488) );
  AND U2232 ( .A(p_input[9331]), .B(p_input[39331]), .Z(n1487) );
  AND U2233 ( .A(n1489), .B(n1490), .Z(o[9330]) );
  AND U2234 ( .A(p_input[29330]), .B(p_input[19330]), .Z(n1490) );
  AND U2235 ( .A(p_input[9330]), .B(p_input[39330]), .Z(n1489) );
  AND U2236 ( .A(n1491), .B(n1492), .Z(o[932]) );
  AND U2237 ( .A(p_input[20932]), .B(p_input[10932]), .Z(n1492) );
  AND U2238 ( .A(p_input[932]), .B(p_input[30932]), .Z(n1491) );
  AND U2239 ( .A(n1493), .B(n1494), .Z(o[9329]) );
  AND U2240 ( .A(p_input[29329]), .B(p_input[19329]), .Z(n1494) );
  AND U2241 ( .A(p_input[9329]), .B(p_input[39329]), .Z(n1493) );
  AND U2242 ( .A(n1495), .B(n1496), .Z(o[9328]) );
  AND U2243 ( .A(p_input[29328]), .B(p_input[19328]), .Z(n1496) );
  AND U2244 ( .A(p_input[9328]), .B(p_input[39328]), .Z(n1495) );
  AND U2245 ( .A(n1497), .B(n1498), .Z(o[9327]) );
  AND U2246 ( .A(p_input[29327]), .B(p_input[19327]), .Z(n1498) );
  AND U2247 ( .A(p_input[9327]), .B(p_input[39327]), .Z(n1497) );
  AND U2248 ( .A(n1499), .B(n1500), .Z(o[9326]) );
  AND U2249 ( .A(p_input[29326]), .B(p_input[19326]), .Z(n1500) );
  AND U2250 ( .A(p_input[9326]), .B(p_input[39326]), .Z(n1499) );
  AND U2251 ( .A(n1501), .B(n1502), .Z(o[9325]) );
  AND U2252 ( .A(p_input[29325]), .B(p_input[19325]), .Z(n1502) );
  AND U2253 ( .A(p_input[9325]), .B(p_input[39325]), .Z(n1501) );
  AND U2254 ( .A(n1503), .B(n1504), .Z(o[9324]) );
  AND U2255 ( .A(p_input[29324]), .B(p_input[19324]), .Z(n1504) );
  AND U2256 ( .A(p_input[9324]), .B(p_input[39324]), .Z(n1503) );
  AND U2257 ( .A(n1505), .B(n1506), .Z(o[9323]) );
  AND U2258 ( .A(p_input[29323]), .B(p_input[19323]), .Z(n1506) );
  AND U2259 ( .A(p_input[9323]), .B(p_input[39323]), .Z(n1505) );
  AND U2260 ( .A(n1507), .B(n1508), .Z(o[9322]) );
  AND U2261 ( .A(p_input[29322]), .B(p_input[19322]), .Z(n1508) );
  AND U2262 ( .A(p_input[9322]), .B(p_input[39322]), .Z(n1507) );
  AND U2263 ( .A(n1509), .B(n1510), .Z(o[9321]) );
  AND U2264 ( .A(p_input[29321]), .B(p_input[19321]), .Z(n1510) );
  AND U2265 ( .A(p_input[9321]), .B(p_input[39321]), .Z(n1509) );
  AND U2266 ( .A(n1511), .B(n1512), .Z(o[9320]) );
  AND U2267 ( .A(p_input[29320]), .B(p_input[19320]), .Z(n1512) );
  AND U2268 ( .A(p_input[9320]), .B(p_input[39320]), .Z(n1511) );
  AND U2269 ( .A(n1513), .B(n1514), .Z(o[931]) );
  AND U2270 ( .A(p_input[20931]), .B(p_input[10931]), .Z(n1514) );
  AND U2271 ( .A(p_input[931]), .B(p_input[30931]), .Z(n1513) );
  AND U2272 ( .A(n1515), .B(n1516), .Z(o[9319]) );
  AND U2273 ( .A(p_input[29319]), .B(p_input[19319]), .Z(n1516) );
  AND U2274 ( .A(p_input[9319]), .B(p_input[39319]), .Z(n1515) );
  AND U2275 ( .A(n1517), .B(n1518), .Z(o[9318]) );
  AND U2276 ( .A(p_input[29318]), .B(p_input[19318]), .Z(n1518) );
  AND U2277 ( .A(p_input[9318]), .B(p_input[39318]), .Z(n1517) );
  AND U2278 ( .A(n1519), .B(n1520), .Z(o[9317]) );
  AND U2279 ( .A(p_input[29317]), .B(p_input[19317]), .Z(n1520) );
  AND U2280 ( .A(p_input[9317]), .B(p_input[39317]), .Z(n1519) );
  AND U2281 ( .A(n1521), .B(n1522), .Z(o[9316]) );
  AND U2282 ( .A(p_input[29316]), .B(p_input[19316]), .Z(n1522) );
  AND U2283 ( .A(p_input[9316]), .B(p_input[39316]), .Z(n1521) );
  AND U2284 ( .A(n1523), .B(n1524), .Z(o[9315]) );
  AND U2285 ( .A(p_input[29315]), .B(p_input[19315]), .Z(n1524) );
  AND U2286 ( .A(p_input[9315]), .B(p_input[39315]), .Z(n1523) );
  AND U2287 ( .A(n1525), .B(n1526), .Z(o[9314]) );
  AND U2288 ( .A(p_input[29314]), .B(p_input[19314]), .Z(n1526) );
  AND U2289 ( .A(p_input[9314]), .B(p_input[39314]), .Z(n1525) );
  AND U2290 ( .A(n1527), .B(n1528), .Z(o[9313]) );
  AND U2291 ( .A(p_input[29313]), .B(p_input[19313]), .Z(n1528) );
  AND U2292 ( .A(p_input[9313]), .B(p_input[39313]), .Z(n1527) );
  AND U2293 ( .A(n1529), .B(n1530), .Z(o[9312]) );
  AND U2294 ( .A(p_input[29312]), .B(p_input[19312]), .Z(n1530) );
  AND U2295 ( .A(p_input[9312]), .B(p_input[39312]), .Z(n1529) );
  AND U2296 ( .A(n1531), .B(n1532), .Z(o[9311]) );
  AND U2297 ( .A(p_input[29311]), .B(p_input[19311]), .Z(n1532) );
  AND U2298 ( .A(p_input[9311]), .B(p_input[39311]), .Z(n1531) );
  AND U2299 ( .A(n1533), .B(n1534), .Z(o[9310]) );
  AND U2300 ( .A(p_input[29310]), .B(p_input[19310]), .Z(n1534) );
  AND U2301 ( .A(p_input[9310]), .B(p_input[39310]), .Z(n1533) );
  AND U2302 ( .A(n1535), .B(n1536), .Z(o[930]) );
  AND U2303 ( .A(p_input[20930]), .B(p_input[10930]), .Z(n1536) );
  AND U2304 ( .A(p_input[930]), .B(p_input[30930]), .Z(n1535) );
  AND U2305 ( .A(n1537), .B(n1538), .Z(o[9309]) );
  AND U2306 ( .A(p_input[29309]), .B(p_input[19309]), .Z(n1538) );
  AND U2307 ( .A(p_input[9309]), .B(p_input[39309]), .Z(n1537) );
  AND U2308 ( .A(n1539), .B(n1540), .Z(o[9308]) );
  AND U2309 ( .A(p_input[29308]), .B(p_input[19308]), .Z(n1540) );
  AND U2310 ( .A(p_input[9308]), .B(p_input[39308]), .Z(n1539) );
  AND U2311 ( .A(n1541), .B(n1542), .Z(o[9307]) );
  AND U2312 ( .A(p_input[29307]), .B(p_input[19307]), .Z(n1542) );
  AND U2313 ( .A(p_input[9307]), .B(p_input[39307]), .Z(n1541) );
  AND U2314 ( .A(n1543), .B(n1544), .Z(o[9306]) );
  AND U2315 ( .A(p_input[29306]), .B(p_input[19306]), .Z(n1544) );
  AND U2316 ( .A(p_input[9306]), .B(p_input[39306]), .Z(n1543) );
  AND U2317 ( .A(n1545), .B(n1546), .Z(o[9305]) );
  AND U2318 ( .A(p_input[29305]), .B(p_input[19305]), .Z(n1546) );
  AND U2319 ( .A(p_input[9305]), .B(p_input[39305]), .Z(n1545) );
  AND U2320 ( .A(n1547), .B(n1548), .Z(o[9304]) );
  AND U2321 ( .A(p_input[29304]), .B(p_input[19304]), .Z(n1548) );
  AND U2322 ( .A(p_input[9304]), .B(p_input[39304]), .Z(n1547) );
  AND U2323 ( .A(n1549), .B(n1550), .Z(o[9303]) );
  AND U2324 ( .A(p_input[29303]), .B(p_input[19303]), .Z(n1550) );
  AND U2325 ( .A(p_input[9303]), .B(p_input[39303]), .Z(n1549) );
  AND U2326 ( .A(n1551), .B(n1552), .Z(o[9302]) );
  AND U2327 ( .A(p_input[29302]), .B(p_input[19302]), .Z(n1552) );
  AND U2328 ( .A(p_input[9302]), .B(p_input[39302]), .Z(n1551) );
  AND U2329 ( .A(n1553), .B(n1554), .Z(o[9301]) );
  AND U2330 ( .A(p_input[29301]), .B(p_input[19301]), .Z(n1554) );
  AND U2331 ( .A(p_input[9301]), .B(p_input[39301]), .Z(n1553) );
  AND U2332 ( .A(n1555), .B(n1556), .Z(o[9300]) );
  AND U2333 ( .A(p_input[29300]), .B(p_input[19300]), .Z(n1556) );
  AND U2334 ( .A(p_input[9300]), .B(p_input[39300]), .Z(n1555) );
  AND U2335 ( .A(n1557), .B(n1558), .Z(o[92]) );
  AND U2336 ( .A(p_input[20092]), .B(p_input[10092]), .Z(n1558) );
  AND U2337 ( .A(p_input[92]), .B(p_input[30092]), .Z(n1557) );
  AND U2338 ( .A(n1559), .B(n1560), .Z(o[929]) );
  AND U2339 ( .A(p_input[20929]), .B(p_input[10929]), .Z(n1560) );
  AND U2340 ( .A(p_input[929]), .B(p_input[30929]), .Z(n1559) );
  AND U2341 ( .A(n1561), .B(n1562), .Z(o[9299]) );
  AND U2342 ( .A(p_input[29299]), .B(p_input[19299]), .Z(n1562) );
  AND U2343 ( .A(p_input[9299]), .B(p_input[39299]), .Z(n1561) );
  AND U2344 ( .A(n1563), .B(n1564), .Z(o[9298]) );
  AND U2345 ( .A(p_input[29298]), .B(p_input[19298]), .Z(n1564) );
  AND U2346 ( .A(p_input[9298]), .B(p_input[39298]), .Z(n1563) );
  AND U2347 ( .A(n1565), .B(n1566), .Z(o[9297]) );
  AND U2348 ( .A(p_input[29297]), .B(p_input[19297]), .Z(n1566) );
  AND U2349 ( .A(p_input[9297]), .B(p_input[39297]), .Z(n1565) );
  AND U2350 ( .A(n1567), .B(n1568), .Z(o[9296]) );
  AND U2351 ( .A(p_input[29296]), .B(p_input[19296]), .Z(n1568) );
  AND U2352 ( .A(p_input[9296]), .B(p_input[39296]), .Z(n1567) );
  AND U2353 ( .A(n1569), .B(n1570), .Z(o[9295]) );
  AND U2354 ( .A(p_input[29295]), .B(p_input[19295]), .Z(n1570) );
  AND U2355 ( .A(p_input[9295]), .B(p_input[39295]), .Z(n1569) );
  AND U2356 ( .A(n1571), .B(n1572), .Z(o[9294]) );
  AND U2357 ( .A(p_input[29294]), .B(p_input[19294]), .Z(n1572) );
  AND U2358 ( .A(p_input[9294]), .B(p_input[39294]), .Z(n1571) );
  AND U2359 ( .A(n1573), .B(n1574), .Z(o[9293]) );
  AND U2360 ( .A(p_input[29293]), .B(p_input[19293]), .Z(n1574) );
  AND U2361 ( .A(p_input[9293]), .B(p_input[39293]), .Z(n1573) );
  AND U2362 ( .A(n1575), .B(n1576), .Z(o[9292]) );
  AND U2363 ( .A(p_input[29292]), .B(p_input[19292]), .Z(n1576) );
  AND U2364 ( .A(p_input[9292]), .B(p_input[39292]), .Z(n1575) );
  AND U2365 ( .A(n1577), .B(n1578), .Z(o[9291]) );
  AND U2366 ( .A(p_input[29291]), .B(p_input[19291]), .Z(n1578) );
  AND U2367 ( .A(p_input[9291]), .B(p_input[39291]), .Z(n1577) );
  AND U2368 ( .A(n1579), .B(n1580), .Z(o[9290]) );
  AND U2369 ( .A(p_input[29290]), .B(p_input[19290]), .Z(n1580) );
  AND U2370 ( .A(p_input[9290]), .B(p_input[39290]), .Z(n1579) );
  AND U2371 ( .A(n1581), .B(n1582), .Z(o[928]) );
  AND U2372 ( .A(p_input[20928]), .B(p_input[10928]), .Z(n1582) );
  AND U2373 ( .A(p_input[928]), .B(p_input[30928]), .Z(n1581) );
  AND U2374 ( .A(n1583), .B(n1584), .Z(o[9289]) );
  AND U2375 ( .A(p_input[29289]), .B(p_input[19289]), .Z(n1584) );
  AND U2376 ( .A(p_input[9289]), .B(p_input[39289]), .Z(n1583) );
  AND U2377 ( .A(n1585), .B(n1586), .Z(o[9288]) );
  AND U2378 ( .A(p_input[29288]), .B(p_input[19288]), .Z(n1586) );
  AND U2379 ( .A(p_input[9288]), .B(p_input[39288]), .Z(n1585) );
  AND U2380 ( .A(n1587), .B(n1588), .Z(o[9287]) );
  AND U2381 ( .A(p_input[29287]), .B(p_input[19287]), .Z(n1588) );
  AND U2382 ( .A(p_input[9287]), .B(p_input[39287]), .Z(n1587) );
  AND U2383 ( .A(n1589), .B(n1590), .Z(o[9286]) );
  AND U2384 ( .A(p_input[29286]), .B(p_input[19286]), .Z(n1590) );
  AND U2385 ( .A(p_input[9286]), .B(p_input[39286]), .Z(n1589) );
  AND U2386 ( .A(n1591), .B(n1592), .Z(o[9285]) );
  AND U2387 ( .A(p_input[29285]), .B(p_input[19285]), .Z(n1592) );
  AND U2388 ( .A(p_input[9285]), .B(p_input[39285]), .Z(n1591) );
  AND U2389 ( .A(n1593), .B(n1594), .Z(o[9284]) );
  AND U2390 ( .A(p_input[29284]), .B(p_input[19284]), .Z(n1594) );
  AND U2391 ( .A(p_input[9284]), .B(p_input[39284]), .Z(n1593) );
  AND U2392 ( .A(n1595), .B(n1596), .Z(o[9283]) );
  AND U2393 ( .A(p_input[29283]), .B(p_input[19283]), .Z(n1596) );
  AND U2394 ( .A(p_input[9283]), .B(p_input[39283]), .Z(n1595) );
  AND U2395 ( .A(n1597), .B(n1598), .Z(o[9282]) );
  AND U2396 ( .A(p_input[29282]), .B(p_input[19282]), .Z(n1598) );
  AND U2397 ( .A(p_input[9282]), .B(p_input[39282]), .Z(n1597) );
  AND U2398 ( .A(n1599), .B(n1600), .Z(o[9281]) );
  AND U2399 ( .A(p_input[29281]), .B(p_input[19281]), .Z(n1600) );
  AND U2400 ( .A(p_input[9281]), .B(p_input[39281]), .Z(n1599) );
  AND U2401 ( .A(n1601), .B(n1602), .Z(o[9280]) );
  AND U2402 ( .A(p_input[29280]), .B(p_input[19280]), .Z(n1602) );
  AND U2403 ( .A(p_input[9280]), .B(p_input[39280]), .Z(n1601) );
  AND U2404 ( .A(n1603), .B(n1604), .Z(o[927]) );
  AND U2405 ( .A(p_input[20927]), .B(p_input[10927]), .Z(n1604) );
  AND U2406 ( .A(p_input[927]), .B(p_input[30927]), .Z(n1603) );
  AND U2407 ( .A(n1605), .B(n1606), .Z(o[9279]) );
  AND U2408 ( .A(p_input[29279]), .B(p_input[19279]), .Z(n1606) );
  AND U2409 ( .A(p_input[9279]), .B(p_input[39279]), .Z(n1605) );
  AND U2410 ( .A(n1607), .B(n1608), .Z(o[9278]) );
  AND U2411 ( .A(p_input[29278]), .B(p_input[19278]), .Z(n1608) );
  AND U2412 ( .A(p_input[9278]), .B(p_input[39278]), .Z(n1607) );
  AND U2413 ( .A(n1609), .B(n1610), .Z(o[9277]) );
  AND U2414 ( .A(p_input[29277]), .B(p_input[19277]), .Z(n1610) );
  AND U2415 ( .A(p_input[9277]), .B(p_input[39277]), .Z(n1609) );
  AND U2416 ( .A(n1611), .B(n1612), .Z(o[9276]) );
  AND U2417 ( .A(p_input[29276]), .B(p_input[19276]), .Z(n1612) );
  AND U2418 ( .A(p_input[9276]), .B(p_input[39276]), .Z(n1611) );
  AND U2419 ( .A(n1613), .B(n1614), .Z(o[9275]) );
  AND U2420 ( .A(p_input[29275]), .B(p_input[19275]), .Z(n1614) );
  AND U2421 ( .A(p_input[9275]), .B(p_input[39275]), .Z(n1613) );
  AND U2422 ( .A(n1615), .B(n1616), .Z(o[9274]) );
  AND U2423 ( .A(p_input[29274]), .B(p_input[19274]), .Z(n1616) );
  AND U2424 ( .A(p_input[9274]), .B(p_input[39274]), .Z(n1615) );
  AND U2425 ( .A(n1617), .B(n1618), .Z(o[9273]) );
  AND U2426 ( .A(p_input[29273]), .B(p_input[19273]), .Z(n1618) );
  AND U2427 ( .A(p_input[9273]), .B(p_input[39273]), .Z(n1617) );
  AND U2428 ( .A(n1619), .B(n1620), .Z(o[9272]) );
  AND U2429 ( .A(p_input[29272]), .B(p_input[19272]), .Z(n1620) );
  AND U2430 ( .A(p_input[9272]), .B(p_input[39272]), .Z(n1619) );
  AND U2431 ( .A(n1621), .B(n1622), .Z(o[9271]) );
  AND U2432 ( .A(p_input[29271]), .B(p_input[19271]), .Z(n1622) );
  AND U2433 ( .A(p_input[9271]), .B(p_input[39271]), .Z(n1621) );
  AND U2434 ( .A(n1623), .B(n1624), .Z(o[9270]) );
  AND U2435 ( .A(p_input[29270]), .B(p_input[19270]), .Z(n1624) );
  AND U2436 ( .A(p_input[9270]), .B(p_input[39270]), .Z(n1623) );
  AND U2437 ( .A(n1625), .B(n1626), .Z(o[926]) );
  AND U2438 ( .A(p_input[20926]), .B(p_input[10926]), .Z(n1626) );
  AND U2439 ( .A(p_input[926]), .B(p_input[30926]), .Z(n1625) );
  AND U2440 ( .A(n1627), .B(n1628), .Z(o[9269]) );
  AND U2441 ( .A(p_input[29269]), .B(p_input[19269]), .Z(n1628) );
  AND U2442 ( .A(p_input[9269]), .B(p_input[39269]), .Z(n1627) );
  AND U2443 ( .A(n1629), .B(n1630), .Z(o[9268]) );
  AND U2444 ( .A(p_input[29268]), .B(p_input[19268]), .Z(n1630) );
  AND U2445 ( .A(p_input[9268]), .B(p_input[39268]), .Z(n1629) );
  AND U2446 ( .A(n1631), .B(n1632), .Z(o[9267]) );
  AND U2447 ( .A(p_input[29267]), .B(p_input[19267]), .Z(n1632) );
  AND U2448 ( .A(p_input[9267]), .B(p_input[39267]), .Z(n1631) );
  AND U2449 ( .A(n1633), .B(n1634), .Z(o[9266]) );
  AND U2450 ( .A(p_input[29266]), .B(p_input[19266]), .Z(n1634) );
  AND U2451 ( .A(p_input[9266]), .B(p_input[39266]), .Z(n1633) );
  AND U2452 ( .A(n1635), .B(n1636), .Z(o[9265]) );
  AND U2453 ( .A(p_input[29265]), .B(p_input[19265]), .Z(n1636) );
  AND U2454 ( .A(p_input[9265]), .B(p_input[39265]), .Z(n1635) );
  AND U2455 ( .A(n1637), .B(n1638), .Z(o[9264]) );
  AND U2456 ( .A(p_input[29264]), .B(p_input[19264]), .Z(n1638) );
  AND U2457 ( .A(p_input[9264]), .B(p_input[39264]), .Z(n1637) );
  AND U2458 ( .A(n1639), .B(n1640), .Z(o[9263]) );
  AND U2459 ( .A(p_input[29263]), .B(p_input[19263]), .Z(n1640) );
  AND U2460 ( .A(p_input[9263]), .B(p_input[39263]), .Z(n1639) );
  AND U2461 ( .A(n1641), .B(n1642), .Z(o[9262]) );
  AND U2462 ( .A(p_input[29262]), .B(p_input[19262]), .Z(n1642) );
  AND U2463 ( .A(p_input[9262]), .B(p_input[39262]), .Z(n1641) );
  AND U2464 ( .A(n1643), .B(n1644), .Z(o[9261]) );
  AND U2465 ( .A(p_input[29261]), .B(p_input[19261]), .Z(n1644) );
  AND U2466 ( .A(p_input[9261]), .B(p_input[39261]), .Z(n1643) );
  AND U2467 ( .A(n1645), .B(n1646), .Z(o[9260]) );
  AND U2468 ( .A(p_input[29260]), .B(p_input[19260]), .Z(n1646) );
  AND U2469 ( .A(p_input[9260]), .B(p_input[39260]), .Z(n1645) );
  AND U2470 ( .A(n1647), .B(n1648), .Z(o[925]) );
  AND U2471 ( .A(p_input[20925]), .B(p_input[10925]), .Z(n1648) );
  AND U2472 ( .A(p_input[925]), .B(p_input[30925]), .Z(n1647) );
  AND U2473 ( .A(n1649), .B(n1650), .Z(o[9259]) );
  AND U2474 ( .A(p_input[29259]), .B(p_input[19259]), .Z(n1650) );
  AND U2475 ( .A(p_input[9259]), .B(p_input[39259]), .Z(n1649) );
  AND U2476 ( .A(n1651), .B(n1652), .Z(o[9258]) );
  AND U2477 ( .A(p_input[29258]), .B(p_input[19258]), .Z(n1652) );
  AND U2478 ( .A(p_input[9258]), .B(p_input[39258]), .Z(n1651) );
  AND U2479 ( .A(n1653), .B(n1654), .Z(o[9257]) );
  AND U2480 ( .A(p_input[29257]), .B(p_input[19257]), .Z(n1654) );
  AND U2481 ( .A(p_input[9257]), .B(p_input[39257]), .Z(n1653) );
  AND U2482 ( .A(n1655), .B(n1656), .Z(o[9256]) );
  AND U2483 ( .A(p_input[29256]), .B(p_input[19256]), .Z(n1656) );
  AND U2484 ( .A(p_input[9256]), .B(p_input[39256]), .Z(n1655) );
  AND U2485 ( .A(n1657), .B(n1658), .Z(o[9255]) );
  AND U2486 ( .A(p_input[29255]), .B(p_input[19255]), .Z(n1658) );
  AND U2487 ( .A(p_input[9255]), .B(p_input[39255]), .Z(n1657) );
  AND U2488 ( .A(n1659), .B(n1660), .Z(o[9254]) );
  AND U2489 ( .A(p_input[29254]), .B(p_input[19254]), .Z(n1660) );
  AND U2490 ( .A(p_input[9254]), .B(p_input[39254]), .Z(n1659) );
  AND U2491 ( .A(n1661), .B(n1662), .Z(o[9253]) );
  AND U2492 ( .A(p_input[29253]), .B(p_input[19253]), .Z(n1662) );
  AND U2493 ( .A(p_input[9253]), .B(p_input[39253]), .Z(n1661) );
  AND U2494 ( .A(n1663), .B(n1664), .Z(o[9252]) );
  AND U2495 ( .A(p_input[29252]), .B(p_input[19252]), .Z(n1664) );
  AND U2496 ( .A(p_input[9252]), .B(p_input[39252]), .Z(n1663) );
  AND U2497 ( .A(n1665), .B(n1666), .Z(o[9251]) );
  AND U2498 ( .A(p_input[29251]), .B(p_input[19251]), .Z(n1666) );
  AND U2499 ( .A(p_input[9251]), .B(p_input[39251]), .Z(n1665) );
  AND U2500 ( .A(n1667), .B(n1668), .Z(o[9250]) );
  AND U2501 ( .A(p_input[29250]), .B(p_input[19250]), .Z(n1668) );
  AND U2502 ( .A(p_input[9250]), .B(p_input[39250]), .Z(n1667) );
  AND U2503 ( .A(n1669), .B(n1670), .Z(o[924]) );
  AND U2504 ( .A(p_input[20924]), .B(p_input[10924]), .Z(n1670) );
  AND U2505 ( .A(p_input[924]), .B(p_input[30924]), .Z(n1669) );
  AND U2506 ( .A(n1671), .B(n1672), .Z(o[9249]) );
  AND U2507 ( .A(p_input[29249]), .B(p_input[19249]), .Z(n1672) );
  AND U2508 ( .A(p_input[9249]), .B(p_input[39249]), .Z(n1671) );
  AND U2509 ( .A(n1673), .B(n1674), .Z(o[9248]) );
  AND U2510 ( .A(p_input[29248]), .B(p_input[19248]), .Z(n1674) );
  AND U2511 ( .A(p_input[9248]), .B(p_input[39248]), .Z(n1673) );
  AND U2512 ( .A(n1675), .B(n1676), .Z(o[9247]) );
  AND U2513 ( .A(p_input[29247]), .B(p_input[19247]), .Z(n1676) );
  AND U2514 ( .A(p_input[9247]), .B(p_input[39247]), .Z(n1675) );
  AND U2515 ( .A(n1677), .B(n1678), .Z(o[9246]) );
  AND U2516 ( .A(p_input[29246]), .B(p_input[19246]), .Z(n1678) );
  AND U2517 ( .A(p_input[9246]), .B(p_input[39246]), .Z(n1677) );
  AND U2518 ( .A(n1679), .B(n1680), .Z(o[9245]) );
  AND U2519 ( .A(p_input[29245]), .B(p_input[19245]), .Z(n1680) );
  AND U2520 ( .A(p_input[9245]), .B(p_input[39245]), .Z(n1679) );
  AND U2521 ( .A(n1681), .B(n1682), .Z(o[9244]) );
  AND U2522 ( .A(p_input[29244]), .B(p_input[19244]), .Z(n1682) );
  AND U2523 ( .A(p_input[9244]), .B(p_input[39244]), .Z(n1681) );
  AND U2524 ( .A(n1683), .B(n1684), .Z(o[9243]) );
  AND U2525 ( .A(p_input[29243]), .B(p_input[19243]), .Z(n1684) );
  AND U2526 ( .A(p_input[9243]), .B(p_input[39243]), .Z(n1683) );
  AND U2527 ( .A(n1685), .B(n1686), .Z(o[9242]) );
  AND U2528 ( .A(p_input[29242]), .B(p_input[19242]), .Z(n1686) );
  AND U2529 ( .A(p_input[9242]), .B(p_input[39242]), .Z(n1685) );
  AND U2530 ( .A(n1687), .B(n1688), .Z(o[9241]) );
  AND U2531 ( .A(p_input[29241]), .B(p_input[19241]), .Z(n1688) );
  AND U2532 ( .A(p_input[9241]), .B(p_input[39241]), .Z(n1687) );
  AND U2533 ( .A(n1689), .B(n1690), .Z(o[9240]) );
  AND U2534 ( .A(p_input[29240]), .B(p_input[19240]), .Z(n1690) );
  AND U2535 ( .A(p_input[9240]), .B(p_input[39240]), .Z(n1689) );
  AND U2536 ( .A(n1691), .B(n1692), .Z(o[923]) );
  AND U2537 ( .A(p_input[20923]), .B(p_input[10923]), .Z(n1692) );
  AND U2538 ( .A(p_input[923]), .B(p_input[30923]), .Z(n1691) );
  AND U2539 ( .A(n1693), .B(n1694), .Z(o[9239]) );
  AND U2540 ( .A(p_input[29239]), .B(p_input[19239]), .Z(n1694) );
  AND U2541 ( .A(p_input[9239]), .B(p_input[39239]), .Z(n1693) );
  AND U2542 ( .A(n1695), .B(n1696), .Z(o[9238]) );
  AND U2543 ( .A(p_input[29238]), .B(p_input[19238]), .Z(n1696) );
  AND U2544 ( .A(p_input[9238]), .B(p_input[39238]), .Z(n1695) );
  AND U2545 ( .A(n1697), .B(n1698), .Z(o[9237]) );
  AND U2546 ( .A(p_input[29237]), .B(p_input[19237]), .Z(n1698) );
  AND U2547 ( .A(p_input[9237]), .B(p_input[39237]), .Z(n1697) );
  AND U2548 ( .A(n1699), .B(n1700), .Z(o[9236]) );
  AND U2549 ( .A(p_input[29236]), .B(p_input[19236]), .Z(n1700) );
  AND U2550 ( .A(p_input[9236]), .B(p_input[39236]), .Z(n1699) );
  AND U2551 ( .A(n1701), .B(n1702), .Z(o[9235]) );
  AND U2552 ( .A(p_input[29235]), .B(p_input[19235]), .Z(n1702) );
  AND U2553 ( .A(p_input[9235]), .B(p_input[39235]), .Z(n1701) );
  AND U2554 ( .A(n1703), .B(n1704), .Z(o[9234]) );
  AND U2555 ( .A(p_input[29234]), .B(p_input[19234]), .Z(n1704) );
  AND U2556 ( .A(p_input[9234]), .B(p_input[39234]), .Z(n1703) );
  AND U2557 ( .A(n1705), .B(n1706), .Z(o[9233]) );
  AND U2558 ( .A(p_input[29233]), .B(p_input[19233]), .Z(n1706) );
  AND U2559 ( .A(p_input[9233]), .B(p_input[39233]), .Z(n1705) );
  AND U2560 ( .A(n1707), .B(n1708), .Z(o[9232]) );
  AND U2561 ( .A(p_input[29232]), .B(p_input[19232]), .Z(n1708) );
  AND U2562 ( .A(p_input[9232]), .B(p_input[39232]), .Z(n1707) );
  AND U2563 ( .A(n1709), .B(n1710), .Z(o[9231]) );
  AND U2564 ( .A(p_input[29231]), .B(p_input[19231]), .Z(n1710) );
  AND U2565 ( .A(p_input[9231]), .B(p_input[39231]), .Z(n1709) );
  AND U2566 ( .A(n1711), .B(n1712), .Z(o[9230]) );
  AND U2567 ( .A(p_input[29230]), .B(p_input[19230]), .Z(n1712) );
  AND U2568 ( .A(p_input[9230]), .B(p_input[39230]), .Z(n1711) );
  AND U2569 ( .A(n1713), .B(n1714), .Z(o[922]) );
  AND U2570 ( .A(p_input[20922]), .B(p_input[10922]), .Z(n1714) );
  AND U2571 ( .A(p_input[922]), .B(p_input[30922]), .Z(n1713) );
  AND U2572 ( .A(n1715), .B(n1716), .Z(o[9229]) );
  AND U2573 ( .A(p_input[29229]), .B(p_input[19229]), .Z(n1716) );
  AND U2574 ( .A(p_input[9229]), .B(p_input[39229]), .Z(n1715) );
  AND U2575 ( .A(n1717), .B(n1718), .Z(o[9228]) );
  AND U2576 ( .A(p_input[29228]), .B(p_input[19228]), .Z(n1718) );
  AND U2577 ( .A(p_input[9228]), .B(p_input[39228]), .Z(n1717) );
  AND U2578 ( .A(n1719), .B(n1720), .Z(o[9227]) );
  AND U2579 ( .A(p_input[29227]), .B(p_input[19227]), .Z(n1720) );
  AND U2580 ( .A(p_input[9227]), .B(p_input[39227]), .Z(n1719) );
  AND U2581 ( .A(n1721), .B(n1722), .Z(o[9226]) );
  AND U2582 ( .A(p_input[29226]), .B(p_input[19226]), .Z(n1722) );
  AND U2583 ( .A(p_input[9226]), .B(p_input[39226]), .Z(n1721) );
  AND U2584 ( .A(n1723), .B(n1724), .Z(o[9225]) );
  AND U2585 ( .A(p_input[29225]), .B(p_input[19225]), .Z(n1724) );
  AND U2586 ( .A(p_input[9225]), .B(p_input[39225]), .Z(n1723) );
  AND U2587 ( .A(n1725), .B(n1726), .Z(o[9224]) );
  AND U2588 ( .A(p_input[29224]), .B(p_input[19224]), .Z(n1726) );
  AND U2589 ( .A(p_input[9224]), .B(p_input[39224]), .Z(n1725) );
  AND U2590 ( .A(n1727), .B(n1728), .Z(o[9223]) );
  AND U2591 ( .A(p_input[29223]), .B(p_input[19223]), .Z(n1728) );
  AND U2592 ( .A(p_input[9223]), .B(p_input[39223]), .Z(n1727) );
  AND U2593 ( .A(n1729), .B(n1730), .Z(o[9222]) );
  AND U2594 ( .A(p_input[29222]), .B(p_input[19222]), .Z(n1730) );
  AND U2595 ( .A(p_input[9222]), .B(p_input[39222]), .Z(n1729) );
  AND U2596 ( .A(n1731), .B(n1732), .Z(o[9221]) );
  AND U2597 ( .A(p_input[29221]), .B(p_input[19221]), .Z(n1732) );
  AND U2598 ( .A(p_input[9221]), .B(p_input[39221]), .Z(n1731) );
  AND U2599 ( .A(n1733), .B(n1734), .Z(o[9220]) );
  AND U2600 ( .A(p_input[29220]), .B(p_input[19220]), .Z(n1734) );
  AND U2601 ( .A(p_input[9220]), .B(p_input[39220]), .Z(n1733) );
  AND U2602 ( .A(n1735), .B(n1736), .Z(o[921]) );
  AND U2603 ( .A(p_input[20921]), .B(p_input[10921]), .Z(n1736) );
  AND U2604 ( .A(p_input[921]), .B(p_input[30921]), .Z(n1735) );
  AND U2605 ( .A(n1737), .B(n1738), .Z(o[9219]) );
  AND U2606 ( .A(p_input[29219]), .B(p_input[19219]), .Z(n1738) );
  AND U2607 ( .A(p_input[9219]), .B(p_input[39219]), .Z(n1737) );
  AND U2608 ( .A(n1739), .B(n1740), .Z(o[9218]) );
  AND U2609 ( .A(p_input[29218]), .B(p_input[19218]), .Z(n1740) );
  AND U2610 ( .A(p_input[9218]), .B(p_input[39218]), .Z(n1739) );
  AND U2611 ( .A(n1741), .B(n1742), .Z(o[9217]) );
  AND U2612 ( .A(p_input[29217]), .B(p_input[19217]), .Z(n1742) );
  AND U2613 ( .A(p_input[9217]), .B(p_input[39217]), .Z(n1741) );
  AND U2614 ( .A(n1743), .B(n1744), .Z(o[9216]) );
  AND U2615 ( .A(p_input[29216]), .B(p_input[19216]), .Z(n1744) );
  AND U2616 ( .A(p_input[9216]), .B(p_input[39216]), .Z(n1743) );
  AND U2617 ( .A(n1745), .B(n1746), .Z(o[9215]) );
  AND U2618 ( .A(p_input[29215]), .B(p_input[19215]), .Z(n1746) );
  AND U2619 ( .A(p_input[9215]), .B(p_input[39215]), .Z(n1745) );
  AND U2620 ( .A(n1747), .B(n1748), .Z(o[9214]) );
  AND U2621 ( .A(p_input[29214]), .B(p_input[19214]), .Z(n1748) );
  AND U2622 ( .A(p_input[9214]), .B(p_input[39214]), .Z(n1747) );
  AND U2623 ( .A(n1749), .B(n1750), .Z(o[9213]) );
  AND U2624 ( .A(p_input[29213]), .B(p_input[19213]), .Z(n1750) );
  AND U2625 ( .A(p_input[9213]), .B(p_input[39213]), .Z(n1749) );
  AND U2626 ( .A(n1751), .B(n1752), .Z(o[9212]) );
  AND U2627 ( .A(p_input[29212]), .B(p_input[19212]), .Z(n1752) );
  AND U2628 ( .A(p_input[9212]), .B(p_input[39212]), .Z(n1751) );
  AND U2629 ( .A(n1753), .B(n1754), .Z(o[9211]) );
  AND U2630 ( .A(p_input[29211]), .B(p_input[19211]), .Z(n1754) );
  AND U2631 ( .A(p_input[9211]), .B(p_input[39211]), .Z(n1753) );
  AND U2632 ( .A(n1755), .B(n1756), .Z(o[9210]) );
  AND U2633 ( .A(p_input[29210]), .B(p_input[19210]), .Z(n1756) );
  AND U2634 ( .A(p_input[9210]), .B(p_input[39210]), .Z(n1755) );
  AND U2635 ( .A(n1757), .B(n1758), .Z(o[920]) );
  AND U2636 ( .A(p_input[20920]), .B(p_input[10920]), .Z(n1758) );
  AND U2637 ( .A(p_input[920]), .B(p_input[30920]), .Z(n1757) );
  AND U2638 ( .A(n1759), .B(n1760), .Z(o[9209]) );
  AND U2639 ( .A(p_input[29209]), .B(p_input[19209]), .Z(n1760) );
  AND U2640 ( .A(p_input[9209]), .B(p_input[39209]), .Z(n1759) );
  AND U2641 ( .A(n1761), .B(n1762), .Z(o[9208]) );
  AND U2642 ( .A(p_input[29208]), .B(p_input[19208]), .Z(n1762) );
  AND U2643 ( .A(p_input[9208]), .B(p_input[39208]), .Z(n1761) );
  AND U2644 ( .A(n1763), .B(n1764), .Z(o[9207]) );
  AND U2645 ( .A(p_input[29207]), .B(p_input[19207]), .Z(n1764) );
  AND U2646 ( .A(p_input[9207]), .B(p_input[39207]), .Z(n1763) );
  AND U2647 ( .A(n1765), .B(n1766), .Z(o[9206]) );
  AND U2648 ( .A(p_input[29206]), .B(p_input[19206]), .Z(n1766) );
  AND U2649 ( .A(p_input[9206]), .B(p_input[39206]), .Z(n1765) );
  AND U2650 ( .A(n1767), .B(n1768), .Z(o[9205]) );
  AND U2651 ( .A(p_input[29205]), .B(p_input[19205]), .Z(n1768) );
  AND U2652 ( .A(p_input[9205]), .B(p_input[39205]), .Z(n1767) );
  AND U2653 ( .A(n1769), .B(n1770), .Z(o[9204]) );
  AND U2654 ( .A(p_input[29204]), .B(p_input[19204]), .Z(n1770) );
  AND U2655 ( .A(p_input[9204]), .B(p_input[39204]), .Z(n1769) );
  AND U2656 ( .A(n1771), .B(n1772), .Z(o[9203]) );
  AND U2657 ( .A(p_input[29203]), .B(p_input[19203]), .Z(n1772) );
  AND U2658 ( .A(p_input[9203]), .B(p_input[39203]), .Z(n1771) );
  AND U2659 ( .A(n1773), .B(n1774), .Z(o[9202]) );
  AND U2660 ( .A(p_input[29202]), .B(p_input[19202]), .Z(n1774) );
  AND U2661 ( .A(p_input[9202]), .B(p_input[39202]), .Z(n1773) );
  AND U2662 ( .A(n1775), .B(n1776), .Z(o[9201]) );
  AND U2663 ( .A(p_input[29201]), .B(p_input[19201]), .Z(n1776) );
  AND U2664 ( .A(p_input[9201]), .B(p_input[39201]), .Z(n1775) );
  AND U2665 ( .A(n1777), .B(n1778), .Z(o[9200]) );
  AND U2666 ( .A(p_input[29200]), .B(p_input[19200]), .Z(n1778) );
  AND U2667 ( .A(p_input[9200]), .B(p_input[39200]), .Z(n1777) );
  AND U2668 ( .A(n1779), .B(n1780), .Z(o[91]) );
  AND U2669 ( .A(p_input[20091]), .B(p_input[10091]), .Z(n1780) );
  AND U2670 ( .A(p_input[91]), .B(p_input[30091]), .Z(n1779) );
  AND U2671 ( .A(n1781), .B(n1782), .Z(o[919]) );
  AND U2672 ( .A(p_input[20919]), .B(p_input[10919]), .Z(n1782) );
  AND U2673 ( .A(p_input[919]), .B(p_input[30919]), .Z(n1781) );
  AND U2674 ( .A(n1783), .B(n1784), .Z(o[9199]) );
  AND U2675 ( .A(p_input[29199]), .B(p_input[19199]), .Z(n1784) );
  AND U2676 ( .A(p_input[9199]), .B(p_input[39199]), .Z(n1783) );
  AND U2677 ( .A(n1785), .B(n1786), .Z(o[9198]) );
  AND U2678 ( .A(p_input[29198]), .B(p_input[19198]), .Z(n1786) );
  AND U2679 ( .A(p_input[9198]), .B(p_input[39198]), .Z(n1785) );
  AND U2680 ( .A(n1787), .B(n1788), .Z(o[9197]) );
  AND U2681 ( .A(p_input[29197]), .B(p_input[19197]), .Z(n1788) );
  AND U2682 ( .A(p_input[9197]), .B(p_input[39197]), .Z(n1787) );
  AND U2683 ( .A(n1789), .B(n1790), .Z(o[9196]) );
  AND U2684 ( .A(p_input[29196]), .B(p_input[19196]), .Z(n1790) );
  AND U2685 ( .A(p_input[9196]), .B(p_input[39196]), .Z(n1789) );
  AND U2686 ( .A(n1791), .B(n1792), .Z(o[9195]) );
  AND U2687 ( .A(p_input[29195]), .B(p_input[19195]), .Z(n1792) );
  AND U2688 ( .A(p_input[9195]), .B(p_input[39195]), .Z(n1791) );
  AND U2689 ( .A(n1793), .B(n1794), .Z(o[9194]) );
  AND U2690 ( .A(p_input[29194]), .B(p_input[19194]), .Z(n1794) );
  AND U2691 ( .A(p_input[9194]), .B(p_input[39194]), .Z(n1793) );
  AND U2692 ( .A(n1795), .B(n1796), .Z(o[9193]) );
  AND U2693 ( .A(p_input[29193]), .B(p_input[19193]), .Z(n1796) );
  AND U2694 ( .A(p_input[9193]), .B(p_input[39193]), .Z(n1795) );
  AND U2695 ( .A(n1797), .B(n1798), .Z(o[9192]) );
  AND U2696 ( .A(p_input[29192]), .B(p_input[19192]), .Z(n1798) );
  AND U2697 ( .A(p_input[9192]), .B(p_input[39192]), .Z(n1797) );
  AND U2698 ( .A(n1799), .B(n1800), .Z(o[9191]) );
  AND U2699 ( .A(p_input[29191]), .B(p_input[19191]), .Z(n1800) );
  AND U2700 ( .A(p_input[9191]), .B(p_input[39191]), .Z(n1799) );
  AND U2701 ( .A(n1801), .B(n1802), .Z(o[9190]) );
  AND U2702 ( .A(p_input[29190]), .B(p_input[19190]), .Z(n1802) );
  AND U2703 ( .A(p_input[9190]), .B(p_input[39190]), .Z(n1801) );
  AND U2704 ( .A(n1803), .B(n1804), .Z(o[918]) );
  AND U2705 ( .A(p_input[20918]), .B(p_input[10918]), .Z(n1804) );
  AND U2706 ( .A(p_input[918]), .B(p_input[30918]), .Z(n1803) );
  AND U2707 ( .A(n1805), .B(n1806), .Z(o[9189]) );
  AND U2708 ( .A(p_input[29189]), .B(p_input[19189]), .Z(n1806) );
  AND U2709 ( .A(p_input[9189]), .B(p_input[39189]), .Z(n1805) );
  AND U2710 ( .A(n1807), .B(n1808), .Z(o[9188]) );
  AND U2711 ( .A(p_input[29188]), .B(p_input[19188]), .Z(n1808) );
  AND U2712 ( .A(p_input[9188]), .B(p_input[39188]), .Z(n1807) );
  AND U2713 ( .A(n1809), .B(n1810), .Z(o[9187]) );
  AND U2714 ( .A(p_input[29187]), .B(p_input[19187]), .Z(n1810) );
  AND U2715 ( .A(p_input[9187]), .B(p_input[39187]), .Z(n1809) );
  AND U2716 ( .A(n1811), .B(n1812), .Z(o[9186]) );
  AND U2717 ( .A(p_input[29186]), .B(p_input[19186]), .Z(n1812) );
  AND U2718 ( .A(p_input[9186]), .B(p_input[39186]), .Z(n1811) );
  AND U2719 ( .A(n1813), .B(n1814), .Z(o[9185]) );
  AND U2720 ( .A(p_input[29185]), .B(p_input[19185]), .Z(n1814) );
  AND U2721 ( .A(p_input[9185]), .B(p_input[39185]), .Z(n1813) );
  AND U2722 ( .A(n1815), .B(n1816), .Z(o[9184]) );
  AND U2723 ( .A(p_input[29184]), .B(p_input[19184]), .Z(n1816) );
  AND U2724 ( .A(p_input[9184]), .B(p_input[39184]), .Z(n1815) );
  AND U2725 ( .A(n1817), .B(n1818), .Z(o[9183]) );
  AND U2726 ( .A(p_input[29183]), .B(p_input[19183]), .Z(n1818) );
  AND U2727 ( .A(p_input[9183]), .B(p_input[39183]), .Z(n1817) );
  AND U2728 ( .A(n1819), .B(n1820), .Z(o[9182]) );
  AND U2729 ( .A(p_input[29182]), .B(p_input[19182]), .Z(n1820) );
  AND U2730 ( .A(p_input[9182]), .B(p_input[39182]), .Z(n1819) );
  AND U2731 ( .A(n1821), .B(n1822), .Z(o[9181]) );
  AND U2732 ( .A(p_input[29181]), .B(p_input[19181]), .Z(n1822) );
  AND U2733 ( .A(p_input[9181]), .B(p_input[39181]), .Z(n1821) );
  AND U2734 ( .A(n1823), .B(n1824), .Z(o[9180]) );
  AND U2735 ( .A(p_input[29180]), .B(p_input[19180]), .Z(n1824) );
  AND U2736 ( .A(p_input[9180]), .B(p_input[39180]), .Z(n1823) );
  AND U2737 ( .A(n1825), .B(n1826), .Z(o[917]) );
  AND U2738 ( .A(p_input[20917]), .B(p_input[10917]), .Z(n1826) );
  AND U2739 ( .A(p_input[917]), .B(p_input[30917]), .Z(n1825) );
  AND U2740 ( .A(n1827), .B(n1828), .Z(o[9179]) );
  AND U2741 ( .A(p_input[29179]), .B(p_input[19179]), .Z(n1828) );
  AND U2742 ( .A(p_input[9179]), .B(p_input[39179]), .Z(n1827) );
  AND U2743 ( .A(n1829), .B(n1830), .Z(o[9178]) );
  AND U2744 ( .A(p_input[29178]), .B(p_input[19178]), .Z(n1830) );
  AND U2745 ( .A(p_input[9178]), .B(p_input[39178]), .Z(n1829) );
  AND U2746 ( .A(n1831), .B(n1832), .Z(o[9177]) );
  AND U2747 ( .A(p_input[29177]), .B(p_input[19177]), .Z(n1832) );
  AND U2748 ( .A(p_input[9177]), .B(p_input[39177]), .Z(n1831) );
  AND U2749 ( .A(n1833), .B(n1834), .Z(o[9176]) );
  AND U2750 ( .A(p_input[29176]), .B(p_input[19176]), .Z(n1834) );
  AND U2751 ( .A(p_input[9176]), .B(p_input[39176]), .Z(n1833) );
  AND U2752 ( .A(n1835), .B(n1836), .Z(o[9175]) );
  AND U2753 ( .A(p_input[29175]), .B(p_input[19175]), .Z(n1836) );
  AND U2754 ( .A(p_input[9175]), .B(p_input[39175]), .Z(n1835) );
  AND U2755 ( .A(n1837), .B(n1838), .Z(o[9174]) );
  AND U2756 ( .A(p_input[29174]), .B(p_input[19174]), .Z(n1838) );
  AND U2757 ( .A(p_input[9174]), .B(p_input[39174]), .Z(n1837) );
  AND U2758 ( .A(n1839), .B(n1840), .Z(o[9173]) );
  AND U2759 ( .A(p_input[29173]), .B(p_input[19173]), .Z(n1840) );
  AND U2760 ( .A(p_input[9173]), .B(p_input[39173]), .Z(n1839) );
  AND U2761 ( .A(n1841), .B(n1842), .Z(o[9172]) );
  AND U2762 ( .A(p_input[29172]), .B(p_input[19172]), .Z(n1842) );
  AND U2763 ( .A(p_input[9172]), .B(p_input[39172]), .Z(n1841) );
  AND U2764 ( .A(n1843), .B(n1844), .Z(o[9171]) );
  AND U2765 ( .A(p_input[29171]), .B(p_input[19171]), .Z(n1844) );
  AND U2766 ( .A(p_input[9171]), .B(p_input[39171]), .Z(n1843) );
  AND U2767 ( .A(n1845), .B(n1846), .Z(o[9170]) );
  AND U2768 ( .A(p_input[29170]), .B(p_input[19170]), .Z(n1846) );
  AND U2769 ( .A(p_input[9170]), .B(p_input[39170]), .Z(n1845) );
  AND U2770 ( .A(n1847), .B(n1848), .Z(o[916]) );
  AND U2771 ( .A(p_input[20916]), .B(p_input[10916]), .Z(n1848) );
  AND U2772 ( .A(p_input[916]), .B(p_input[30916]), .Z(n1847) );
  AND U2773 ( .A(n1849), .B(n1850), .Z(o[9169]) );
  AND U2774 ( .A(p_input[29169]), .B(p_input[19169]), .Z(n1850) );
  AND U2775 ( .A(p_input[9169]), .B(p_input[39169]), .Z(n1849) );
  AND U2776 ( .A(n1851), .B(n1852), .Z(o[9168]) );
  AND U2777 ( .A(p_input[29168]), .B(p_input[19168]), .Z(n1852) );
  AND U2778 ( .A(p_input[9168]), .B(p_input[39168]), .Z(n1851) );
  AND U2779 ( .A(n1853), .B(n1854), .Z(o[9167]) );
  AND U2780 ( .A(p_input[29167]), .B(p_input[19167]), .Z(n1854) );
  AND U2781 ( .A(p_input[9167]), .B(p_input[39167]), .Z(n1853) );
  AND U2782 ( .A(n1855), .B(n1856), .Z(o[9166]) );
  AND U2783 ( .A(p_input[29166]), .B(p_input[19166]), .Z(n1856) );
  AND U2784 ( .A(p_input[9166]), .B(p_input[39166]), .Z(n1855) );
  AND U2785 ( .A(n1857), .B(n1858), .Z(o[9165]) );
  AND U2786 ( .A(p_input[29165]), .B(p_input[19165]), .Z(n1858) );
  AND U2787 ( .A(p_input[9165]), .B(p_input[39165]), .Z(n1857) );
  AND U2788 ( .A(n1859), .B(n1860), .Z(o[9164]) );
  AND U2789 ( .A(p_input[29164]), .B(p_input[19164]), .Z(n1860) );
  AND U2790 ( .A(p_input[9164]), .B(p_input[39164]), .Z(n1859) );
  AND U2791 ( .A(n1861), .B(n1862), .Z(o[9163]) );
  AND U2792 ( .A(p_input[29163]), .B(p_input[19163]), .Z(n1862) );
  AND U2793 ( .A(p_input[9163]), .B(p_input[39163]), .Z(n1861) );
  AND U2794 ( .A(n1863), .B(n1864), .Z(o[9162]) );
  AND U2795 ( .A(p_input[29162]), .B(p_input[19162]), .Z(n1864) );
  AND U2796 ( .A(p_input[9162]), .B(p_input[39162]), .Z(n1863) );
  AND U2797 ( .A(n1865), .B(n1866), .Z(o[9161]) );
  AND U2798 ( .A(p_input[29161]), .B(p_input[19161]), .Z(n1866) );
  AND U2799 ( .A(p_input[9161]), .B(p_input[39161]), .Z(n1865) );
  AND U2800 ( .A(n1867), .B(n1868), .Z(o[9160]) );
  AND U2801 ( .A(p_input[29160]), .B(p_input[19160]), .Z(n1868) );
  AND U2802 ( .A(p_input[9160]), .B(p_input[39160]), .Z(n1867) );
  AND U2803 ( .A(n1869), .B(n1870), .Z(o[915]) );
  AND U2804 ( .A(p_input[20915]), .B(p_input[10915]), .Z(n1870) );
  AND U2805 ( .A(p_input[915]), .B(p_input[30915]), .Z(n1869) );
  AND U2806 ( .A(n1871), .B(n1872), .Z(o[9159]) );
  AND U2807 ( .A(p_input[29159]), .B(p_input[19159]), .Z(n1872) );
  AND U2808 ( .A(p_input[9159]), .B(p_input[39159]), .Z(n1871) );
  AND U2809 ( .A(n1873), .B(n1874), .Z(o[9158]) );
  AND U2810 ( .A(p_input[29158]), .B(p_input[19158]), .Z(n1874) );
  AND U2811 ( .A(p_input[9158]), .B(p_input[39158]), .Z(n1873) );
  AND U2812 ( .A(n1875), .B(n1876), .Z(o[9157]) );
  AND U2813 ( .A(p_input[29157]), .B(p_input[19157]), .Z(n1876) );
  AND U2814 ( .A(p_input[9157]), .B(p_input[39157]), .Z(n1875) );
  AND U2815 ( .A(n1877), .B(n1878), .Z(o[9156]) );
  AND U2816 ( .A(p_input[29156]), .B(p_input[19156]), .Z(n1878) );
  AND U2817 ( .A(p_input[9156]), .B(p_input[39156]), .Z(n1877) );
  AND U2818 ( .A(n1879), .B(n1880), .Z(o[9155]) );
  AND U2819 ( .A(p_input[29155]), .B(p_input[19155]), .Z(n1880) );
  AND U2820 ( .A(p_input[9155]), .B(p_input[39155]), .Z(n1879) );
  AND U2821 ( .A(n1881), .B(n1882), .Z(o[9154]) );
  AND U2822 ( .A(p_input[29154]), .B(p_input[19154]), .Z(n1882) );
  AND U2823 ( .A(p_input[9154]), .B(p_input[39154]), .Z(n1881) );
  AND U2824 ( .A(n1883), .B(n1884), .Z(o[9153]) );
  AND U2825 ( .A(p_input[29153]), .B(p_input[19153]), .Z(n1884) );
  AND U2826 ( .A(p_input[9153]), .B(p_input[39153]), .Z(n1883) );
  AND U2827 ( .A(n1885), .B(n1886), .Z(o[9152]) );
  AND U2828 ( .A(p_input[29152]), .B(p_input[19152]), .Z(n1886) );
  AND U2829 ( .A(p_input[9152]), .B(p_input[39152]), .Z(n1885) );
  AND U2830 ( .A(n1887), .B(n1888), .Z(o[9151]) );
  AND U2831 ( .A(p_input[29151]), .B(p_input[19151]), .Z(n1888) );
  AND U2832 ( .A(p_input[9151]), .B(p_input[39151]), .Z(n1887) );
  AND U2833 ( .A(n1889), .B(n1890), .Z(o[9150]) );
  AND U2834 ( .A(p_input[29150]), .B(p_input[19150]), .Z(n1890) );
  AND U2835 ( .A(p_input[9150]), .B(p_input[39150]), .Z(n1889) );
  AND U2836 ( .A(n1891), .B(n1892), .Z(o[914]) );
  AND U2837 ( .A(p_input[20914]), .B(p_input[10914]), .Z(n1892) );
  AND U2838 ( .A(p_input[914]), .B(p_input[30914]), .Z(n1891) );
  AND U2839 ( .A(n1893), .B(n1894), .Z(o[9149]) );
  AND U2840 ( .A(p_input[29149]), .B(p_input[19149]), .Z(n1894) );
  AND U2841 ( .A(p_input[9149]), .B(p_input[39149]), .Z(n1893) );
  AND U2842 ( .A(n1895), .B(n1896), .Z(o[9148]) );
  AND U2843 ( .A(p_input[29148]), .B(p_input[19148]), .Z(n1896) );
  AND U2844 ( .A(p_input[9148]), .B(p_input[39148]), .Z(n1895) );
  AND U2845 ( .A(n1897), .B(n1898), .Z(o[9147]) );
  AND U2846 ( .A(p_input[29147]), .B(p_input[19147]), .Z(n1898) );
  AND U2847 ( .A(p_input[9147]), .B(p_input[39147]), .Z(n1897) );
  AND U2848 ( .A(n1899), .B(n1900), .Z(o[9146]) );
  AND U2849 ( .A(p_input[29146]), .B(p_input[19146]), .Z(n1900) );
  AND U2850 ( .A(p_input[9146]), .B(p_input[39146]), .Z(n1899) );
  AND U2851 ( .A(n1901), .B(n1902), .Z(o[9145]) );
  AND U2852 ( .A(p_input[29145]), .B(p_input[19145]), .Z(n1902) );
  AND U2853 ( .A(p_input[9145]), .B(p_input[39145]), .Z(n1901) );
  AND U2854 ( .A(n1903), .B(n1904), .Z(o[9144]) );
  AND U2855 ( .A(p_input[29144]), .B(p_input[19144]), .Z(n1904) );
  AND U2856 ( .A(p_input[9144]), .B(p_input[39144]), .Z(n1903) );
  AND U2857 ( .A(n1905), .B(n1906), .Z(o[9143]) );
  AND U2858 ( .A(p_input[29143]), .B(p_input[19143]), .Z(n1906) );
  AND U2859 ( .A(p_input[9143]), .B(p_input[39143]), .Z(n1905) );
  AND U2860 ( .A(n1907), .B(n1908), .Z(o[9142]) );
  AND U2861 ( .A(p_input[29142]), .B(p_input[19142]), .Z(n1908) );
  AND U2862 ( .A(p_input[9142]), .B(p_input[39142]), .Z(n1907) );
  AND U2863 ( .A(n1909), .B(n1910), .Z(o[9141]) );
  AND U2864 ( .A(p_input[29141]), .B(p_input[19141]), .Z(n1910) );
  AND U2865 ( .A(p_input[9141]), .B(p_input[39141]), .Z(n1909) );
  AND U2866 ( .A(n1911), .B(n1912), .Z(o[9140]) );
  AND U2867 ( .A(p_input[29140]), .B(p_input[19140]), .Z(n1912) );
  AND U2868 ( .A(p_input[9140]), .B(p_input[39140]), .Z(n1911) );
  AND U2869 ( .A(n1913), .B(n1914), .Z(o[913]) );
  AND U2870 ( .A(p_input[20913]), .B(p_input[10913]), .Z(n1914) );
  AND U2871 ( .A(p_input[913]), .B(p_input[30913]), .Z(n1913) );
  AND U2872 ( .A(n1915), .B(n1916), .Z(o[9139]) );
  AND U2873 ( .A(p_input[29139]), .B(p_input[19139]), .Z(n1916) );
  AND U2874 ( .A(p_input[9139]), .B(p_input[39139]), .Z(n1915) );
  AND U2875 ( .A(n1917), .B(n1918), .Z(o[9138]) );
  AND U2876 ( .A(p_input[29138]), .B(p_input[19138]), .Z(n1918) );
  AND U2877 ( .A(p_input[9138]), .B(p_input[39138]), .Z(n1917) );
  AND U2878 ( .A(n1919), .B(n1920), .Z(o[9137]) );
  AND U2879 ( .A(p_input[29137]), .B(p_input[19137]), .Z(n1920) );
  AND U2880 ( .A(p_input[9137]), .B(p_input[39137]), .Z(n1919) );
  AND U2881 ( .A(n1921), .B(n1922), .Z(o[9136]) );
  AND U2882 ( .A(p_input[29136]), .B(p_input[19136]), .Z(n1922) );
  AND U2883 ( .A(p_input[9136]), .B(p_input[39136]), .Z(n1921) );
  AND U2884 ( .A(n1923), .B(n1924), .Z(o[9135]) );
  AND U2885 ( .A(p_input[29135]), .B(p_input[19135]), .Z(n1924) );
  AND U2886 ( .A(p_input[9135]), .B(p_input[39135]), .Z(n1923) );
  AND U2887 ( .A(n1925), .B(n1926), .Z(o[9134]) );
  AND U2888 ( .A(p_input[29134]), .B(p_input[19134]), .Z(n1926) );
  AND U2889 ( .A(p_input[9134]), .B(p_input[39134]), .Z(n1925) );
  AND U2890 ( .A(n1927), .B(n1928), .Z(o[9133]) );
  AND U2891 ( .A(p_input[29133]), .B(p_input[19133]), .Z(n1928) );
  AND U2892 ( .A(p_input[9133]), .B(p_input[39133]), .Z(n1927) );
  AND U2893 ( .A(n1929), .B(n1930), .Z(o[9132]) );
  AND U2894 ( .A(p_input[29132]), .B(p_input[19132]), .Z(n1930) );
  AND U2895 ( .A(p_input[9132]), .B(p_input[39132]), .Z(n1929) );
  AND U2896 ( .A(n1931), .B(n1932), .Z(o[9131]) );
  AND U2897 ( .A(p_input[29131]), .B(p_input[19131]), .Z(n1932) );
  AND U2898 ( .A(p_input[9131]), .B(p_input[39131]), .Z(n1931) );
  AND U2899 ( .A(n1933), .B(n1934), .Z(o[9130]) );
  AND U2900 ( .A(p_input[29130]), .B(p_input[19130]), .Z(n1934) );
  AND U2901 ( .A(p_input[9130]), .B(p_input[39130]), .Z(n1933) );
  AND U2902 ( .A(n1935), .B(n1936), .Z(o[912]) );
  AND U2903 ( .A(p_input[20912]), .B(p_input[10912]), .Z(n1936) );
  AND U2904 ( .A(p_input[912]), .B(p_input[30912]), .Z(n1935) );
  AND U2905 ( .A(n1937), .B(n1938), .Z(o[9129]) );
  AND U2906 ( .A(p_input[29129]), .B(p_input[19129]), .Z(n1938) );
  AND U2907 ( .A(p_input[9129]), .B(p_input[39129]), .Z(n1937) );
  AND U2908 ( .A(n1939), .B(n1940), .Z(o[9128]) );
  AND U2909 ( .A(p_input[29128]), .B(p_input[19128]), .Z(n1940) );
  AND U2910 ( .A(p_input[9128]), .B(p_input[39128]), .Z(n1939) );
  AND U2911 ( .A(n1941), .B(n1942), .Z(o[9127]) );
  AND U2912 ( .A(p_input[29127]), .B(p_input[19127]), .Z(n1942) );
  AND U2913 ( .A(p_input[9127]), .B(p_input[39127]), .Z(n1941) );
  AND U2914 ( .A(n1943), .B(n1944), .Z(o[9126]) );
  AND U2915 ( .A(p_input[29126]), .B(p_input[19126]), .Z(n1944) );
  AND U2916 ( .A(p_input[9126]), .B(p_input[39126]), .Z(n1943) );
  AND U2917 ( .A(n1945), .B(n1946), .Z(o[9125]) );
  AND U2918 ( .A(p_input[29125]), .B(p_input[19125]), .Z(n1946) );
  AND U2919 ( .A(p_input[9125]), .B(p_input[39125]), .Z(n1945) );
  AND U2920 ( .A(n1947), .B(n1948), .Z(o[9124]) );
  AND U2921 ( .A(p_input[29124]), .B(p_input[19124]), .Z(n1948) );
  AND U2922 ( .A(p_input[9124]), .B(p_input[39124]), .Z(n1947) );
  AND U2923 ( .A(n1949), .B(n1950), .Z(o[9123]) );
  AND U2924 ( .A(p_input[29123]), .B(p_input[19123]), .Z(n1950) );
  AND U2925 ( .A(p_input[9123]), .B(p_input[39123]), .Z(n1949) );
  AND U2926 ( .A(n1951), .B(n1952), .Z(o[9122]) );
  AND U2927 ( .A(p_input[29122]), .B(p_input[19122]), .Z(n1952) );
  AND U2928 ( .A(p_input[9122]), .B(p_input[39122]), .Z(n1951) );
  AND U2929 ( .A(n1953), .B(n1954), .Z(o[9121]) );
  AND U2930 ( .A(p_input[29121]), .B(p_input[19121]), .Z(n1954) );
  AND U2931 ( .A(p_input[9121]), .B(p_input[39121]), .Z(n1953) );
  AND U2932 ( .A(n1955), .B(n1956), .Z(o[9120]) );
  AND U2933 ( .A(p_input[29120]), .B(p_input[19120]), .Z(n1956) );
  AND U2934 ( .A(p_input[9120]), .B(p_input[39120]), .Z(n1955) );
  AND U2935 ( .A(n1957), .B(n1958), .Z(o[911]) );
  AND U2936 ( .A(p_input[20911]), .B(p_input[10911]), .Z(n1958) );
  AND U2937 ( .A(p_input[911]), .B(p_input[30911]), .Z(n1957) );
  AND U2938 ( .A(n1959), .B(n1960), .Z(o[9119]) );
  AND U2939 ( .A(p_input[29119]), .B(p_input[19119]), .Z(n1960) );
  AND U2940 ( .A(p_input[9119]), .B(p_input[39119]), .Z(n1959) );
  AND U2941 ( .A(n1961), .B(n1962), .Z(o[9118]) );
  AND U2942 ( .A(p_input[29118]), .B(p_input[19118]), .Z(n1962) );
  AND U2943 ( .A(p_input[9118]), .B(p_input[39118]), .Z(n1961) );
  AND U2944 ( .A(n1963), .B(n1964), .Z(o[9117]) );
  AND U2945 ( .A(p_input[29117]), .B(p_input[19117]), .Z(n1964) );
  AND U2946 ( .A(p_input[9117]), .B(p_input[39117]), .Z(n1963) );
  AND U2947 ( .A(n1965), .B(n1966), .Z(o[9116]) );
  AND U2948 ( .A(p_input[29116]), .B(p_input[19116]), .Z(n1966) );
  AND U2949 ( .A(p_input[9116]), .B(p_input[39116]), .Z(n1965) );
  AND U2950 ( .A(n1967), .B(n1968), .Z(o[9115]) );
  AND U2951 ( .A(p_input[29115]), .B(p_input[19115]), .Z(n1968) );
  AND U2952 ( .A(p_input[9115]), .B(p_input[39115]), .Z(n1967) );
  AND U2953 ( .A(n1969), .B(n1970), .Z(o[9114]) );
  AND U2954 ( .A(p_input[29114]), .B(p_input[19114]), .Z(n1970) );
  AND U2955 ( .A(p_input[9114]), .B(p_input[39114]), .Z(n1969) );
  AND U2956 ( .A(n1971), .B(n1972), .Z(o[9113]) );
  AND U2957 ( .A(p_input[29113]), .B(p_input[19113]), .Z(n1972) );
  AND U2958 ( .A(p_input[9113]), .B(p_input[39113]), .Z(n1971) );
  AND U2959 ( .A(n1973), .B(n1974), .Z(o[9112]) );
  AND U2960 ( .A(p_input[29112]), .B(p_input[19112]), .Z(n1974) );
  AND U2961 ( .A(p_input[9112]), .B(p_input[39112]), .Z(n1973) );
  AND U2962 ( .A(n1975), .B(n1976), .Z(o[9111]) );
  AND U2963 ( .A(p_input[29111]), .B(p_input[19111]), .Z(n1976) );
  AND U2964 ( .A(p_input[9111]), .B(p_input[39111]), .Z(n1975) );
  AND U2965 ( .A(n1977), .B(n1978), .Z(o[9110]) );
  AND U2966 ( .A(p_input[29110]), .B(p_input[19110]), .Z(n1978) );
  AND U2967 ( .A(p_input[9110]), .B(p_input[39110]), .Z(n1977) );
  AND U2968 ( .A(n1979), .B(n1980), .Z(o[910]) );
  AND U2969 ( .A(p_input[20910]), .B(p_input[10910]), .Z(n1980) );
  AND U2970 ( .A(p_input[910]), .B(p_input[30910]), .Z(n1979) );
  AND U2971 ( .A(n1981), .B(n1982), .Z(o[9109]) );
  AND U2972 ( .A(p_input[29109]), .B(p_input[19109]), .Z(n1982) );
  AND U2973 ( .A(p_input[9109]), .B(p_input[39109]), .Z(n1981) );
  AND U2974 ( .A(n1983), .B(n1984), .Z(o[9108]) );
  AND U2975 ( .A(p_input[29108]), .B(p_input[19108]), .Z(n1984) );
  AND U2976 ( .A(p_input[9108]), .B(p_input[39108]), .Z(n1983) );
  AND U2977 ( .A(n1985), .B(n1986), .Z(o[9107]) );
  AND U2978 ( .A(p_input[29107]), .B(p_input[19107]), .Z(n1986) );
  AND U2979 ( .A(p_input[9107]), .B(p_input[39107]), .Z(n1985) );
  AND U2980 ( .A(n1987), .B(n1988), .Z(o[9106]) );
  AND U2981 ( .A(p_input[29106]), .B(p_input[19106]), .Z(n1988) );
  AND U2982 ( .A(p_input[9106]), .B(p_input[39106]), .Z(n1987) );
  AND U2983 ( .A(n1989), .B(n1990), .Z(o[9105]) );
  AND U2984 ( .A(p_input[29105]), .B(p_input[19105]), .Z(n1990) );
  AND U2985 ( .A(p_input[9105]), .B(p_input[39105]), .Z(n1989) );
  AND U2986 ( .A(n1991), .B(n1992), .Z(o[9104]) );
  AND U2987 ( .A(p_input[29104]), .B(p_input[19104]), .Z(n1992) );
  AND U2988 ( .A(p_input[9104]), .B(p_input[39104]), .Z(n1991) );
  AND U2989 ( .A(n1993), .B(n1994), .Z(o[9103]) );
  AND U2990 ( .A(p_input[29103]), .B(p_input[19103]), .Z(n1994) );
  AND U2991 ( .A(p_input[9103]), .B(p_input[39103]), .Z(n1993) );
  AND U2992 ( .A(n1995), .B(n1996), .Z(o[9102]) );
  AND U2993 ( .A(p_input[29102]), .B(p_input[19102]), .Z(n1996) );
  AND U2994 ( .A(p_input[9102]), .B(p_input[39102]), .Z(n1995) );
  AND U2995 ( .A(n1997), .B(n1998), .Z(o[9101]) );
  AND U2996 ( .A(p_input[29101]), .B(p_input[19101]), .Z(n1998) );
  AND U2997 ( .A(p_input[9101]), .B(p_input[39101]), .Z(n1997) );
  AND U2998 ( .A(n1999), .B(n2000), .Z(o[9100]) );
  AND U2999 ( .A(p_input[29100]), .B(p_input[19100]), .Z(n2000) );
  AND U3000 ( .A(p_input[9100]), .B(p_input[39100]), .Z(n1999) );
  AND U3001 ( .A(n2001), .B(n2002), .Z(o[90]) );
  AND U3002 ( .A(p_input[20090]), .B(p_input[10090]), .Z(n2002) );
  AND U3003 ( .A(p_input[90]), .B(p_input[30090]), .Z(n2001) );
  AND U3004 ( .A(n2003), .B(n2004), .Z(o[909]) );
  AND U3005 ( .A(p_input[20909]), .B(p_input[10909]), .Z(n2004) );
  AND U3006 ( .A(p_input[909]), .B(p_input[30909]), .Z(n2003) );
  AND U3007 ( .A(n2005), .B(n2006), .Z(o[9099]) );
  AND U3008 ( .A(p_input[29099]), .B(p_input[19099]), .Z(n2006) );
  AND U3009 ( .A(p_input[9099]), .B(p_input[39099]), .Z(n2005) );
  AND U3010 ( .A(n2007), .B(n2008), .Z(o[9098]) );
  AND U3011 ( .A(p_input[29098]), .B(p_input[19098]), .Z(n2008) );
  AND U3012 ( .A(p_input[9098]), .B(p_input[39098]), .Z(n2007) );
  AND U3013 ( .A(n2009), .B(n2010), .Z(o[9097]) );
  AND U3014 ( .A(p_input[29097]), .B(p_input[19097]), .Z(n2010) );
  AND U3015 ( .A(p_input[9097]), .B(p_input[39097]), .Z(n2009) );
  AND U3016 ( .A(n2011), .B(n2012), .Z(o[9096]) );
  AND U3017 ( .A(p_input[29096]), .B(p_input[19096]), .Z(n2012) );
  AND U3018 ( .A(p_input[9096]), .B(p_input[39096]), .Z(n2011) );
  AND U3019 ( .A(n2013), .B(n2014), .Z(o[9095]) );
  AND U3020 ( .A(p_input[29095]), .B(p_input[19095]), .Z(n2014) );
  AND U3021 ( .A(p_input[9095]), .B(p_input[39095]), .Z(n2013) );
  AND U3022 ( .A(n2015), .B(n2016), .Z(o[9094]) );
  AND U3023 ( .A(p_input[29094]), .B(p_input[19094]), .Z(n2016) );
  AND U3024 ( .A(p_input[9094]), .B(p_input[39094]), .Z(n2015) );
  AND U3025 ( .A(n2017), .B(n2018), .Z(o[9093]) );
  AND U3026 ( .A(p_input[29093]), .B(p_input[19093]), .Z(n2018) );
  AND U3027 ( .A(p_input[9093]), .B(p_input[39093]), .Z(n2017) );
  AND U3028 ( .A(n2019), .B(n2020), .Z(o[9092]) );
  AND U3029 ( .A(p_input[29092]), .B(p_input[19092]), .Z(n2020) );
  AND U3030 ( .A(p_input[9092]), .B(p_input[39092]), .Z(n2019) );
  AND U3031 ( .A(n2021), .B(n2022), .Z(o[9091]) );
  AND U3032 ( .A(p_input[29091]), .B(p_input[19091]), .Z(n2022) );
  AND U3033 ( .A(p_input[9091]), .B(p_input[39091]), .Z(n2021) );
  AND U3034 ( .A(n2023), .B(n2024), .Z(o[9090]) );
  AND U3035 ( .A(p_input[29090]), .B(p_input[19090]), .Z(n2024) );
  AND U3036 ( .A(p_input[9090]), .B(p_input[39090]), .Z(n2023) );
  AND U3037 ( .A(n2025), .B(n2026), .Z(o[908]) );
  AND U3038 ( .A(p_input[20908]), .B(p_input[10908]), .Z(n2026) );
  AND U3039 ( .A(p_input[908]), .B(p_input[30908]), .Z(n2025) );
  AND U3040 ( .A(n2027), .B(n2028), .Z(o[9089]) );
  AND U3041 ( .A(p_input[29089]), .B(p_input[19089]), .Z(n2028) );
  AND U3042 ( .A(p_input[9089]), .B(p_input[39089]), .Z(n2027) );
  AND U3043 ( .A(n2029), .B(n2030), .Z(o[9088]) );
  AND U3044 ( .A(p_input[29088]), .B(p_input[19088]), .Z(n2030) );
  AND U3045 ( .A(p_input[9088]), .B(p_input[39088]), .Z(n2029) );
  AND U3046 ( .A(n2031), .B(n2032), .Z(o[9087]) );
  AND U3047 ( .A(p_input[29087]), .B(p_input[19087]), .Z(n2032) );
  AND U3048 ( .A(p_input[9087]), .B(p_input[39087]), .Z(n2031) );
  AND U3049 ( .A(n2033), .B(n2034), .Z(o[9086]) );
  AND U3050 ( .A(p_input[29086]), .B(p_input[19086]), .Z(n2034) );
  AND U3051 ( .A(p_input[9086]), .B(p_input[39086]), .Z(n2033) );
  AND U3052 ( .A(n2035), .B(n2036), .Z(o[9085]) );
  AND U3053 ( .A(p_input[29085]), .B(p_input[19085]), .Z(n2036) );
  AND U3054 ( .A(p_input[9085]), .B(p_input[39085]), .Z(n2035) );
  AND U3055 ( .A(n2037), .B(n2038), .Z(o[9084]) );
  AND U3056 ( .A(p_input[29084]), .B(p_input[19084]), .Z(n2038) );
  AND U3057 ( .A(p_input[9084]), .B(p_input[39084]), .Z(n2037) );
  AND U3058 ( .A(n2039), .B(n2040), .Z(o[9083]) );
  AND U3059 ( .A(p_input[29083]), .B(p_input[19083]), .Z(n2040) );
  AND U3060 ( .A(p_input[9083]), .B(p_input[39083]), .Z(n2039) );
  AND U3061 ( .A(n2041), .B(n2042), .Z(o[9082]) );
  AND U3062 ( .A(p_input[29082]), .B(p_input[19082]), .Z(n2042) );
  AND U3063 ( .A(p_input[9082]), .B(p_input[39082]), .Z(n2041) );
  AND U3064 ( .A(n2043), .B(n2044), .Z(o[9081]) );
  AND U3065 ( .A(p_input[29081]), .B(p_input[19081]), .Z(n2044) );
  AND U3066 ( .A(p_input[9081]), .B(p_input[39081]), .Z(n2043) );
  AND U3067 ( .A(n2045), .B(n2046), .Z(o[9080]) );
  AND U3068 ( .A(p_input[29080]), .B(p_input[19080]), .Z(n2046) );
  AND U3069 ( .A(p_input[9080]), .B(p_input[39080]), .Z(n2045) );
  AND U3070 ( .A(n2047), .B(n2048), .Z(o[907]) );
  AND U3071 ( .A(p_input[20907]), .B(p_input[10907]), .Z(n2048) );
  AND U3072 ( .A(p_input[907]), .B(p_input[30907]), .Z(n2047) );
  AND U3073 ( .A(n2049), .B(n2050), .Z(o[9079]) );
  AND U3074 ( .A(p_input[29079]), .B(p_input[19079]), .Z(n2050) );
  AND U3075 ( .A(p_input[9079]), .B(p_input[39079]), .Z(n2049) );
  AND U3076 ( .A(n2051), .B(n2052), .Z(o[9078]) );
  AND U3077 ( .A(p_input[29078]), .B(p_input[19078]), .Z(n2052) );
  AND U3078 ( .A(p_input[9078]), .B(p_input[39078]), .Z(n2051) );
  AND U3079 ( .A(n2053), .B(n2054), .Z(o[9077]) );
  AND U3080 ( .A(p_input[29077]), .B(p_input[19077]), .Z(n2054) );
  AND U3081 ( .A(p_input[9077]), .B(p_input[39077]), .Z(n2053) );
  AND U3082 ( .A(n2055), .B(n2056), .Z(o[9076]) );
  AND U3083 ( .A(p_input[29076]), .B(p_input[19076]), .Z(n2056) );
  AND U3084 ( .A(p_input[9076]), .B(p_input[39076]), .Z(n2055) );
  AND U3085 ( .A(n2057), .B(n2058), .Z(o[9075]) );
  AND U3086 ( .A(p_input[29075]), .B(p_input[19075]), .Z(n2058) );
  AND U3087 ( .A(p_input[9075]), .B(p_input[39075]), .Z(n2057) );
  AND U3088 ( .A(n2059), .B(n2060), .Z(o[9074]) );
  AND U3089 ( .A(p_input[29074]), .B(p_input[19074]), .Z(n2060) );
  AND U3090 ( .A(p_input[9074]), .B(p_input[39074]), .Z(n2059) );
  AND U3091 ( .A(n2061), .B(n2062), .Z(o[9073]) );
  AND U3092 ( .A(p_input[29073]), .B(p_input[19073]), .Z(n2062) );
  AND U3093 ( .A(p_input[9073]), .B(p_input[39073]), .Z(n2061) );
  AND U3094 ( .A(n2063), .B(n2064), .Z(o[9072]) );
  AND U3095 ( .A(p_input[29072]), .B(p_input[19072]), .Z(n2064) );
  AND U3096 ( .A(p_input[9072]), .B(p_input[39072]), .Z(n2063) );
  AND U3097 ( .A(n2065), .B(n2066), .Z(o[9071]) );
  AND U3098 ( .A(p_input[29071]), .B(p_input[19071]), .Z(n2066) );
  AND U3099 ( .A(p_input[9071]), .B(p_input[39071]), .Z(n2065) );
  AND U3100 ( .A(n2067), .B(n2068), .Z(o[9070]) );
  AND U3101 ( .A(p_input[29070]), .B(p_input[19070]), .Z(n2068) );
  AND U3102 ( .A(p_input[9070]), .B(p_input[39070]), .Z(n2067) );
  AND U3103 ( .A(n2069), .B(n2070), .Z(o[906]) );
  AND U3104 ( .A(p_input[20906]), .B(p_input[10906]), .Z(n2070) );
  AND U3105 ( .A(p_input[906]), .B(p_input[30906]), .Z(n2069) );
  AND U3106 ( .A(n2071), .B(n2072), .Z(o[9069]) );
  AND U3107 ( .A(p_input[29069]), .B(p_input[19069]), .Z(n2072) );
  AND U3108 ( .A(p_input[9069]), .B(p_input[39069]), .Z(n2071) );
  AND U3109 ( .A(n2073), .B(n2074), .Z(o[9068]) );
  AND U3110 ( .A(p_input[29068]), .B(p_input[19068]), .Z(n2074) );
  AND U3111 ( .A(p_input[9068]), .B(p_input[39068]), .Z(n2073) );
  AND U3112 ( .A(n2075), .B(n2076), .Z(o[9067]) );
  AND U3113 ( .A(p_input[29067]), .B(p_input[19067]), .Z(n2076) );
  AND U3114 ( .A(p_input[9067]), .B(p_input[39067]), .Z(n2075) );
  AND U3115 ( .A(n2077), .B(n2078), .Z(o[9066]) );
  AND U3116 ( .A(p_input[29066]), .B(p_input[19066]), .Z(n2078) );
  AND U3117 ( .A(p_input[9066]), .B(p_input[39066]), .Z(n2077) );
  AND U3118 ( .A(n2079), .B(n2080), .Z(o[9065]) );
  AND U3119 ( .A(p_input[29065]), .B(p_input[19065]), .Z(n2080) );
  AND U3120 ( .A(p_input[9065]), .B(p_input[39065]), .Z(n2079) );
  AND U3121 ( .A(n2081), .B(n2082), .Z(o[9064]) );
  AND U3122 ( .A(p_input[29064]), .B(p_input[19064]), .Z(n2082) );
  AND U3123 ( .A(p_input[9064]), .B(p_input[39064]), .Z(n2081) );
  AND U3124 ( .A(n2083), .B(n2084), .Z(o[9063]) );
  AND U3125 ( .A(p_input[29063]), .B(p_input[19063]), .Z(n2084) );
  AND U3126 ( .A(p_input[9063]), .B(p_input[39063]), .Z(n2083) );
  AND U3127 ( .A(n2085), .B(n2086), .Z(o[9062]) );
  AND U3128 ( .A(p_input[29062]), .B(p_input[19062]), .Z(n2086) );
  AND U3129 ( .A(p_input[9062]), .B(p_input[39062]), .Z(n2085) );
  AND U3130 ( .A(n2087), .B(n2088), .Z(o[9061]) );
  AND U3131 ( .A(p_input[29061]), .B(p_input[19061]), .Z(n2088) );
  AND U3132 ( .A(p_input[9061]), .B(p_input[39061]), .Z(n2087) );
  AND U3133 ( .A(n2089), .B(n2090), .Z(o[9060]) );
  AND U3134 ( .A(p_input[29060]), .B(p_input[19060]), .Z(n2090) );
  AND U3135 ( .A(p_input[9060]), .B(p_input[39060]), .Z(n2089) );
  AND U3136 ( .A(n2091), .B(n2092), .Z(o[905]) );
  AND U3137 ( .A(p_input[20905]), .B(p_input[10905]), .Z(n2092) );
  AND U3138 ( .A(p_input[905]), .B(p_input[30905]), .Z(n2091) );
  AND U3139 ( .A(n2093), .B(n2094), .Z(o[9059]) );
  AND U3140 ( .A(p_input[29059]), .B(p_input[19059]), .Z(n2094) );
  AND U3141 ( .A(p_input[9059]), .B(p_input[39059]), .Z(n2093) );
  AND U3142 ( .A(n2095), .B(n2096), .Z(o[9058]) );
  AND U3143 ( .A(p_input[29058]), .B(p_input[19058]), .Z(n2096) );
  AND U3144 ( .A(p_input[9058]), .B(p_input[39058]), .Z(n2095) );
  AND U3145 ( .A(n2097), .B(n2098), .Z(o[9057]) );
  AND U3146 ( .A(p_input[29057]), .B(p_input[19057]), .Z(n2098) );
  AND U3147 ( .A(p_input[9057]), .B(p_input[39057]), .Z(n2097) );
  AND U3148 ( .A(n2099), .B(n2100), .Z(o[9056]) );
  AND U3149 ( .A(p_input[29056]), .B(p_input[19056]), .Z(n2100) );
  AND U3150 ( .A(p_input[9056]), .B(p_input[39056]), .Z(n2099) );
  AND U3151 ( .A(n2101), .B(n2102), .Z(o[9055]) );
  AND U3152 ( .A(p_input[29055]), .B(p_input[19055]), .Z(n2102) );
  AND U3153 ( .A(p_input[9055]), .B(p_input[39055]), .Z(n2101) );
  AND U3154 ( .A(n2103), .B(n2104), .Z(o[9054]) );
  AND U3155 ( .A(p_input[29054]), .B(p_input[19054]), .Z(n2104) );
  AND U3156 ( .A(p_input[9054]), .B(p_input[39054]), .Z(n2103) );
  AND U3157 ( .A(n2105), .B(n2106), .Z(o[9053]) );
  AND U3158 ( .A(p_input[29053]), .B(p_input[19053]), .Z(n2106) );
  AND U3159 ( .A(p_input[9053]), .B(p_input[39053]), .Z(n2105) );
  AND U3160 ( .A(n2107), .B(n2108), .Z(o[9052]) );
  AND U3161 ( .A(p_input[29052]), .B(p_input[19052]), .Z(n2108) );
  AND U3162 ( .A(p_input[9052]), .B(p_input[39052]), .Z(n2107) );
  AND U3163 ( .A(n2109), .B(n2110), .Z(o[9051]) );
  AND U3164 ( .A(p_input[29051]), .B(p_input[19051]), .Z(n2110) );
  AND U3165 ( .A(p_input[9051]), .B(p_input[39051]), .Z(n2109) );
  AND U3166 ( .A(n2111), .B(n2112), .Z(o[9050]) );
  AND U3167 ( .A(p_input[29050]), .B(p_input[19050]), .Z(n2112) );
  AND U3168 ( .A(p_input[9050]), .B(p_input[39050]), .Z(n2111) );
  AND U3169 ( .A(n2113), .B(n2114), .Z(o[904]) );
  AND U3170 ( .A(p_input[20904]), .B(p_input[10904]), .Z(n2114) );
  AND U3171 ( .A(p_input[904]), .B(p_input[30904]), .Z(n2113) );
  AND U3172 ( .A(n2115), .B(n2116), .Z(o[9049]) );
  AND U3173 ( .A(p_input[29049]), .B(p_input[19049]), .Z(n2116) );
  AND U3174 ( .A(p_input[9049]), .B(p_input[39049]), .Z(n2115) );
  AND U3175 ( .A(n2117), .B(n2118), .Z(o[9048]) );
  AND U3176 ( .A(p_input[29048]), .B(p_input[19048]), .Z(n2118) );
  AND U3177 ( .A(p_input[9048]), .B(p_input[39048]), .Z(n2117) );
  AND U3178 ( .A(n2119), .B(n2120), .Z(o[9047]) );
  AND U3179 ( .A(p_input[29047]), .B(p_input[19047]), .Z(n2120) );
  AND U3180 ( .A(p_input[9047]), .B(p_input[39047]), .Z(n2119) );
  AND U3181 ( .A(n2121), .B(n2122), .Z(o[9046]) );
  AND U3182 ( .A(p_input[29046]), .B(p_input[19046]), .Z(n2122) );
  AND U3183 ( .A(p_input[9046]), .B(p_input[39046]), .Z(n2121) );
  AND U3184 ( .A(n2123), .B(n2124), .Z(o[9045]) );
  AND U3185 ( .A(p_input[29045]), .B(p_input[19045]), .Z(n2124) );
  AND U3186 ( .A(p_input[9045]), .B(p_input[39045]), .Z(n2123) );
  AND U3187 ( .A(n2125), .B(n2126), .Z(o[9044]) );
  AND U3188 ( .A(p_input[29044]), .B(p_input[19044]), .Z(n2126) );
  AND U3189 ( .A(p_input[9044]), .B(p_input[39044]), .Z(n2125) );
  AND U3190 ( .A(n2127), .B(n2128), .Z(o[9043]) );
  AND U3191 ( .A(p_input[29043]), .B(p_input[19043]), .Z(n2128) );
  AND U3192 ( .A(p_input[9043]), .B(p_input[39043]), .Z(n2127) );
  AND U3193 ( .A(n2129), .B(n2130), .Z(o[9042]) );
  AND U3194 ( .A(p_input[29042]), .B(p_input[19042]), .Z(n2130) );
  AND U3195 ( .A(p_input[9042]), .B(p_input[39042]), .Z(n2129) );
  AND U3196 ( .A(n2131), .B(n2132), .Z(o[9041]) );
  AND U3197 ( .A(p_input[29041]), .B(p_input[19041]), .Z(n2132) );
  AND U3198 ( .A(p_input[9041]), .B(p_input[39041]), .Z(n2131) );
  AND U3199 ( .A(n2133), .B(n2134), .Z(o[9040]) );
  AND U3200 ( .A(p_input[29040]), .B(p_input[19040]), .Z(n2134) );
  AND U3201 ( .A(p_input[9040]), .B(p_input[39040]), .Z(n2133) );
  AND U3202 ( .A(n2135), .B(n2136), .Z(o[903]) );
  AND U3203 ( .A(p_input[20903]), .B(p_input[10903]), .Z(n2136) );
  AND U3204 ( .A(p_input[903]), .B(p_input[30903]), .Z(n2135) );
  AND U3205 ( .A(n2137), .B(n2138), .Z(o[9039]) );
  AND U3206 ( .A(p_input[29039]), .B(p_input[19039]), .Z(n2138) );
  AND U3207 ( .A(p_input[9039]), .B(p_input[39039]), .Z(n2137) );
  AND U3208 ( .A(n2139), .B(n2140), .Z(o[9038]) );
  AND U3209 ( .A(p_input[29038]), .B(p_input[19038]), .Z(n2140) );
  AND U3210 ( .A(p_input[9038]), .B(p_input[39038]), .Z(n2139) );
  AND U3211 ( .A(n2141), .B(n2142), .Z(o[9037]) );
  AND U3212 ( .A(p_input[29037]), .B(p_input[19037]), .Z(n2142) );
  AND U3213 ( .A(p_input[9037]), .B(p_input[39037]), .Z(n2141) );
  AND U3214 ( .A(n2143), .B(n2144), .Z(o[9036]) );
  AND U3215 ( .A(p_input[29036]), .B(p_input[19036]), .Z(n2144) );
  AND U3216 ( .A(p_input[9036]), .B(p_input[39036]), .Z(n2143) );
  AND U3217 ( .A(n2145), .B(n2146), .Z(o[9035]) );
  AND U3218 ( .A(p_input[29035]), .B(p_input[19035]), .Z(n2146) );
  AND U3219 ( .A(p_input[9035]), .B(p_input[39035]), .Z(n2145) );
  AND U3220 ( .A(n2147), .B(n2148), .Z(o[9034]) );
  AND U3221 ( .A(p_input[29034]), .B(p_input[19034]), .Z(n2148) );
  AND U3222 ( .A(p_input[9034]), .B(p_input[39034]), .Z(n2147) );
  AND U3223 ( .A(n2149), .B(n2150), .Z(o[9033]) );
  AND U3224 ( .A(p_input[29033]), .B(p_input[19033]), .Z(n2150) );
  AND U3225 ( .A(p_input[9033]), .B(p_input[39033]), .Z(n2149) );
  AND U3226 ( .A(n2151), .B(n2152), .Z(o[9032]) );
  AND U3227 ( .A(p_input[29032]), .B(p_input[19032]), .Z(n2152) );
  AND U3228 ( .A(p_input[9032]), .B(p_input[39032]), .Z(n2151) );
  AND U3229 ( .A(n2153), .B(n2154), .Z(o[9031]) );
  AND U3230 ( .A(p_input[29031]), .B(p_input[19031]), .Z(n2154) );
  AND U3231 ( .A(p_input[9031]), .B(p_input[39031]), .Z(n2153) );
  AND U3232 ( .A(n2155), .B(n2156), .Z(o[9030]) );
  AND U3233 ( .A(p_input[29030]), .B(p_input[19030]), .Z(n2156) );
  AND U3234 ( .A(p_input[9030]), .B(p_input[39030]), .Z(n2155) );
  AND U3235 ( .A(n2157), .B(n2158), .Z(o[902]) );
  AND U3236 ( .A(p_input[20902]), .B(p_input[10902]), .Z(n2158) );
  AND U3237 ( .A(p_input[902]), .B(p_input[30902]), .Z(n2157) );
  AND U3238 ( .A(n2159), .B(n2160), .Z(o[9029]) );
  AND U3239 ( .A(p_input[29029]), .B(p_input[19029]), .Z(n2160) );
  AND U3240 ( .A(p_input[9029]), .B(p_input[39029]), .Z(n2159) );
  AND U3241 ( .A(n2161), .B(n2162), .Z(o[9028]) );
  AND U3242 ( .A(p_input[29028]), .B(p_input[19028]), .Z(n2162) );
  AND U3243 ( .A(p_input[9028]), .B(p_input[39028]), .Z(n2161) );
  AND U3244 ( .A(n2163), .B(n2164), .Z(o[9027]) );
  AND U3245 ( .A(p_input[29027]), .B(p_input[19027]), .Z(n2164) );
  AND U3246 ( .A(p_input[9027]), .B(p_input[39027]), .Z(n2163) );
  AND U3247 ( .A(n2165), .B(n2166), .Z(o[9026]) );
  AND U3248 ( .A(p_input[29026]), .B(p_input[19026]), .Z(n2166) );
  AND U3249 ( .A(p_input[9026]), .B(p_input[39026]), .Z(n2165) );
  AND U3250 ( .A(n2167), .B(n2168), .Z(o[9025]) );
  AND U3251 ( .A(p_input[29025]), .B(p_input[19025]), .Z(n2168) );
  AND U3252 ( .A(p_input[9025]), .B(p_input[39025]), .Z(n2167) );
  AND U3253 ( .A(n2169), .B(n2170), .Z(o[9024]) );
  AND U3254 ( .A(p_input[29024]), .B(p_input[19024]), .Z(n2170) );
  AND U3255 ( .A(p_input[9024]), .B(p_input[39024]), .Z(n2169) );
  AND U3256 ( .A(n2171), .B(n2172), .Z(o[9023]) );
  AND U3257 ( .A(p_input[29023]), .B(p_input[19023]), .Z(n2172) );
  AND U3258 ( .A(p_input[9023]), .B(p_input[39023]), .Z(n2171) );
  AND U3259 ( .A(n2173), .B(n2174), .Z(o[9022]) );
  AND U3260 ( .A(p_input[29022]), .B(p_input[19022]), .Z(n2174) );
  AND U3261 ( .A(p_input[9022]), .B(p_input[39022]), .Z(n2173) );
  AND U3262 ( .A(n2175), .B(n2176), .Z(o[9021]) );
  AND U3263 ( .A(p_input[29021]), .B(p_input[19021]), .Z(n2176) );
  AND U3264 ( .A(p_input[9021]), .B(p_input[39021]), .Z(n2175) );
  AND U3265 ( .A(n2177), .B(n2178), .Z(o[9020]) );
  AND U3266 ( .A(p_input[29020]), .B(p_input[19020]), .Z(n2178) );
  AND U3267 ( .A(p_input[9020]), .B(p_input[39020]), .Z(n2177) );
  AND U3268 ( .A(n2179), .B(n2180), .Z(o[901]) );
  AND U3269 ( .A(p_input[20901]), .B(p_input[10901]), .Z(n2180) );
  AND U3270 ( .A(p_input[901]), .B(p_input[30901]), .Z(n2179) );
  AND U3271 ( .A(n2181), .B(n2182), .Z(o[9019]) );
  AND U3272 ( .A(p_input[29019]), .B(p_input[19019]), .Z(n2182) );
  AND U3273 ( .A(p_input[9019]), .B(p_input[39019]), .Z(n2181) );
  AND U3274 ( .A(n2183), .B(n2184), .Z(o[9018]) );
  AND U3275 ( .A(p_input[29018]), .B(p_input[19018]), .Z(n2184) );
  AND U3276 ( .A(p_input[9018]), .B(p_input[39018]), .Z(n2183) );
  AND U3277 ( .A(n2185), .B(n2186), .Z(o[9017]) );
  AND U3278 ( .A(p_input[29017]), .B(p_input[19017]), .Z(n2186) );
  AND U3279 ( .A(p_input[9017]), .B(p_input[39017]), .Z(n2185) );
  AND U3280 ( .A(n2187), .B(n2188), .Z(o[9016]) );
  AND U3281 ( .A(p_input[29016]), .B(p_input[19016]), .Z(n2188) );
  AND U3282 ( .A(p_input[9016]), .B(p_input[39016]), .Z(n2187) );
  AND U3283 ( .A(n2189), .B(n2190), .Z(o[9015]) );
  AND U3284 ( .A(p_input[29015]), .B(p_input[19015]), .Z(n2190) );
  AND U3285 ( .A(p_input[9015]), .B(p_input[39015]), .Z(n2189) );
  AND U3286 ( .A(n2191), .B(n2192), .Z(o[9014]) );
  AND U3287 ( .A(p_input[29014]), .B(p_input[19014]), .Z(n2192) );
  AND U3288 ( .A(p_input[9014]), .B(p_input[39014]), .Z(n2191) );
  AND U3289 ( .A(n2193), .B(n2194), .Z(o[9013]) );
  AND U3290 ( .A(p_input[29013]), .B(p_input[19013]), .Z(n2194) );
  AND U3291 ( .A(p_input[9013]), .B(p_input[39013]), .Z(n2193) );
  AND U3292 ( .A(n2195), .B(n2196), .Z(o[9012]) );
  AND U3293 ( .A(p_input[29012]), .B(p_input[19012]), .Z(n2196) );
  AND U3294 ( .A(p_input[9012]), .B(p_input[39012]), .Z(n2195) );
  AND U3295 ( .A(n2197), .B(n2198), .Z(o[9011]) );
  AND U3296 ( .A(p_input[29011]), .B(p_input[19011]), .Z(n2198) );
  AND U3297 ( .A(p_input[9011]), .B(p_input[39011]), .Z(n2197) );
  AND U3298 ( .A(n2199), .B(n2200), .Z(o[9010]) );
  AND U3299 ( .A(p_input[29010]), .B(p_input[19010]), .Z(n2200) );
  AND U3300 ( .A(p_input[9010]), .B(p_input[39010]), .Z(n2199) );
  AND U3301 ( .A(n2201), .B(n2202), .Z(o[900]) );
  AND U3302 ( .A(p_input[20900]), .B(p_input[10900]), .Z(n2202) );
  AND U3303 ( .A(p_input[900]), .B(p_input[30900]), .Z(n2201) );
  AND U3304 ( .A(n2203), .B(n2204), .Z(o[9009]) );
  AND U3305 ( .A(p_input[29009]), .B(p_input[19009]), .Z(n2204) );
  AND U3306 ( .A(p_input[9009]), .B(p_input[39009]), .Z(n2203) );
  AND U3307 ( .A(n2205), .B(n2206), .Z(o[9008]) );
  AND U3308 ( .A(p_input[29008]), .B(p_input[19008]), .Z(n2206) );
  AND U3309 ( .A(p_input[9008]), .B(p_input[39008]), .Z(n2205) );
  AND U3310 ( .A(n2207), .B(n2208), .Z(o[9007]) );
  AND U3311 ( .A(p_input[29007]), .B(p_input[19007]), .Z(n2208) );
  AND U3312 ( .A(p_input[9007]), .B(p_input[39007]), .Z(n2207) );
  AND U3313 ( .A(n2209), .B(n2210), .Z(o[9006]) );
  AND U3314 ( .A(p_input[29006]), .B(p_input[19006]), .Z(n2210) );
  AND U3315 ( .A(p_input[9006]), .B(p_input[39006]), .Z(n2209) );
  AND U3316 ( .A(n2211), .B(n2212), .Z(o[9005]) );
  AND U3317 ( .A(p_input[29005]), .B(p_input[19005]), .Z(n2212) );
  AND U3318 ( .A(p_input[9005]), .B(p_input[39005]), .Z(n2211) );
  AND U3319 ( .A(n2213), .B(n2214), .Z(o[9004]) );
  AND U3320 ( .A(p_input[29004]), .B(p_input[19004]), .Z(n2214) );
  AND U3321 ( .A(p_input[9004]), .B(p_input[39004]), .Z(n2213) );
  AND U3322 ( .A(n2215), .B(n2216), .Z(o[9003]) );
  AND U3323 ( .A(p_input[29003]), .B(p_input[19003]), .Z(n2216) );
  AND U3324 ( .A(p_input[9003]), .B(p_input[39003]), .Z(n2215) );
  AND U3325 ( .A(n2217), .B(n2218), .Z(o[9002]) );
  AND U3326 ( .A(p_input[29002]), .B(p_input[19002]), .Z(n2218) );
  AND U3327 ( .A(p_input[9002]), .B(p_input[39002]), .Z(n2217) );
  AND U3328 ( .A(n2219), .B(n2220), .Z(o[9001]) );
  AND U3329 ( .A(p_input[29001]), .B(p_input[19001]), .Z(n2220) );
  AND U3330 ( .A(p_input[9001]), .B(p_input[39001]), .Z(n2219) );
  AND U3331 ( .A(n2221), .B(n2222), .Z(o[9000]) );
  AND U3332 ( .A(p_input[29000]), .B(p_input[19000]), .Z(n2222) );
  AND U3333 ( .A(p_input[9000]), .B(p_input[39000]), .Z(n2221) );
  AND U3334 ( .A(n2223), .B(n2224), .Z(o[8]) );
  AND U3335 ( .A(p_input[20008]), .B(p_input[10008]), .Z(n2224) );
  AND U3336 ( .A(p_input[8]), .B(p_input[30008]), .Z(n2223) );
  AND U3337 ( .A(n2225), .B(n2226), .Z(o[89]) );
  AND U3338 ( .A(p_input[20089]), .B(p_input[10089]), .Z(n2226) );
  AND U3339 ( .A(p_input[89]), .B(p_input[30089]), .Z(n2225) );
  AND U3340 ( .A(n2227), .B(n2228), .Z(o[899]) );
  AND U3341 ( .A(p_input[20899]), .B(p_input[10899]), .Z(n2228) );
  AND U3342 ( .A(p_input[899]), .B(p_input[30899]), .Z(n2227) );
  AND U3343 ( .A(n2229), .B(n2230), .Z(o[8999]) );
  AND U3344 ( .A(p_input[28999]), .B(p_input[18999]), .Z(n2230) );
  AND U3345 ( .A(p_input[8999]), .B(p_input[38999]), .Z(n2229) );
  AND U3346 ( .A(n2231), .B(n2232), .Z(o[8998]) );
  AND U3347 ( .A(p_input[28998]), .B(p_input[18998]), .Z(n2232) );
  AND U3348 ( .A(p_input[8998]), .B(p_input[38998]), .Z(n2231) );
  AND U3349 ( .A(n2233), .B(n2234), .Z(o[8997]) );
  AND U3350 ( .A(p_input[28997]), .B(p_input[18997]), .Z(n2234) );
  AND U3351 ( .A(p_input[8997]), .B(p_input[38997]), .Z(n2233) );
  AND U3352 ( .A(n2235), .B(n2236), .Z(o[8996]) );
  AND U3353 ( .A(p_input[28996]), .B(p_input[18996]), .Z(n2236) );
  AND U3354 ( .A(p_input[8996]), .B(p_input[38996]), .Z(n2235) );
  AND U3355 ( .A(n2237), .B(n2238), .Z(o[8995]) );
  AND U3356 ( .A(p_input[28995]), .B(p_input[18995]), .Z(n2238) );
  AND U3357 ( .A(p_input[8995]), .B(p_input[38995]), .Z(n2237) );
  AND U3358 ( .A(n2239), .B(n2240), .Z(o[8994]) );
  AND U3359 ( .A(p_input[28994]), .B(p_input[18994]), .Z(n2240) );
  AND U3360 ( .A(p_input[8994]), .B(p_input[38994]), .Z(n2239) );
  AND U3361 ( .A(n2241), .B(n2242), .Z(o[8993]) );
  AND U3362 ( .A(p_input[28993]), .B(p_input[18993]), .Z(n2242) );
  AND U3363 ( .A(p_input[8993]), .B(p_input[38993]), .Z(n2241) );
  AND U3364 ( .A(n2243), .B(n2244), .Z(o[8992]) );
  AND U3365 ( .A(p_input[28992]), .B(p_input[18992]), .Z(n2244) );
  AND U3366 ( .A(p_input[8992]), .B(p_input[38992]), .Z(n2243) );
  AND U3367 ( .A(n2245), .B(n2246), .Z(o[8991]) );
  AND U3368 ( .A(p_input[28991]), .B(p_input[18991]), .Z(n2246) );
  AND U3369 ( .A(p_input[8991]), .B(p_input[38991]), .Z(n2245) );
  AND U3370 ( .A(n2247), .B(n2248), .Z(o[8990]) );
  AND U3371 ( .A(p_input[28990]), .B(p_input[18990]), .Z(n2248) );
  AND U3372 ( .A(p_input[8990]), .B(p_input[38990]), .Z(n2247) );
  AND U3373 ( .A(n2249), .B(n2250), .Z(o[898]) );
  AND U3374 ( .A(p_input[20898]), .B(p_input[10898]), .Z(n2250) );
  AND U3375 ( .A(p_input[898]), .B(p_input[30898]), .Z(n2249) );
  AND U3376 ( .A(n2251), .B(n2252), .Z(o[8989]) );
  AND U3377 ( .A(p_input[28989]), .B(p_input[18989]), .Z(n2252) );
  AND U3378 ( .A(p_input[8989]), .B(p_input[38989]), .Z(n2251) );
  AND U3379 ( .A(n2253), .B(n2254), .Z(o[8988]) );
  AND U3380 ( .A(p_input[28988]), .B(p_input[18988]), .Z(n2254) );
  AND U3381 ( .A(p_input[8988]), .B(p_input[38988]), .Z(n2253) );
  AND U3382 ( .A(n2255), .B(n2256), .Z(o[8987]) );
  AND U3383 ( .A(p_input[28987]), .B(p_input[18987]), .Z(n2256) );
  AND U3384 ( .A(p_input[8987]), .B(p_input[38987]), .Z(n2255) );
  AND U3385 ( .A(n2257), .B(n2258), .Z(o[8986]) );
  AND U3386 ( .A(p_input[28986]), .B(p_input[18986]), .Z(n2258) );
  AND U3387 ( .A(p_input[8986]), .B(p_input[38986]), .Z(n2257) );
  AND U3388 ( .A(n2259), .B(n2260), .Z(o[8985]) );
  AND U3389 ( .A(p_input[28985]), .B(p_input[18985]), .Z(n2260) );
  AND U3390 ( .A(p_input[8985]), .B(p_input[38985]), .Z(n2259) );
  AND U3391 ( .A(n2261), .B(n2262), .Z(o[8984]) );
  AND U3392 ( .A(p_input[28984]), .B(p_input[18984]), .Z(n2262) );
  AND U3393 ( .A(p_input[8984]), .B(p_input[38984]), .Z(n2261) );
  AND U3394 ( .A(n2263), .B(n2264), .Z(o[8983]) );
  AND U3395 ( .A(p_input[28983]), .B(p_input[18983]), .Z(n2264) );
  AND U3396 ( .A(p_input[8983]), .B(p_input[38983]), .Z(n2263) );
  AND U3397 ( .A(n2265), .B(n2266), .Z(o[8982]) );
  AND U3398 ( .A(p_input[28982]), .B(p_input[18982]), .Z(n2266) );
  AND U3399 ( .A(p_input[8982]), .B(p_input[38982]), .Z(n2265) );
  AND U3400 ( .A(n2267), .B(n2268), .Z(o[8981]) );
  AND U3401 ( .A(p_input[28981]), .B(p_input[18981]), .Z(n2268) );
  AND U3402 ( .A(p_input[8981]), .B(p_input[38981]), .Z(n2267) );
  AND U3403 ( .A(n2269), .B(n2270), .Z(o[8980]) );
  AND U3404 ( .A(p_input[28980]), .B(p_input[18980]), .Z(n2270) );
  AND U3405 ( .A(p_input[8980]), .B(p_input[38980]), .Z(n2269) );
  AND U3406 ( .A(n2271), .B(n2272), .Z(o[897]) );
  AND U3407 ( .A(p_input[20897]), .B(p_input[10897]), .Z(n2272) );
  AND U3408 ( .A(p_input[897]), .B(p_input[30897]), .Z(n2271) );
  AND U3409 ( .A(n2273), .B(n2274), .Z(o[8979]) );
  AND U3410 ( .A(p_input[28979]), .B(p_input[18979]), .Z(n2274) );
  AND U3411 ( .A(p_input[8979]), .B(p_input[38979]), .Z(n2273) );
  AND U3412 ( .A(n2275), .B(n2276), .Z(o[8978]) );
  AND U3413 ( .A(p_input[28978]), .B(p_input[18978]), .Z(n2276) );
  AND U3414 ( .A(p_input[8978]), .B(p_input[38978]), .Z(n2275) );
  AND U3415 ( .A(n2277), .B(n2278), .Z(o[8977]) );
  AND U3416 ( .A(p_input[28977]), .B(p_input[18977]), .Z(n2278) );
  AND U3417 ( .A(p_input[8977]), .B(p_input[38977]), .Z(n2277) );
  AND U3418 ( .A(n2279), .B(n2280), .Z(o[8976]) );
  AND U3419 ( .A(p_input[28976]), .B(p_input[18976]), .Z(n2280) );
  AND U3420 ( .A(p_input[8976]), .B(p_input[38976]), .Z(n2279) );
  AND U3421 ( .A(n2281), .B(n2282), .Z(o[8975]) );
  AND U3422 ( .A(p_input[28975]), .B(p_input[18975]), .Z(n2282) );
  AND U3423 ( .A(p_input[8975]), .B(p_input[38975]), .Z(n2281) );
  AND U3424 ( .A(n2283), .B(n2284), .Z(o[8974]) );
  AND U3425 ( .A(p_input[28974]), .B(p_input[18974]), .Z(n2284) );
  AND U3426 ( .A(p_input[8974]), .B(p_input[38974]), .Z(n2283) );
  AND U3427 ( .A(n2285), .B(n2286), .Z(o[8973]) );
  AND U3428 ( .A(p_input[28973]), .B(p_input[18973]), .Z(n2286) );
  AND U3429 ( .A(p_input[8973]), .B(p_input[38973]), .Z(n2285) );
  AND U3430 ( .A(n2287), .B(n2288), .Z(o[8972]) );
  AND U3431 ( .A(p_input[28972]), .B(p_input[18972]), .Z(n2288) );
  AND U3432 ( .A(p_input[8972]), .B(p_input[38972]), .Z(n2287) );
  AND U3433 ( .A(n2289), .B(n2290), .Z(o[8971]) );
  AND U3434 ( .A(p_input[28971]), .B(p_input[18971]), .Z(n2290) );
  AND U3435 ( .A(p_input[8971]), .B(p_input[38971]), .Z(n2289) );
  AND U3436 ( .A(n2291), .B(n2292), .Z(o[8970]) );
  AND U3437 ( .A(p_input[28970]), .B(p_input[18970]), .Z(n2292) );
  AND U3438 ( .A(p_input[8970]), .B(p_input[38970]), .Z(n2291) );
  AND U3439 ( .A(n2293), .B(n2294), .Z(o[896]) );
  AND U3440 ( .A(p_input[20896]), .B(p_input[10896]), .Z(n2294) );
  AND U3441 ( .A(p_input[896]), .B(p_input[30896]), .Z(n2293) );
  AND U3442 ( .A(n2295), .B(n2296), .Z(o[8969]) );
  AND U3443 ( .A(p_input[28969]), .B(p_input[18969]), .Z(n2296) );
  AND U3444 ( .A(p_input[8969]), .B(p_input[38969]), .Z(n2295) );
  AND U3445 ( .A(n2297), .B(n2298), .Z(o[8968]) );
  AND U3446 ( .A(p_input[28968]), .B(p_input[18968]), .Z(n2298) );
  AND U3447 ( .A(p_input[8968]), .B(p_input[38968]), .Z(n2297) );
  AND U3448 ( .A(n2299), .B(n2300), .Z(o[8967]) );
  AND U3449 ( .A(p_input[28967]), .B(p_input[18967]), .Z(n2300) );
  AND U3450 ( .A(p_input[8967]), .B(p_input[38967]), .Z(n2299) );
  AND U3451 ( .A(n2301), .B(n2302), .Z(o[8966]) );
  AND U3452 ( .A(p_input[28966]), .B(p_input[18966]), .Z(n2302) );
  AND U3453 ( .A(p_input[8966]), .B(p_input[38966]), .Z(n2301) );
  AND U3454 ( .A(n2303), .B(n2304), .Z(o[8965]) );
  AND U3455 ( .A(p_input[28965]), .B(p_input[18965]), .Z(n2304) );
  AND U3456 ( .A(p_input[8965]), .B(p_input[38965]), .Z(n2303) );
  AND U3457 ( .A(n2305), .B(n2306), .Z(o[8964]) );
  AND U3458 ( .A(p_input[28964]), .B(p_input[18964]), .Z(n2306) );
  AND U3459 ( .A(p_input[8964]), .B(p_input[38964]), .Z(n2305) );
  AND U3460 ( .A(n2307), .B(n2308), .Z(o[8963]) );
  AND U3461 ( .A(p_input[28963]), .B(p_input[18963]), .Z(n2308) );
  AND U3462 ( .A(p_input[8963]), .B(p_input[38963]), .Z(n2307) );
  AND U3463 ( .A(n2309), .B(n2310), .Z(o[8962]) );
  AND U3464 ( .A(p_input[28962]), .B(p_input[18962]), .Z(n2310) );
  AND U3465 ( .A(p_input[8962]), .B(p_input[38962]), .Z(n2309) );
  AND U3466 ( .A(n2311), .B(n2312), .Z(o[8961]) );
  AND U3467 ( .A(p_input[28961]), .B(p_input[18961]), .Z(n2312) );
  AND U3468 ( .A(p_input[8961]), .B(p_input[38961]), .Z(n2311) );
  AND U3469 ( .A(n2313), .B(n2314), .Z(o[8960]) );
  AND U3470 ( .A(p_input[28960]), .B(p_input[18960]), .Z(n2314) );
  AND U3471 ( .A(p_input[8960]), .B(p_input[38960]), .Z(n2313) );
  AND U3472 ( .A(n2315), .B(n2316), .Z(o[895]) );
  AND U3473 ( .A(p_input[20895]), .B(p_input[10895]), .Z(n2316) );
  AND U3474 ( .A(p_input[895]), .B(p_input[30895]), .Z(n2315) );
  AND U3475 ( .A(n2317), .B(n2318), .Z(o[8959]) );
  AND U3476 ( .A(p_input[28959]), .B(p_input[18959]), .Z(n2318) );
  AND U3477 ( .A(p_input[8959]), .B(p_input[38959]), .Z(n2317) );
  AND U3478 ( .A(n2319), .B(n2320), .Z(o[8958]) );
  AND U3479 ( .A(p_input[28958]), .B(p_input[18958]), .Z(n2320) );
  AND U3480 ( .A(p_input[8958]), .B(p_input[38958]), .Z(n2319) );
  AND U3481 ( .A(n2321), .B(n2322), .Z(o[8957]) );
  AND U3482 ( .A(p_input[28957]), .B(p_input[18957]), .Z(n2322) );
  AND U3483 ( .A(p_input[8957]), .B(p_input[38957]), .Z(n2321) );
  AND U3484 ( .A(n2323), .B(n2324), .Z(o[8956]) );
  AND U3485 ( .A(p_input[28956]), .B(p_input[18956]), .Z(n2324) );
  AND U3486 ( .A(p_input[8956]), .B(p_input[38956]), .Z(n2323) );
  AND U3487 ( .A(n2325), .B(n2326), .Z(o[8955]) );
  AND U3488 ( .A(p_input[28955]), .B(p_input[18955]), .Z(n2326) );
  AND U3489 ( .A(p_input[8955]), .B(p_input[38955]), .Z(n2325) );
  AND U3490 ( .A(n2327), .B(n2328), .Z(o[8954]) );
  AND U3491 ( .A(p_input[28954]), .B(p_input[18954]), .Z(n2328) );
  AND U3492 ( .A(p_input[8954]), .B(p_input[38954]), .Z(n2327) );
  AND U3493 ( .A(n2329), .B(n2330), .Z(o[8953]) );
  AND U3494 ( .A(p_input[28953]), .B(p_input[18953]), .Z(n2330) );
  AND U3495 ( .A(p_input[8953]), .B(p_input[38953]), .Z(n2329) );
  AND U3496 ( .A(n2331), .B(n2332), .Z(o[8952]) );
  AND U3497 ( .A(p_input[28952]), .B(p_input[18952]), .Z(n2332) );
  AND U3498 ( .A(p_input[8952]), .B(p_input[38952]), .Z(n2331) );
  AND U3499 ( .A(n2333), .B(n2334), .Z(o[8951]) );
  AND U3500 ( .A(p_input[28951]), .B(p_input[18951]), .Z(n2334) );
  AND U3501 ( .A(p_input[8951]), .B(p_input[38951]), .Z(n2333) );
  AND U3502 ( .A(n2335), .B(n2336), .Z(o[8950]) );
  AND U3503 ( .A(p_input[28950]), .B(p_input[18950]), .Z(n2336) );
  AND U3504 ( .A(p_input[8950]), .B(p_input[38950]), .Z(n2335) );
  AND U3505 ( .A(n2337), .B(n2338), .Z(o[894]) );
  AND U3506 ( .A(p_input[20894]), .B(p_input[10894]), .Z(n2338) );
  AND U3507 ( .A(p_input[894]), .B(p_input[30894]), .Z(n2337) );
  AND U3508 ( .A(n2339), .B(n2340), .Z(o[8949]) );
  AND U3509 ( .A(p_input[28949]), .B(p_input[18949]), .Z(n2340) );
  AND U3510 ( .A(p_input[8949]), .B(p_input[38949]), .Z(n2339) );
  AND U3511 ( .A(n2341), .B(n2342), .Z(o[8948]) );
  AND U3512 ( .A(p_input[28948]), .B(p_input[18948]), .Z(n2342) );
  AND U3513 ( .A(p_input[8948]), .B(p_input[38948]), .Z(n2341) );
  AND U3514 ( .A(n2343), .B(n2344), .Z(o[8947]) );
  AND U3515 ( .A(p_input[28947]), .B(p_input[18947]), .Z(n2344) );
  AND U3516 ( .A(p_input[8947]), .B(p_input[38947]), .Z(n2343) );
  AND U3517 ( .A(n2345), .B(n2346), .Z(o[8946]) );
  AND U3518 ( .A(p_input[28946]), .B(p_input[18946]), .Z(n2346) );
  AND U3519 ( .A(p_input[8946]), .B(p_input[38946]), .Z(n2345) );
  AND U3520 ( .A(n2347), .B(n2348), .Z(o[8945]) );
  AND U3521 ( .A(p_input[28945]), .B(p_input[18945]), .Z(n2348) );
  AND U3522 ( .A(p_input[8945]), .B(p_input[38945]), .Z(n2347) );
  AND U3523 ( .A(n2349), .B(n2350), .Z(o[8944]) );
  AND U3524 ( .A(p_input[28944]), .B(p_input[18944]), .Z(n2350) );
  AND U3525 ( .A(p_input[8944]), .B(p_input[38944]), .Z(n2349) );
  AND U3526 ( .A(n2351), .B(n2352), .Z(o[8943]) );
  AND U3527 ( .A(p_input[28943]), .B(p_input[18943]), .Z(n2352) );
  AND U3528 ( .A(p_input[8943]), .B(p_input[38943]), .Z(n2351) );
  AND U3529 ( .A(n2353), .B(n2354), .Z(o[8942]) );
  AND U3530 ( .A(p_input[28942]), .B(p_input[18942]), .Z(n2354) );
  AND U3531 ( .A(p_input[8942]), .B(p_input[38942]), .Z(n2353) );
  AND U3532 ( .A(n2355), .B(n2356), .Z(o[8941]) );
  AND U3533 ( .A(p_input[28941]), .B(p_input[18941]), .Z(n2356) );
  AND U3534 ( .A(p_input[8941]), .B(p_input[38941]), .Z(n2355) );
  AND U3535 ( .A(n2357), .B(n2358), .Z(o[8940]) );
  AND U3536 ( .A(p_input[28940]), .B(p_input[18940]), .Z(n2358) );
  AND U3537 ( .A(p_input[8940]), .B(p_input[38940]), .Z(n2357) );
  AND U3538 ( .A(n2359), .B(n2360), .Z(o[893]) );
  AND U3539 ( .A(p_input[20893]), .B(p_input[10893]), .Z(n2360) );
  AND U3540 ( .A(p_input[893]), .B(p_input[30893]), .Z(n2359) );
  AND U3541 ( .A(n2361), .B(n2362), .Z(o[8939]) );
  AND U3542 ( .A(p_input[28939]), .B(p_input[18939]), .Z(n2362) );
  AND U3543 ( .A(p_input[8939]), .B(p_input[38939]), .Z(n2361) );
  AND U3544 ( .A(n2363), .B(n2364), .Z(o[8938]) );
  AND U3545 ( .A(p_input[28938]), .B(p_input[18938]), .Z(n2364) );
  AND U3546 ( .A(p_input[8938]), .B(p_input[38938]), .Z(n2363) );
  AND U3547 ( .A(n2365), .B(n2366), .Z(o[8937]) );
  AND U3548 ( .A(p_input[28937]), .B(p_input[18937]), .Z(n2366) );
  AND U3549 ( .A(p_input[8937]), .B(p_input[38937]), .Z(n2365) );
  AND U3550 ( .A(n2367), .B(n2368), .Z(o[8936]) );
  AND U3551 ( .A(p_input[28936]), .B(p_input[18936]), .Z(n2368) );
  AND U3552 ( .A(p_input[8936]), .B(p_input[38936]), .Z(n2367) );
  AND U3553 ( .A(n2369), .B(n2370), .Z(o[8935]) );
  AND U3554 ( .A(p_input[28935]), .B(p_input[18935]), .Z(n2370) );
  AND U3555 ( .A(p_input[8935]), .B(p_input[38935]), .Z(n2369) );
  AND U3556 ( .A(n2371), .B(n2372), .Z(o[8934]) );
  AND U3557 ( .A(p_input[28934]), .B(p_input[18934]), .Z(n2372) );
  AND U3558 ( .A(p_input[8934]), .B(p_input[38934]), .Z(n2371) );
  AND U3559 ( .A(n2373), .B(n2374), .Z(o[8933]) );
  AND U3560 ( .A(p_input[28933]), .B(p_input[18933]), .Z(n2374) );
  AND U3561 ( .A(p_input[8933]), .B(p_input[38933]), .Z(n2373) );
  AND U3562 ( .A(n2375), .B(n2376), .Z(o[8932]) );
  AND U3563 ( .A(p_input[28932]), .B(p_input[18932]), .Z(n2376) );
  AND U3564 ( .A(p_input[8932]), .B(p_input[38932]), .Z(n2375) );
  AND U3565 ( .A(n2377), .B(n2378), .Z(o[8931]) );
  AND U3566 ( .A(p_input[28931]), .B(p_input[18931]), .Z(n2378) );
  AND U3567 ( .A(p_input[8931]), .B(p_input[38931]), .Z(n2377) );
  AND U3568 ( .A(n2379), .B(n2380), .Z(o[8930]) );
  AND U3569 ( .A(p_input[28930]), .B(p_input[18930]), .Z(n2380) );
  AND U3570 ( .A(p_input[8930]), .B(p_input[38930]), .Z(n2379) );
  AND U3571 ( .A(n2381), .B(n2382), .Z(o[892]) );
  AND U3572 ( .A(p_input[20892]), .B(p_input[10892]), .Z(n2382) );
  AND U3573 ( .A(p_input[892]), .B(p_input[30892]), .Z(n2381) );
  AND U3574 ( .A(n2383), .B(n2384), .Z(o[8929]) );
  AND U3575 ( .A(p_input[28929]), .B(p_input[18929]), .Z(n2384) );
  AND U3576 ( .A(p_input[8929]), .B(p_input[38929]), .Z(n2383) );
  AND U3577 ( .A(n2385), .B(n2386), .Z(o[8928]) );
  AND U3578 ( .A(p_input[28928]), .B(p_input[18928]), .Z(n2386) );
  AND U3579 ( .A(p_input[8928]), .B(p_input[38928]), .Z(n2385) );
  AND U3580 ( .A(n2387), .B(n2388), .Z(o[8927]) );
  AND U3581 ( .A(p_input[28927]), .B(p_input[18927]), .Z(n2388) );
  AND U3582 ( .A(p_input[8927]), .B(p_input[38927]), .Z(n2387) );
  AND U3583 ( .A(n2389), .B(n2390), .Z(o[8926]) );
  AND U3584 ( .A(p_input[28926]), .B(p_input[18926]), .Z(n2390) );
  AND U3585 ( .A(p_input[8926]), .B(p_input[38926]), .Z(n2389) );
  AND U3586 ( .A(n2391), .B(n2392), .Z(o[8925]) );
  AND U3587 ( .A(p_input[28925]), .B(p_input[18925]), .Z(n2392) );
  AND U3588 ( .A(p_input[8925]), .B(p_input[38925]), .Z(n2391) );
  AND U3589 ( .A(n2393), .B(n2394), .Z(o[8924]) );
  AND U3590 ( .A(p_input[28924]), .B(p_input[18924]), .Z(n2394) );
  AND U3591 ( .A(p_input[8924]), .B(p_input[38924]), .Z(n2393) );
  AND U3592 ( .A(n2395), .B(n2396), .Z(o[8923]) );
  AND U3593 ( .A(p_input[28923]), .B(p_input[18923]), .Z(n2396) );
  AND U3594 ( .A(p_input[8923]), .B(p_input[38923]), .Z(n2395) );
  AND U3595 ( .A(n2397), .B(n2398), .Z(o[8922]) );
  AND U3596 ( .A(p_input[28922]), .B(p_input[18922]), .Z(n2398) );
  AND U3597 ( .A(p_input[8922]), .B(p_input[38922]), .Z(n2397) );
  AND U3598 ( .A(n2399), .B(n2400), .Z(o[8921]) );
  AND U3599 ( .A(p_input[28921]), .B(p_input[18921]), .Z(n2400) );
  AND U3600 ( .A(p_input[8921]), .B(p_input[38921]), .Z(n2399) );
  AND U3601 ( .A(n2401), .B(n2402), .Z(o[8920]) );
  AND U3602 ( .A(p_input[28920]), .B(p_input[18920]), .Z(n2402) );
  AND U3603 ( .A(p_input[8920]), .B(p_input[38920]), .Z(n2401) );
  AND U3604 ( .A(n2403), .B(n2404), .Z(o[891]) );
  AND U3605 ( .A(p_input[20891]), .B(p_input[10891]), .Z(n2404) );
  AND U3606 ( .A(p_input[891]), .B(p_input[30891]), .Z(n2403) );
  AND U3607 ( .A(n2405), .B(n2406), .Z(o[8919]) );
  AND U3608 ( .A(p_input[28919]), .B(p_input[18919]), .Z(n2406) );
  AND U3609 ( .A(p_input[8919]), .B(p_input[38919]), .Z(n2405) );
  AND U3610 ( .A(n2407), .B(n2408), .Z(o[8918]) );
  AND U3611 ( .A(p_input[28918]), .B(p_input[18918]), .Z(n2408) );
  AND U3612 ( .A(p_input[8918]), .B(p_input[38918]), .Z(n2407) );
  AND U3613 ( .A(n2409), .B(n2410), .Z(o[8917]) );
  AND U3614 ( .A(p_input[28917]), .B(p_input[18917]), .Z(n2410) );
  AND U3615 ( .A(p_input[8917]), .B(p_input[38917]), .Z(n2409) );
  AND U3616 ( .A(n2411), .B(n2412), .Z(o[8916]) );
  AND U3617 ( .A(p_input[28916]), .B(p_input[18916]), .Z(n2412) );
  AND U3618 ( .A(p_input[8916]), .B(p_input[38916]), .Z(n2411) );
  AND U3619 ( .A(n2413), .B(n2414), .Z(o[8915]) );
  AND U3620 ( .A(p_input[28915]), .B(p_input[18915]), .Z(n2414) );
  AND U3621 ( .A(p_input[8915]), .B(p_input[38915]), .Z(n2413) );
  AND U3622 ( .A(n2415), .B(n2416), .Z(o[8914]) );
  AND U3623 ( .A(p_input[28914]), .B(p_input[18914]), .Z(n2416) );
  AND U3624 ( .A(p_input[8914]), .B(p_input[38914]), .Z(n2415) );
  AND U3625 ( .A(n2417), .B(n2418), .Z(o[8913]) );
  AND U3626 ( .A(p_input[28913]), .B(p_input[18913]), .Z(n2418) );
  AND U3627 ( .A(p_input[8913]), .B(p_input[38913]), .Z(n2417) );
  AND U3628 ( .A(n2419), .B(n2420), .Z(o[8912]) );
  AND U3629 ( .A(p_input[28912]), .B(p_input[18912]), .Z(n2420) );
  AND U3630 ( .A(p_input[8912]), .B(p_input[38912]), .Z(n2419) );
  AND U3631 ( .A(n2421), .B(n2422), .Z(o[8911]) );
  AND U3632 ( .A(p_input[28911]), .B(p_input[18911]), .Z(n2422) );
  AND U3633 ( .A(p_input[8911]), .B(p_input[38911]), .Z(n2421) );
  AND U3634 ( .A(n2423), .B(n2424), .Z(o[8910]) );
  AND U3635 ( .A(p_input[28910]), .B(p_input[18910]), .Z(n2424) );
  AND U3636 ( .A(p_input[8910]), .B(p_input[38910]), .Z(n2423) );
  AND U3637 ( .A(n2425), .B(n2426), .Z(o[890]) );
  AND U3638 ( .A(p_input[20890]), .B(p_input[10890]), .Z(n2426) );
  AND U3639 ( .A(p_input[890]), .B(p_input[30890]), .Z(n2425) );
  AND U3640 ( .A(n2427), .B(n2428), .Z(o[8909]) );
  AND U3641 ( .A(p_input[28909]), .B(p_input[18909]), .Z(n2428) );
  AND U3642 ( .A(p_input[8909]), .B(p_input[38909]), .Z(n2427) );
  AND U3643 ( .A(n2429), .B(n2430), .Z(o[8908]) );
  AND U3644 ( .A(p_input[28908]), .B(p_input[18908]), .Z(n2430) );
  AND U3645 ( .A(p_input[8908]), .B(p_input[38908]), .Z(n2429) );
  AND U3646 ( .A(n2431), .B(n2432), .Z(o[8907]) );
  AND U3647 ( .A(p_input[28907]), .B(p_input[18907]), .Z(n2432) );
  AND U3648 ( .A(p_input[8907]), .B(p_input[38907]), .Z(n2431) );
  AND U3649 ( .A(n2433), .B(n2434), .Z(o[8906]) );
  AND U3650 ( .A(p_input[28906]), .B(p_input[18906]), .Z(n2434) );
  AND U3651 ( .A(p_input[8906]), .B(p_input[38906]), .Z(n2433) );
  AND U3652 ( .A(n2435), .B(n2436), .Z(o[8905]) );
  AND U3653 ( .A(p_input[28905]), .B(p_input[18905]), .Z(n2436) );
  AND U3654 ( .A(p_input[8905]), .B(p_input[38905]), .Z(n2435) );
  AND U3655 ( .A(n2437), .B(n2438), .Z(o[8904]) );
  AND U3656 ( .A(p_input[28904]), .B(p_input[18904]), .Z(n2438) );
  AND U3657 ( .A(p_input[8904]), .B(p_input[38904]), .Z(n2437) );
  AND U3658 ( .A(n2439), .B(n2440), .Z(o[8903]) );
  AND U3659 ( .A(p_input[28903]), .B(p_input[18903]), .Z(n2440) );
  AND U3660 ( .A(p_input[8903]), .B(p_input[38903]), .Z(n2439) );
  AND U3661 ( .A(n2441), .B(n2442), .Z(o[8902]) );
  AND U3662 ( .A(p_input[28902]), .B(p_input[18902]), .Z(n2442) );
  AND U3663 ( .A(p_input[8902]), .B(p_input[38902]), .Z(n2441) );
  AND U3664 ( .A(n2443), .B(n2444), .Z(o[8901]) );
  AND U3665 ( .A(p_input[28901]), .B(p_input[18901]), .Z(n2444) );
  AND U3666 ( .A(p_input[8901]), .B(p_input[38901]), .Z(n2443) );
  AND U3667 ( .A(n2445), .B(n2446), .Z(o[8900]) );
  AND U3668 ( .A(p_input[28900]), .B(p_input[18900]), .Z(n2446) );
  AND U3669 ( .A(p_input[8900]), .B(p_input[38900]), .Z(n2445) );
  AND U3670 ( .A(n2447), .B(n2448), .Z(o[88]) );
  AND U3671 ( .A(p_input[20088]), .B(p_input[10088]), .Z(n2448) );
  AND U3672 ( .A(p_input[88]), .B(p_input[30088]), .Z(n2447) );
  AND U3673 ( .A(n2449), .B(n2450), .Z(o[889]) );
  AND U3674 ( .A(p_input[20889]), .B(p_input[10889]), .Z(n2450) );
  AND U3675 ( .A(p_input[889]), .B(p_input[30889]), .Z(n2449) );
  AND U3676 ( .A(n2451), .B(n2452), .Z(o[8899]) );
  AND U3677 ( .A(p_input[28899]), .B(p_input[18899]), .Z(n2452) );
  AND U3678 ( .A(p_input[8899]), .B(p_input[38899]), .Z(n2451) );
  AND U3679 ( .A(n2453), .B(n2454), .Z(o[8898]) );
  AND U3680 ( .A(p_input[28898]), .B(p_input[18898]), .Z(n2454) );
  AND U3681 ( .A(p_input[8898]), .B(p_input[38898]), .Z(n2453) );
  AND U3682 ( .A(n2455), .B(n2456), .Z(o[8897]) );
  AND U3683 ( .A(p_input[28897]), .B(p_input[18897]), .Z(n2456) );
  AND U3684 ( .A(p_input[8897]), .B(p_input[38897]), .Z(n2455) );
  AND U3685 ( .A(n2457), .B(n2458), .Z(o[8896]) );
  AND U3686 ( .A(p_input[28896]), .B(p_input[18896]), .Z(n2458) );
  AND U3687 ( .A(p_input[8896]), .B(p_input[38896]), .Z(n2457) );
  AND U3688 ( .A(n2459), .B(n2460), .Z(o[8895]) );
  AND U3689 ( .A(p_input[28895]), .B(p_input[18895]), .Z(n2460) );
  AND U3690 ( .A(p_input[8895]), .B(p_input[38895]), .Z(n2459) );
  AND U3691 ( .A(n2461), .B(n2462), .Z(o[8894]) );
  AND U3692 ( .A(p_input[28894]), .B(p_input[18894]), .Z(n2462) );
  AND U3693 ( .A(p_input[8894]), .B(p_input[38894]), .Z(n2461) );
  AND U3694 ( .A(n2463), .B(n2464), .Z(o[8893]) );
  AND U3695 ( .A(p_input[28893]), .B(p_input[18893]), .Z(n2464) );
  AND U3696 ( .A(p_input[8893]), .B(p_input[38893]), .Z(n2463) );
  AND U3697 ( .A(n2465), .B(n2466), .Z(o[8892]) );
  AND U3698 ( .A(p_input[28892]), .B(p_input[18892]), .Z(n2466) );
  AND U3699 ( .A(p_input[8892]), .B(p_input[38892]), .Z(n2465) );
  AND U3700 ( .A(n2467), .B(n2468), .Z(o[8891]) );
  AND U3701 ( .A(p_input[28891]), .B(p_input[18891]), .Z(n2468) );
  AND U3702 ( .A(p_input[8891]), .B(p_input[38891]), .Z(n2467) );
  AND U3703 ( .A(n2469), .B(n2470), .Z(o[8890]) );
  AND U3704 ( .A(p_input[28890]), .B(p_input[18890]), .Z(n2470) );
  AND U3705 ( .A(p_input[8890]), .B(p_input[38890]), .Z(n2469) );
  AND U3706 ( .A(n2471), .B(n2472), .Z(o[888]) );
  AND U3707 ( .A(p_input[20888]), .B(p_input[10888]), .Z(n2472) );
  AND U3708 ( .A(p_input[888]), .B(p_input[30888]), .Z(n2471) );
  AND U3709 ( .A(n2473), .B(n2474), .Z(o[8889]) );
  AND U3710 ( .A(p_input[28889]), .B(p_input[18889]), .Z(n2474) );
  AND U3711 ( .A(p_input[8889]), .B(p_input[38889]), .Z(n2473) );
  AND U3712 ( .A(n2475), .B(n2476), .Z(o[8888]) );
  AND U3713 ( .A(p_input[28888]), .B(p_input[18888]), .Z(n2476) );
  AND U3714 ( .A(p_input[8888]), .B(p_input[38888]), .Z(n2475) );
  AND U3715 ( .A(n2477), .B(n2478), .Z(o[8887]) );
  AND U3716 ( .A(p_input[28887]), .B(p_input[18887]), .Z(n2478) );
  AND U3717 ( .A(p_input[8887]), .B(p_input[38887]), .Z(n2477) );
  AND U3718 ( .A(n2479), .B(n2480), .Z(o[8886]) );
  AND U3719 ( .A(p_input[28886]), .B(p_input[18886]), .Z(n2480) );
  AND U3720 ( .A(p_input[8886]), .B(p_input[38886]), .Z(n2479) );
  AND U3721 ( .A(n2481), .B(n2482), .Z(o[8885]) );
  AND U3722 ( .A(p_input[28885]), .B(p_input[18885]), .Z(n2482) );
  AND U3723 ( .A(p_input[8885]), .B(p_input[38885]), .Z(n2481) );
  AND U3724 ( .A(n2483), .B(n2484), .Z(o[8884]) );
  AND U3725 ( .A(p_input[28884]), .B(p_input[18884]), .Z(n2484) );
  AND U3726 ( .A(p_input[8884]), .B(p_input[38884]), .Z(n2483) );
  AND U3727 ( .A(n2485), .B(n2486), .Z(o[8883]) );
  AND U3728 ( .A(p_input[28883]), .B(p_input[18883]), .Z(n2486) );
  AND U3729 ( .A(p_input[8883]), .B(p_input[38883]), .Z(n2485) );
  AND U3730 ( .A(n2487), .B(n2488), .Z(o[8882]) );
  AND U3731 ( .A(p_input[28882]), .B(p_input[18882]), .Z(n2488) );
  AND U3732 ( .A(p_input[8882]), .B(p_input[38882]), .Z(n2487) );
  AND U3733 ( .A(n2489), .B(n2490), .Z(o[8881]) );
  AND U3734 ( .A(p_input[28881]), .B(p_input[18881]), .Z(n2490) );
  AND U3735 ( .A(p_input[8881]), .B(p_input[38881]), .Z(n2489) );
  AND U3736 ( .A(n2491), .B(n2492), .Z(o[8880]) );
  AND U3737 ( .A(p_input[28880]), .B(p_input[18880]), .Z(n2492) );
  AND U3738 ( .A(p_input[8880]), .B(p_input[38880]), .Z(n2491) );
  AND U3739 ( .A(n2493), .B(n2494), .Z(o[887]) );
  AND U3740 ( .A(p_input[20887]), .B(p_input[10887]), .Z(n2494) );
  AND U3741 ( .A(p_input[887]), .B(p_input[30887]), .Z(n2493) );
  AND U3742 ( .A(n2495), .B(n2496), .Z(o[8879]) );
  AND U3743 ( .A(p_input[28879]), .B(p_input[18879]), .Z(n2496) );
  AND U3744 ( .A(p_input[8879]), .B(p_input[38879]), .Z(n2495) );
  AND U3745 ( .A(n2497), .B(n2498), .Z(o[8878]) );
  AND U3746 ( .A(p_input[28878]), .B(p_input[18878]), .Z(n2498) );
  AND U3747 ( .A(p_input[8878]), .B(p_input[38878]), .Z(n2497) );
  AND U3748 ( .A(n2499), .B(n2500), .Z(o[8877]) );
  AND U3749 ( .A(p_input[28877]), .B(p_input[18877]), .Z(n2500) );
  AND U3750 ( .A(p_input[8877]), .B(p_input[38877]), .Z(n2499) );
  AND U3751 ( .A(n2501), .B(n2502), .Z(o[8876]) );
  AND U3752 ( .A(p_input[28876]), .B(p_input[18876]), .Z(n2502) );
  AND U3753 ( .A(p_input[8876]), .B(p_input[38876]), .Z(n2501) );
  AND U3754 ( .A(n2503), .B(n2504), .Z(o[8875]) );
  AND U3755 ( .A(p_input[28875]), .B(p_input[18875]), .Z(n2504) );
  AND U3756 ( .A(p_input[8875]), .B(p_input[38875]), .Z(n2503) );
  AND U3757 ( .A(n2505), .B(n2506), .Z(o[8874]) );
  AND U3758 ( .A(p_input[28874]), .B(p_input[18874]), .Z(n2506) );
  AND U3759 ( .A(p_input[8874]), .B(p_input[38874]), .Z(n2505) );
  AND U3760 ( .A(n2507), .B(n2508), .Z(o[8873]) );
  AND U3761 ( .A(p_input[28873]), .B(p_input[18873]), .Z(n2508) );
  AND U3762 ( .A(p_input[8873]), .B(p_input[38873]), .Z(n2507) );
  AND U3763 ( .A(n2509), .B(n2510), .Z(o[8872]) );
  AND U3764 ( .A(p_input[28872]), .B(p_input[18872]), .Z(n2510) );
  AND U3765 ( .A(p_input[8872]), .B(p_input[38872]), .Z(n2509) );
  AND U3766 ( .A(n2511), .B(n2512), .Z(o[8871]) );
  AND U3767 ( .A(p_input[28871]), .B(p_input[18871]), .Z(n2512) );
  AND U3768 ( .A(p_input[8871]), .B(p_input[38871]), .Z(n2511) );
  AND U3769 ( .A(n2513), .B(n2514), .Z(o[8870]) );
  AND U3770 ( .A(p_input[28870]), .B(p_input[18870]), .Z(n2514) );
  AND U3771 ( .A(p_input[8870]), .B(p_input[38870]), .Z(n2513) );
  AND U3772 ( .A(n2515), .B(n2516), .Z(o[886]) );
  AND U3773 ( .A(p_input[20886]), .B(p_input[10886]), .Z(n2516) );
  AND U3774 ( .A(p_input[886]), .B(p_input[30886]), .Z(n2515) );
  AND U3775 ( .A(n2517), .B(n2518), .Z(o[8869]) );
  AND U3776 ( .A(p_input[28869]), .B(p_input[18869]), .Z(n2518) );
  AND U3777 ( .A(p_input[8869]), .B(p_input[38869]), .Z(n2517) );
  AND U3778 ( .A(n2519), .B(n2520), .Z(o[8868]) );
  AND U3779 ( .A(p_input[28868]), .B(p_input[18868]), .Z(n2520) );
  AND U3780 ( .A(p_input[8868]), .B(p_input[38868]), .Z(n2519) );
  AND U3781 ( .A(n2521), .B(n2522), .Z(o[8867]) );
  AND U3782 ( .A(p_input[28867]), .B(p_input[18867]), .Z(n2522) );
  AND U3783 ( .A(p_input[8867]), .B(p_input[38867]), .Z(n2521) );
  AND U3784 ( .A(n2523), .B(n2524), .Z(o[8866]) );
  AND U3785 ( .A(p_input[28866]), .B(p_input[18866]), .Z(n2524) );
  AND U3786 ( .A(p_input[8866]), .B(p_input[38866]), .Z(n2523) );
  AND U3787 ( .A(n2525), .B(n2526), .Z(o[8865]) );
  AND U3788 ( .A(p_input[28865]), .B(p_input[18865]), .Z(n2526) );
  AND U3789 ( .A(p_input[8865]), .B(p_input[38865]), .Z(n2525) );
  AND U3790 ( .A(n2527), .B(n2528), .Z(o[8864]) );
  AND U3791 ( .A(p_input[28864]), .B(p_input[18864]), .Z(n2528) );
  AND U3792 ( .A(p_input[8864]), .B(p_input[38864]), .Z(n2527) );
  AND U3793 ( .A(n2529), .B(n2530), .Z(o[8863]) );
  AND U3794 ( .A(p_input[28863]), .B(p_input[18863]), .Z(n2530) );
  AND U3795 ( .A(p_input[8863]), .B(p_input[38863]), .Z(n2529) );
  AND U3796 ( .A(n2531), .B(n2532), .Z(o[8862]) );
  AND U3797 ( .A(p_input[28862]), .B(p_input[18862]), .Z(n2532) );
  AND U3798 ( .A(p_input[8862]), .B(p_input[38862]), .Z(n2531) );
  AND U3799 ( .A(n2533), .B(n2534), .Z(o[8861]) );
  AND U3800 ( .A(p_input[28861]), .B(p_input[18861]), .Z(n2534) );
  AND U3801 ( .A(p_input[8861]), .B(p_input[38861]), .Z(n2533) );
  AND U3802 ( .A(n2535), .B(n2536), .Z(o[8860]) );
  AND U3803 ( .A(p_input[28860]), .B(p_input[18860]), .Z(n2536) );
  AND U3804 ( .A(p_input[8860]), .B(p_input[38860]), .Z(n2535) );
  AND U3805 ( .A(n2537), .B(n2538), .Z(o[885]) );
  AND U3806 ( .A(p_input[20885]), .B(p_input[10885]), .Z(n2538) );
  AND U3807 ( .A(p_input[885]), .B(p_input[30885]), .Z(n2537) );
  AND U3808 ( .A(n2539), .B(n2540), .Z(o[8859]) );
  AND U3809 ( .A(p_input[28859]), .B(p_input[18859]), .Z(n2540) );
  AND U3810 ( .A(p_input[8859]), .B(p_input[38859]), .Z(n2539) );
  AND U3811 ( .A(n2541), .B(n2542), .Z(o[8858]) );
  AND U3812 ( .A(p_input[28858]), .B(p_input[18858]), .Z(n2542) );
  AND U3813 ( .A(p_input[8858]), .B(p_input[38858]), .Z(n2541) );
  AND U3814 ( .A(n2543), .B(n2544), .Z(o[8857]) );
  AND U3815 ( .A(p_input[28857]), .B(p_input[18857]), .Z(n2544) );
  AND U3816 ( .A(p_input[8857]), .B(p_input[38857]), .Z(n2543) );
  AND U3817 ( .A(n2545), .B(n2546), .Z(o[8856]) );
  AND U3818 ( .A(p_input[28856]), .B(p_input[18856]), .Z(n2546) );
  AND U3819 ( .A(p_input[8856]), .B(p_input[38856]), .Z(n2545) );
  AND U3820 ( .A(n2547), .B(n2548), .Z(o[8855]) );
  AND U3821 ( .A(p_input[28855]), .B(p_input[18855]), .Z(n2548) );
  AND U3822 ( .A(p_input[8855]), .B(p_input[38855]), .Z(n2547) );
  AND U3823 ( .A(n2549), .B(n2550), .Z(o[8854]) );
  AND U3824 ( .A(p_input[28854]), .B(p_input[18854]), .Z(n2550) );
  AND U3825 ( .A(p_input[8854]), .B(p_input[38854]), .Z(n2549) );
  AND U3826 ( .A(n2551), .B(n2552), .Z(o[8853]) );
  AND U3827 ( .A(p_input[28853]), .B(p_input[18853]), .Z(n2552) );
  AND U3828 ( .A(p_input[8853]), .B(p_input[38853]), .Z(n2551) );
  AND U3829 ( .A(n2553), .B(n2554), .Z(o[8852]) );
  AND U3830 ( .A(p_input[28852]), .B(p_input[18852]), .Z(n2554) );
  AND U3831 ( .A(p_input[8852]), .B(p_input[38852]), .Z(n2553) );
  AND U3832 ( .A(n2555), .B(n2556), .Z(o[8851]) );
  AND U3833 ( .A(p_input[28851]), .B(p_input[18851]), .Z(n2556) );
  AND U3834 ( .A(p_input[8851]), .B(p_input[38851]), .Z(n2555) );
  AND U3835 ( .A(n2557), .B(n2558), .Z(o[8850]) );
  AND U3836 ( .A(p_input[28850]), .B(p_input[18850]), .Z(n2558) );
  AND U3837 ( .A(p_input[8850]), .B(p_input[38850]), .Z(n2557) );
  AND U3838 ( .A(n2559), .B(n2560), .Z(o[884]) );
  AND U3839 ( .A(p_input[20884]), .B(p_input[10884]), .Z(n2560) );
  AND U3840 ( .A(p_input[884]), .B(p_input[30884]), .Z(n2559) );
  AND U3841 ( .A(n2561), .B(n2562), .Z(o[8849]) );
  AND U3842 ( .A(p_input[28849]), .B(p_input[18849]), .Z(n2562) );
  AND U3843 ( .A(p_input[8849]), .B(p_input[38849]), .Z(n2561) );
  AND U3844 ( .A(n2563), .B(n2564), .Z(o[8848]) );
  AND U3845 ( .A(p_input[28848]), .B(p_input[18848]), .Z(n2564) );
  AND U3846 ( .A(p_input[8848]), .B(p_input[38848]), .Z(n2563) );
  AND U3847 ( .A(n2565), .B(n2566), .Z(o[8847]) );
  AND U3848 ( .A(p_input[28847]), .B(p_input[18847]), .Z(n2566) );
  AND U3849 ( .A(p_input[8847]), .B(p_input[38847]), .Z(n2565) );
  AND U3850 ( .A(n2567), .B(n2568), .Z(o[8846]) );
  AND U3851 ( .A(p_input[28846]), .B(p_input[18846]), .Z(n2568) );
  AND U3852 ( .A(p_input[8846]), .B(p_input[38846]), .Z(n2567) );
  AND U3853 ( .A(n2569), .B(n2570), .Z(o[8845]) );
  AND U3854 ( .A(p_input[28845]), .B(p_input[18845]), .Z(n2570) );
  AND U3855 ( .A(p_input[8845]), .B(p_input[38845]), .Z(n2569) );
  AND U3856 ( .A(n2571), .B(n2572), .Z(o[8844]) );
  AND U3857 ( .A(p_input[28844]), .B(p_input[18844]), .Z(n2572) );
  AND U3858 ( .A(p_input[8844]), .B(p_input[38844]), .Z(n2571) );
  AND U3859 ( .A(n2573), .B(n2574), .Z(o[8843]) );
  AND U3860 ( .A(p_input[28843]), .B(p_input[18843]), .Z(n2574) );
  AND U3861 ( .A(p_input[8843]), .B(p_input[38843]), .Z(n2573) );
  AND U3862 ( .A(n2575), .B(n2576), .Z(o[8842]) );
  AND U3863 ( .A(p_input[28842]), .B(p_input[18842]), .Z(n2576) );
  AND U3864 ( .A(p_input[8842]), .B(p_input[38842]), .Z(n2575) );
  AND U3865 ( .A(n2577), .B(n2578), .Z(o[8841]) );
  AND U3866 ( .A(p_input[28841]), .B(p_input[18841]), .Z(n2578) );
  AND U3867 ( .A(p_input[8841]), .B(p_input[38841]), .Z(n2577) );
  AND U3868 ( .A(n2579), .B(n2580), .Z(o[8840]) );
  AND U3869 ( .A(p_input[28840]), .B(p_input[18840]), .Z(n2580) );
  AND U3870 ( .A(p_input[8840]), .B(p_input[38840]), .Z(n2579) );
  AND U3871 ( .A(n2581), .B(n2582), .Z(o[883]) );
  AND U3872 ( .A(p_input[20883]), .B(p_input[10883]), .Z(n2582) );
  AND U3873 ( .A(p_input[883]), .B(p_input[30883]), .Z(n2581) );
  AND U3874 ( .A(n2583), .B(n2584), .Z(o[8839]) );
  AND U3875 ( .A(p_input[28839]), .B(p_input[18839]), .Z(n2584) );
  AND U3876 ( .A(p_input[8839]), .B(p_input[38839]), .Z(n2583) );
  AND U3877 ( .A(n2585), .B(n2586), .Z(o[8838]) );
  AND U3878 ( .A(p_input[28838]), .B(p_input[18838]), .Z(n2586) );
  AND U3879 ( .A(p_input[8838]), .B(p_input[38838]), .Z(n2585) );
  AND U3880 ( .A(n2587), .B(n2588), .Z(o[8837]) );
  AND U3881 ( .A(p_input[28837]), .B(p_input[18837]), .Z(n2588) );
  AND U3882 ( .A(p_input[8837]), .B(p_input[38837]), .Z(n2587) );
  AND U3883 ( .A(n2589), .B(n2590), .Z(o[8836]) );
  AND U3884 ( .A(p_input[28836]), .B(p_input[18836]), .Z(n2590) );
  AND U3885 ( .A(p_input[8836]), .B(p_input[38836]), .Z(n2589) );
  AND U3886 ( .A(n2591), .B(n2592), .Z(o[8835]) );
  AND U3887 ( .A(p_input[28835]), .B(p_input[18835]), .Z(n2592) );
  AND U3888 ( .A(p_input[8835]), .B(p_input[38835]), .Z(n2591) );
  AND U3889 ( .A(n2593), .B(n2594), .Z(o[8834]) );
  AND U3890 ( .A(p_input[28834]), .B(p_input[18834]), .Z(n2594) );
  AND U3891 ( .A(p_input[8834]), .B(p_input[38834]), .Z(n2593) );
  AND U3892 ( .A(n2595), .B(n2596), .Z(o[8833]) );
  AND U3893 ( .A(p_input[28833]), .B(p_input[18833]), .Z(n2596) );
  AND U3894 ( .A(p_input[8833]), .B(p_input[38833]), .Z(n2595) );
  AND U3895 ( .A(n2597), .B(n2598), .Z(o[8832]) );
  AND U3896 ( .A(p_input[28832]), .B(p_input[18832]), .Z(n2598) );
  AND U3897 ( .A(p_input[8832]), .B(p_input[38832]), .Z(n2597) );
  AND U3898 ( .A(n2599), .B(n2600), .Z(o[8831]) );
  AND U3899 ( .A(p_input[28831]), .B(p_input[18831]), .Z(n2600) );
  AND U3900 ( .A(p_input[8831]), .B(p_input[38831]), .Z(n2599) );
  AND U3901 ( .A(n2601), .B(n2602), .Z(o[8830]) );
  AND U3902 ( .A(p_input[28830]), .B(p_input[18830]), .Z(n2602) );
  AND U3903 ( .A(p_input[8830]), .B(p_input[38830]), .Z(n2601) );
  AND U3904 ( .A(n2603), .B(n2604), .Z(o[882]) );
  AND U3905 ( .A(p_input[20882]), .B(p_input[10882]), .Z(n2604) );
  AND U3906 ( .A(p_input[882]), .B(p_input[30882]), .Z(n2603) );
  AND U3907 ( .A(n2605), .B(n2606), .Z(o[8829]) );
  AND U3908 ( .A(p_input[28829]), .B(p_input[18829]), .Z(n2606) );
  AND U3909 ( .A(p_input[8829]), .B(p_input[38829]), .Z(n2605) );
  AND U3910 ( .A(n2607), .B(n2608), .Z(o[8828]) );
  AND U3911 ( .A(p_input[28828]), .B(p_input[18828]), .Z(n2608) );
  AND U3912 ( .A(p_input[8828]), .B(p_input[38828]), .Z(n2607) );
  AND U3913 ( .A(n2609), .B(n2610), .Z(o[8827]) );
  AND U3914 ( .A(p_input[28827]), .B(p_input[18827]), .Z(n2610) );
  AND U3915 ( .A(p_input[8827]), .B(p_input[38827]), .Z(n2609) );
  AND U3916 ( .A(n2611), .B(n2612), .Z(o[8826]) );
  AND U3917 ( .A(p_input[28826]), .B(p_input[18826]), .Z(n2612) );
  AND U3918 ( .A(p_input[8826]), .B(p_input[38826]), .Z(n2611) );
  AND U3919 ( .A(n2613), .B(n2614), .Z(o[8825]) );
  AND U3920 ( .A(p_input[28825]), .B(p_input[18825]), .Z(n2614) );
  AND U3921 ( .A(p_input[8825]), .B(p_input[38825]), .Z(n2613) );
  AND U3922 ( .A(n2615), .B(n2616), .Z(o[8824]) );
  AND U3923 ( .A(p_input[28824]), .B(p_input[18824]), .Z(n2616) );
  AND U3924 ( .A(p_input[8824]), .B(p_input[38824]), .Z(n2615) );
  AND U3925 ( .A(n2617), .B(n2618), .Z(o[8823]) );
  AND U3926 ( .A(p_input[28823]), .B(p_input[18823]), .Z(n2618) );
  AND U3927 ( .A(p_input[8823]), .B(p_input[38823]), .Z(n2617) );
  AND U3928 ( .A(n2619), .B(n2620), .Z(o[8822]) );
  AND U3929 ( .A(p_input[28822]), .B(p_input[18822]), .Z(n2620) );
  AND U3930 ( .A(p_input[8822]), .B(p_input[38822]), .Z(n2619) );
  AND U3931 ( .A(n2621), .B(n2622), .Z(o[8821]) );
  AND U3932 ( .A(p_input[28821]), .B(p_input[18821]), .Z(n2622) );
  AND U3933 ( .A(p_input[8821]), .B(p_input[38821]), .Z(n2621) );
  AND U3934 ( .A(n2623), .B(n2624), .Z(o[8820]) );
  AND U3935 ( .A(p_input[28820]), .B(p_input[18820]), .Z(n2624) );
  AND U3936 ( .A(p_input[8820]), .B(p_input[38820]), .Z(n2623) );
  AND U3937 ( .A(n2625), .B(n2626), .Z(o[881]) );
  AND U3938 ( .A(p_input[20881]), .B(p_input[10881]), .Z(n2626) );
  AND U3939 ( .A(p_input[881]), .B(p_input[30881]), .Z(n2625) );
  AND U3940 ( .A(n2627), .B(n2628), .Z(o[8819]) );
  AND U3941 ( .A(p_input[28819]), .B(p_input[18819]), .Z(n2628) );
  AND U3942 ( .A(p_input[8819]), .B(p_input[38819]), .Z(n2627) );
  AND U3943 ( .A(n2629), .B(n2630), .Z(o[8818]) );
  AND U3944 ( .A(p_input[28818]), .B(p_input[18818]), .Z(n2630) );
  AND U3945 ( .A(p_input[8818]), .B(p_input[38818]), .Z(n2629) );
  AND U3946 ( .A(n2631), .B(n2632), .Z(o[8817]) );
  AND U3947 ( .A(p_input[28817]), .B(p_input[18817]), .Z(n2632) );
  AND U3948 ( .A(p_input[8817]), .B(p_input[38817]), .Z(n2631) );
  AND U3949 ( .A(n2633), .B(n2634), .Z(o[8816]) );
  AND U3950 ( .A(p_input[28816]), .B(p_input[18816]), .Z(n2634) );
  AND U3951 ( .A(p_input[8816]), .B(p_input[38816]), .Z(n2633) );
  AND U3952 ( .A(n2635), .B(n2636), .Z(o[8815]) );
  AND U3953 ( .A(p_input[28815]), .B(p_input[18815]), .Z(n2636) );
  AND U3954 ( .A(p_input[8815]), .B(p_input[38815]), .Z(n2635) );
  AND U3955 ( .A(n2637), .B(n2638), .Z(o[8814]) );
  AND U3956 ( .A(p_input[28814]), .B(p_input[18814]), .Z(n2638) );
  AND U3957 ( .A(p_input[8814]), .B(p_input[38814]), .Z(n2637) );
  AND U3958 ( .A(n2639), .B(n2640), .Z(o[8813]) );
  AND U3959 ( .A(p_input[28813]), .B(p_input[18813]), .Z(n2640) );
  AND U3960 ( .A(p_input[8813]), .B(p_input[38813]), .Z(n2639) );
  AND U3961 ( .A(n2641), .B(n2642), .Z(o[8812]) );
  AND U3962 ( .A(p_input[28812]), .B(p_input[18812]), .Z(n2642) );
  AND U3963 ( .A(p_input[8812]), .B(p_input[38812]), .Z(n2641) );
  AND U3964 ( .A(n2643), .B(n2644), .Z(o[8811]) );
  AND U3965 ( .A(p_input[28811]), .B(p_input[18811]), .Z(n2644) );
  AND U3966 ( .A(p_input[8811]), .B(p_input[38811]), .Z(n2643) );
  AND U3967 ( .A(n2645), .B(n2646), .Z(o[8810]) );
  AND U3968 ( .A(p_input[28810]), .B(p_input[18810]), .Z(n2646) );
  AND U3969 ( .A(p_input[8810]), .B(p_input[38810]), .Z(n2645) );
  AND U3970 ( .A(n2647), .B(n2648), .Z(o[880]) );
  AND U3971 ( .A(p_input[20880]), .B(p_input[10880]), .Z(n2648) );
  AND U3972 ( .A(p_input[880]), .B(p_input[30880]), .Z(n2647) );
  AND U3973 ( .A(n2649), .B(n2650), .Z(o[8809]) );
  AND U3974 ( .A(p_input[28809]), .B(p_input[18809]), .Z(n2650) );
  AND U3975 ( .A(p_input[8809]), .B(p_input[38809]), .Z(n2649) );
  AND U3976 ( .A(n2651), .B(n2652), .Z(o[8808]) );
  AND U3977 ( .A(p_input[28808]), .B(p_input[18808]), .Z(n2652) );
  AND U3978 ( .A(p_input[8808]), .B(p_input[38808]), .Z(n2651) );
  AND U3979 ( .A(n2653), .B(n2654), .Z(o[8807]) );
  AND U3980 ( .A(p_input[28807]), .B(p_input[18807]), .Z(n2654) );
  AND U3981 ( .A(p_input[8807]), .B(p_input[38807]), .Z(n2653) );
  AND U3982 ( .A(n2655), .B(n2656), .Z(o[8806]) );
  AND U3983 ( .A(p_input[28806]), .B(p_input[18806]), .Z(n2656) );
  AND U3984 ( .A(p_input[8806]), .B(p_input[38806]), .Z(n2655) );
  AND U3985 ( .A(n2657), .B(n2658), .Z(o[8805]) );
  AND U3986 ( .A(p_input[28805]), .B(p_input[18805]), .Z(n2658) );
  AND U3987 ( .A(p_input[8805]), .B(p_input[38805]), .Z(n2657) );
  AND U3988 ( .A(n2659), .B(n2660), .Z(o[8804]) );
  AND U3989 ( .A(p_input[28804]), .B(p_input[18804]), .Z(n2660) );
  AND U3990 ( .A(p_input[8804]), .B(p_input[38804]), .Z(n2659) );
  AND U3991 ( .A(n2661), .B(n2662), .Z(o[8803]) );
  AND U3992 ( .A(p_input[28803]), .B(p_input[18803]), .Z(n2662) );
  AND U3993 ( .A(p_input[8803]), .B(p_input[38803]), .Z(n2661) );
  AND U3994 ( .A(n2663), .B(n2664), .Z(o[8802]) );
  AND U3995 ( .A(p_input[28802]), .B(p_input[18802]), .Z(n2664) );
  AND U3996 ( .A(p_input[8802]), .B(p_input[38802]), .Z(n2663) );
  AND U3997 ( .A(n2665), .B(n2666), .Z(o[8801]) );
  AND U3998 ( .A(p_input[28801]), .B(p_input[18801]), .Z(n2666) );
  AND U3999 ( .A(p_input[8801]), .B(p_input[38801]), .Z(n2665) );
  AND U4000 ( .A(n2667), .B(n2668), .Z(o[8800]) );
  AND U4001 ( .A(p_input[28800]), .B(p_input[18800]), .Z(n2668) );
  AND U4002 ( .A(p_input[8800]), .B(p_input[38800]), .Z(n2667) );
  AND U4003 ( .A(n2669), .B(n2670), .Z(o[87]) );
  AND U4004 ( .A(p_input[20087]), .B(p_input[10087]), .Z(n2670) );
  AND U4005 ( .A(p_input[87]), .B(p_input[30087]), .Z(n2669) );
  AND U4006 ( .A(n2671), .B(n2672), .Z(o[879]) );
  AND U4007 ( .A(p_input[20879]), .B(p_input[10879]), .Z(n2672) );
  AND U4008 ( .A(p_input[879]), .B(p_input[30879]), .Z(n2671) );
  AND U4009 ( .A(n2673), .B(n2674), .Z(o[8799]) );
  AND U4010 ( .A(p_input[28799]), .B(p_input[18799]), .Z(n2674) );
  AND U4011 ( .A(p_input[8799]), .B(p_input[38799]), .Z(n2673) );
  AND U4012 ( .A(n2675), .B(n2676), .Z(o[8798]) );
  AND U4013 ( .A(p_input[28798]), .B(p_input[18798]), .Z(n2676) );
  AND U4014 ( .A(p_input[8798]), .B(p_input[38798]), .Z(n2675) );
  AND U4015 ( .A(n2677), .B(n2678), .Z(o[8797]) );
  AND U4016 ( .A(p_input[28797]), .B(p_input[18797]), .Z(n2678) );
  AND U4017 ( .A(p_input[8797]), .B(p_input[38797]), .Z(n2677) );
  AND U4018 ( .A(n2679), .B(n2680), .Z(o[8796]) );
  AND U4019 ( .A(p_input[28796]), .B(p_input[18796]), .Z(n2680) );
  AND U4020 ( .A(p_input[8796]), .B(p_input[38796]), .Z(n2679) );
  AND U4021 ( .A(n2681), .B(n2682), .Z(o[8795]) );
  AND U4022 ( .A(p_input[28795]), .B(p_input[18795]), .Z(n2682) );
  AND U4023 ( .A(p_input[8795]), .B(p_input[38795]), .Z(n2681) );
  AND U4024 ( .A(n2683), .B(n2684), .Z(o[8794]) );
  AND U4025 ( .A(p_input[28794]), .B(p_input[18794]), .Z(n2684) );
  AND U4026 ( .A(p_input[8794]), .B(p_input[38794]), .Z(n2683) );
  AND U4027 ( .A(n2685), .B(n2686), .Z(o[8793]) );
  AND U4028 ( .A(p_input[28793]), .B(p_input[18793]), .Z(n2686) );
  AND U4029 ( .A(p_input[8793]), .B(p_input[38793]), .Z(n2685) );
  AND U4030 ( .A(n2687), .B(n2688), .Z(o[8792]) );
  AND U4031 ( .A(p_input[28792]), .B(p_input[18792]), .Z(n2688) );
  AND U4032 ( .A(p_input[8792]), .B(p_input[38792]), .Z(n2687) );
  AND U4033 ( .A(n2689), .B(n2690), .Z(o[8791]) );
  AND U4034 ( .A(p_input[28791]), .B(p_input[18791]), .Z(n2690) );
  AND U4035 ( .A(p_input[8791]), .B(p_input[38791]), .Z(n2689) );
  AND U4036 ( .A(n2691), .B(n2692), .Z(o[8790]) );
  AND U4037 ( .A(p_input[28790]), .B(p_input[18790]), .Z(n2692) );
  AND U4038 ( .A(p_input[8790]), .B(p_input[38790]), .Z(n2691) );
  AND U4039 ( .A(n2693), .B(n2694), .Z(o[878]) );
  AND U4040 ( .A(p_input[20878]), .B(p_input[10878]), .Z(n2694) );
  AND U4041 ( .A(p_input[878]), .B(p_input[30878]), .Z(n2693) );
  AND U4042 ( .A(n2695), .B(n2696), .Z(o[8789]) );
  AND U4043 ( .A(p_input[28789]), .B(p_input[18789]), .Z(n2696) );
  AND U4044 ( .A(p_input[8789]), .B(p_input[38789]), .Z(n2695) );
  AND U4045 ( .A(n2697), .B(n2698), .Z(o[8788]) );
  AND U4046 ( .A(p_input[28788]), .B(p_input[18788]), .Z(n2698) );
  AND U4047 ( .A(p_input[8788]), .B(p_input[38788]), .Z(n2697) );
  AND U4048 ( .A(n2699), .B(n2700), .Z(o[8787]) );
  AND U4049 ( .A(p_input[28787]), .B(p_input[18787]), .Z(n2700) );
  AND U4050 ( .A(p_input[8787]), .B(p_input[38787]), .Z(n2699) );
  AND U4051 ( .A(n2701), .B(n2702), .Z(o[8786]) );
  AND U4052 ( .A(p_input[28786]), .B(p_input[18786]), .Z(n2702) );
  AND U4053 ( .A(p_input[8786]), .B(p_input[38786]), .Z(n2701) );
  AND U4054 ( .A(n2703), .B(n2704), .Z(o[8785]) );
  AND U4055 ( .A(p_input[28785]), .B(p_input[18785]), .Z(n2704) );
  AND U4056 ( .A(p_input[8785]), .B(p_input[38785]), .Z(n2703) );
  AND U4057 ( .A(n2705), .B(n2706), .Z(o[8784]) );
  AND U4058 ( .A(p_input[28784]), .B(p_input[18784]), .Z(n2706) );
  AND U4059 ( .A(p_input[8784]), .B(p_input[38784]), .Z(n2705) );
  AND U4060 ( .A(n2707), .B(n2708), .Z(o[8783]) );
  AND U4061 ( .A(p_input[28783]), .B(p_input[18783]), .Z(n2708) );
  AND U4062 ( .A(p_input[8783]), .B(p_input[38783]), .Z(n2707) );
  AND U4063 ( .A(n2709), .B(n2710), .Z(o[8782]) );
  AND U4064 ( .A(p_input[28782]), .B(p_input[18782]), .Z(n2710) );
  AND U4065 ( .A(p_input[8782]), .B(p_input[38782]), .Z(n2709) );
  AND U4066 ( .A(n2711), .B(n2712), .Z(o[8781]) );
  AND U4067 ( .A(p_input[28781]), .B(p_input[18781]), .Z(n2712) );
  AND U4068 ( .A(p_input[8781]), .B(p_input[38781]), .Z(n2711) );
  AND U4069 ( .A(n2713), .B(n2714), .Z(o[8780]) );
  AND U4070 ( .A(p_input[28780]), .B(p_input[18780]), .Z(n2714) );
  AND U4071 ( .A(p_input[8780]), .B(p_input[38780]), .Z(n2713) );
  AND U4072 ( .A(n2715), .B(n2716), .Z(o[877]) );
  AND U4073 ( .A(p_input[20877]), .B(p_input[10877]), .Z(n2716) );
  AND U4074 ( .A(p_input[877]), .B(p_input[30877]), .Z(n2715) );
  AND U4075 ( .A(n2717), .B(n2718), .Z(o[8779]) );
  AND U4076 ( .A(p_input[28779]), .B(p_input[18779]), .Z(n2718) );
  AND U4077 ( .A(p_input[8779]), .B(p_input[38779]), .Z(n2717) );
  AND U4078 ( .A(n2719), .B(n2720), .Z(o[8778]) );
  AND U4079 ( .A(p_input[28778]), .B(p_input[18778]), .Z(n2720) );
  AND U4080 ( .A(p_input[8778]), .B(p_input[38778]), .Z(n2719) );
  AND U4081 ( .A(n2721), .B(n2722), .Z(o[8777]) );
  AND U4082 ( .A(p_input[28777]), .B(p_input[18777]), .Z(n2722) );
  AND U4083 ( .A(p_input[8777]), .B(p_input[38777]), .Z(n2721) );
  AND U4084 ( .A(n2723), .B(n2724), .Z(o[8776]) );
  AND U4085 ( .A(p_input[28776]), .B(p_input[18776]), .Z(n2724) );
  AND U4086 ( .A(p_input[8776]), .B(p_input[38776]), .Z(n2723) );
  AND U4087 ( .A(n2725), .B(n2726), .Z(o[8775]) );
  AND U4088 ( .A(p_input[28775]), .B(p_input[18775]), .Z(n2726) );
  AND U4089 ( .A(p_input[8775]), .B(p_input[38775]), .Z(n2725) );
  AND U4090 ( .A(n2727), .B(n2728), .Z(o[8774]) );
  AND U4091 ( .A(p_input[28774]), .B(p_input[18774]), .Z(n2728) );
  AND U4092 ( .A(p_input[8774]), .B(p_input[38774]), .Z(n2727) );
  AND U4093 ( .A(n2729), .B(n2730), .Z(o[8773]) );
  AND U4094 ( .A(p_input[28773]), .B(p_input[18773]), .Z(n2730) );
  AND U4095 ( .A(p_input[8773]), .B(p_input[38773]), .Z(n2729) );
  AND U4096 ( .A(n2731), .B(n2732), .Z(o[8772]) );
  AND U4097 ( .A(p_input[28772]), .B(p_input[18772]), .Z(n2732) );
  AND U4098 ( .A(p_input[8772]), .B(p_input[38772]), .Z(n2731) );
  AND U4099 ( .A(n2733), .B(n2734), .Z(o[8771]) );
  AND U4100 ( .A(p_input[28771]), .B(p_input[18771]), .Z(n2734) );
  AND U4101 ( .A(p_input[8771]), .B(p_input[38771]), .Z(n2733) );
  AND U4102 ( .A(n2735), .B(n2736), .Z(o[8770]) );
  AND U4103 ( .A(p_input[28770]), .B(p_input[18770]), .Z(n2736) );
  AND U4104 ( .A(p_input[8770]), .B(p_input[38770]), .Z(n2735) );
  AND U4105 ( .A(n2737), .B(n2738), .Z(o[876]) );
  AND U4106 ( .A(p_input[20876]), .B(p_input[10876]), .Z(n2738) );
  AND U4107 ( .A(p_input[876]), .B(p_input[30876]), .Z(n2737) );
  AND U4108 ( .A(n2739), .B(n2740), .Z(o[8769]) );
  AND U4109 ( .A(p_input[28769]), .B(p_input[18769]), .Z(n2740) );
  AND U4110 ( .A(p_input[8769]), .B(p_input[38769]), .Z(n2739) );
  AND U4111 ( .A(n2741), .B(n2742), .Z(o[8768]) );
  AND U4112 ( .A(p_input[28768]), .B(p_input[18768]), .Z(n2742) );
  AND U4113 ( .A(p_input[8768]), .B(p_input[38768]), .Z(n2741) );
  AND U4114 ( .A(n2743), .B(n2744), .Z(o[8767]) );
  AND U4115 ( .A(p_input[28767]), .B(p_input[18767]), .Z(n2744) );
  AND U4116 ( .A(p_input[8767]), .B(p_input[38767]), .Z(n2743) );
  AND U4117 ( .A(n2745), .B(n2746), .Z(o[8766]) );
  AND U4118 ( .A(p_input[28766]), .B(p_input[18766]), .Z(n2746) );
  AND U4119 ( .A(p_input[8766]), .B(p_input[38766]), .Z(n2745) );
  AND U4120 ( .A(n2747), .B(n2748), .Z(o[8765]) );
  AND U4121 ( .A(p_input[28765]), .B(p_input[18765]), .Z(n2748) );
  AND U4122 ( .A(p_input[8765]), .B(p_input[38765]), .Z(n2747) );
  AND U4123 ( .A(n2749), .B(n2750), .Z(o[8764]) );
  AND U4124 ( .A(p_input[28764]), .B(p_input[18764]), .Z(n2750) );
  AND U4125 ( .A(p_input[8764]), .B(p_input[38764]), .Z(n2749) );
  AND U4126 ( .A(n2751), .B(n2752), .Z(o[8763]) );
  AND U4127 ( .A(p_input[28763]), .B(p_input[18763]), .Z(n2752) );
  AND U4128 ( .A(p_input[8763]), .B(p_input[38763]), .Z(n2751) );
  AND U4129 ( .A(n2753), .B(n2754), .Z(o[8762]) );
  AND U4130 ( .A(p_input[28762]), .B(p_input[18762]), .Z(n2754) );
  AND U4131 ( .A(p_input[8762]), .B(p_input[38762]), .Z(n2753) );
  AND U4132 ( .A(n2755), .B(n2756), .Z(o[8761]) );
  AND U4133 ( .A(p_input[28761]), .B(p_input[18761]), .Z(n2756) );
  AND U4134 ( .A(p_input[8761]), .B(p_input[38761]), .Z(n2755) );
  AND U4135 ( .A(n2757), .B(n2758), .Z(o[8760]) );
  AND U4136 ( .A(p_input[28760]), .B(p_input[18760]), .Z(n2758) );
  AND U4137 ( .A(p_input[8760]), .B(p_input[38760]), .Z(n2757) );
  AND U4138 ( .A(n2759), .B(n2760), .Z(o[875]) );
  AND U4139 ( .A(p_input[20875]), .B(p_input[10875]), .Z(n2760) );
  AND U4140 ( .A(p_input[875]), .B(p_input[30875]), .Z(n2759) );
  AND U4141 ( .A(n2761), .B(n2762), .Z(o[8759]) );
  AND U4142 ( .A(p_input[28759]), .B(p_input[18759]), .Z(n2762) );
  AND U4143 ( .A(p_input[8759]), .B(p_input[38759]), .Z(n2761) );
  AND U4144 ( .A(n2763), .B(n2764), .Z(o[8758]) );
  AND U4145 ( .A(p_input[28758]), .B(p_input[18758]), .Z(n2764) );
  AND U4146 ( .A(p_input[8758]), .B(p_input[38758]), .Z(n2763) );
  AND U4147 ( .A(n2765), .B(n2766), .Z(o[8757]) );
  AND U4148 ( .A(p_input[28757]), .B(p_input[18757]), .Z(n2766) );
  AND U4149 ( .A(p_input[8757]), .B(p_input[38757]), .Z(n2765) );
  AND U4150 ( .A(n2767), .B(n2768), .Z(o[8756]) );
  AND U4151 ( .A(p_input[28756]), .B(p_input[18756]), .Z(n2768) );
  AND U4152 ( .A(p_input[8756]), .B(p_input[38756]), .Z(n2767) );
  AND U4153 ( .A(n2769), .B(n2770), .Z(o[8755]) );
  AND U4154 ( .A(p_input[28755]), .B(p_input[18755]), .Z(n2770) );
  AND U4155 ( .A(p_input[8755]), .B(p_input[38755]), .Z(n2769) );
  AND U4156 ( .A(n2771), .B(n2772), .Z(o[8754]) );
  AND U4157 ( .A(p_input[28754]), .B(p_input[18754]), .Z(n2772) );
  AND U4158 ( .A(p_input[8754]), .B(p_input[38754]), .Z(n2771) );
  AND U4159 ( .A(n2773), .B(n2774), .Z(o[8753]) );
  AND U4160 ( .A(p_input[28753]), .B(p_input[18753]), .Z(n2774) );
  AND U4161 ( .A(p_input[8753]), .B(p_input[38753]), .Z(n2773) );
  AND U4162 ( .A(n2775), .B(n2776), .Z(o[8752]) );
  AND U4163 ( .A(p_input[28752]), .B(p_input[18752]), .Z(n2776) );
  AND U4164 ( .A(p_input[8752]), .B(p_input[38752]), .Z(n2775) );
  AND U4165 ( .A(n2777), .B(n2778), .Z(o[8751]) );
  AND U4166 ( .A(p_input[28751]), .B(p_input[18751]), .Z(n2778) );
  AND U4167 ( .A(p_input[8751]), .B(p_input[38751]), .Z(n2777) );
  AND U4168 ( .A(n2779), .B(n2780), .Z(o[8750]) );
  AND U4169 ( .A(p_input[28750]), .B(p_input[18750]), .Z(n2780) );
  AND U4170 ( .A(p_input[8750]), .B(p_input[38750]), .Z(n2779) );
  AND U4171 ( .A(n2781), .B(n2782), .Z(o[874]) );
  AND U4172 ( .A(p_input[20874]), .B(p_input[10874]), .Z(n2782) );
  AND U4173 ( .A(p_input[874]), .B(p_input[30874]), .Z(n2781) );
  AND U4174 ( .A(n2783), .B(n2784), .Z(o[8749]) );
  AND U4175 ( .A(p_input[28749]), .B(p_input[18749]), .Z(n2784) );
  AND U4176 ( .A(p_input[8749]), .B(p_input[38749]), .Z(n2783) );
  AND U4177 ( .A(n2785), .B(n2786), .Z(o[8748]) );
  AND U4178 ( .A(p_input[28748]), .B(p_input[18748]), .Z(n2786) );
  AND U4179 ( .A(p_input[8748]), .B(p_input[38748]), .Z(n2785) );
  AND U4180 ( .A(n2787), .B(n2788), .Z(o[8747]) );
  AND U4181 ( .A(p_input[28747]), .B(p_input[18747]), .Z(n2788) );
  AND U4182 ( .A(p_input[8747]), .B(p_input[38747]), .Z(n2787) );
  AND U4183 ( .A(n2789), .B(n2790), .Z(o[8746]) );
  AND U4184 ( .A(p_input[28746]), .B(p_input[18746]), .Z(n2790) );
  AND U4185 ( .A(p_input[8746]), .B(p_input[38746]), .Z(n2789) );
  AND U4186 ( .A(n2791), .B(n2792), .Z(o[8745]) );
  AND U4187 ( .A(p_input[28745]), .B(p_input[18745]), .Z(n2792) );
  AND U4188 ( .A(p_input[8745]), .B(p_input[38745]), .Z(n2791) );
  AND U4189 ( .A(n2793), .B(n2794), .Z(o[8744]) );
  AND U4190 ( .A(p_input[28744]), .B(p_input[18744]), .Z(n2794) );
  AND U4191 ( .A(p_input[8744]), .B(p_input[38744]), .Z(n2793) );
  AND U4192 ( .A(n2795), .B(n2796), .Z(o[8743]) );
  AND U4193 ( .A(p_input[28743]), .B(p_input[18743]), .Z(n2796) );
  AND U4194 ( .A(p_input[8743]), .B(p_input[38743]), .Z(n2795) );
  AND U4195 ( .A(n2797), .B(n2798), .Z(o[8742]) );
  AND U4196 ( .A(p_input[28742]), .B(p_input[18742]), .Z(n2798) );
  AND U4197 ( .A(p_input[8742]), .B(p_input[38742]), .Z(n2797) );
  AND U4198 ( .A(n2799), .B(n2800), .Z(o[8741]) );
  AND U4199 ( .A(p_input[28741]), .B(p_input[18741]), .Z(n2800) );
  AND U4200 ( .A(p_input[8741]), .B(p_input[38741]), .Z(n2799) );
  AND U4201 ( .A(n2801), .B(n2802), .Z(o[8740]) );
  AND U4202 ( .A(p_input[28740]), .B(p_input[18740]), .Z(n2802) );
  AND U4203 ( .A(p_input[8740]), .B(p_input[38740]), .Z(n2801) );
  AND U4204 ( .A(n2803), .B(n2804), .Z(o[873]) );
  AND U4205 ( .A(p_input[20873]), .B(p_input[10873]), .Z(n2804) );
  AND U4206 ( .A(p_input[873]), .B(p_input[30873]), .Z(n2803) );
  AND U4207 ( .A(n2805), .B(n2806), .Z(o[8739]) );
  AND U4208 ( .A(p_input[28739]), .B(p_input[18739]), .Z(n2806) );
  AND U4209 ( .A(p_input[8739]), .B(p_input[38739]), .Z(n2805) );
  AND U4210 ( .A(n2807), .B(n2808), .Z(o[8738]) );
  AND U4211 ( .A(p_input[28738]), .B(p_input[18738]), .Z(n2808) );
  AND U4212 ( .A(p_input[8738]), .B(p_input[38738]), .Z(n2807) );
  AND U4213 ( .A(n2809), .B(n2810), .Z(o[8737]) );
  AND U4214 ( .A(p_input[28737]), .B(p_input[18737]), .Z(n2810) );
  AND U4215 ( .A(p_input[8737]), .B(p_input[38737]), .Z(n2809) );
  AND U4216 ( .A(n2811), .B(n2812), .Z(o[8736]) );
  AND U4217 ( .A(p_input[28736]), .B(p_input[18736]), .Z(n2812) );
  AND U4218 ( .A(p_input[8736]), .B(p_input[38736]), .Z(n2811) );
  AND U4219 ( .A(n2813), .B(n2814), .Z(o[8735]) );
  AND U4220 ( .A(p_input[28735]), .B(p_input[18735]), .Z(n2814) );
  AND U4221 ( .A(p_input[8735]), .B(p_input[38735]), .Z(n2813) );
  AND U4222 ( .A(n2815), .B(n2816), .Z(o[8734]) );
  AND U4223 ( .A(p_input[28734]), .B(p_input[18734]), .Z(n2816) );
  AND U4224 ( .A(p_input[8734]), .B(p_input[38734]), .Z(n2815) );
  AND U4225 ( .A(n2817), .B(n2818), .Z(o[8733]) );
  AND U4226 ( .A(p_input[28733]), .B(p_input[18733]), .Z(n2818) );
  AND U4227 ( .A(p_input[8733]), .B(p_input[38733]), .Z(n2817) );
  AND U4228 ( .A(n2819), .B(n2820), .Z(o[8732]) );
  AND U4229 ( .A(p_input[28732]), .B(p_input[18732]), .Z(n2820) );
  AND U4230 ( .A(p_input[8732]), .B(p_input[38732]), .Z(n2819) );
  AND U4231 ( .A(n2821), .B(n2822), .Z(o[8731]) );
  AND U4232 ( .A(p_input[28731]), .B(p_input[18731]), .Z(n2822) );
  AND U4233 ( .A(p_input[8731]), .B(p_input[38731]), .Z(n2821) );
  AND U4234 ( .A(n2823), .B(n2824), .Z(o[8730]) );
  AND U4235 ( .A(p_input[28730]), .B(p_input[18730]), .Z(n2824) );
  AND U4236 ( .A(p_input[8730]), .B(p_input[38730]), .Z(n2823) );
  AND U4237 ( .A(n2825), .B(n2826), .Z(o[872]) );
  AND U4238 ( .A(p_input[20872]), .B(p_input[10872]), .Z(n2826) );
  AND U4239 ( .A(p_input[872]), .B(p_input[30872]), .Z(n2825) );
  AND U4240 ( .A(n2827), .B(n2828), .Z(o[8729]) );
  AND U4241 ( .A(p_input[28729]), .B(p_input[18729]), .Z(n2828) );
  AND U4242 ( .A(p_input[8729]), .B(p_input[38729]), .Z(n2827) );
  AND U4243 ( .A(n2829), .B(n2830), .Z(o[8728]) );
  AND U4244 ( .A(p_input[28728]), .B(p_input[18728]), .Z(n2830) );
  AND U4245 ( .A(p_input[8728]), .B(p_input[38728]), .Z(n2829) );
  AND U4246 ( .A(n2831), .B(n2832), .Z(o[8727]) );
  AND U4247 ( .A(p_input[28727]), .B(p_input[18727]), .Z(n2832) );
  AND U4248 ( .A(p_input[8727]), .B(p_input[38727]), .Z(n2831) );
  AND U4249 ( .A(n2833), .B(n2834), .Z(o[8726]) );
  AND U4250 ( .A(p_input[28726]), .B(p_input[18726]), .Z(n2834) );
  AND U4251 ( .A(p_input[8726]), .B(p_input[38726]), .Z(n2833) );
  AND U4252 ( .A(n2835), .B(n2836), .Z(o[8725]) );
  AND U4253 ( .A(p_input[28725]), .B(p_input[18725]), .Z(n2836) );
  AND U4254 ( .A(p_input[8725]), .B(p_input[38725]), .Z(n2835) );
  AND U4255 ( .A(n2837), .B(n2838), .Z(o[8724]) );
  AND U4256 ( .A(p_input[28724]), .B(p_input[18724]), .Z(n2838) );
  AND U4257 ( .A(p_input[8724]), .B(p_input[38724]), .Z(n2837) );
  AND U4258 ( .A(n2839), .B(n2840), .Z(o[8723]) );
  AND U4259 ( .A(p_input[28723]), .B(p_input[18723]), .Z(n2840) );
  AND U4260 ( .A(p_input[8723]), .B(p_input[38723]), .Z(n2839) );
  AND U4261 ( .A(n2841), .B(n2842), .Z(o[8722]) );
  AND U4262 ( .A(p_input[28722]), .B(p_input[18722]), .Z(n2842) );
  AND U4263 ( .A(p_input[8722]), .B(p_input[38722]), .Z(n2841) );
  AND U4264 ( .A(n2843), .B(n2844), .Z(o[8721]) );
  AND U4265 ( .A(p_input[28721]), .B(p_input[18721]), .Z(n2844) );
  AND U4266 ( .A(p_input[8721]), .B(p_input[38721]), .Z(n2843) );
  AND U4267 ( .A(n2845), .B(n2846), .Z(o[8720]) );
  AND U4268 ( .A(p_input[28720]), .B(p_input[18720]), .Z(n2846) );
  AND U4269 ( .A(p_input[8720]), .B(p_input[38720]), .Z(n2845) );
  AND U4270 ( .A(n2847), .B(n2848), .Z(o[871]) );
  AND U4271 ( .A(p_input[20871]), .B(p_input[10871]), .Z(n2848) );
  AND U4272 ( .A(p_input[871]), .B(p_input[30871]), .Z(n2847) );
  AND U4273 ( .A(n2849), .B(n2850), .Z(o[8719]) );
  AND U4274 ( .A(p_input[28719]), .B(p_input[18719]), .Z(n2850) );
  AND U4275 ( .A(p_input[8719]), .B(p_input[38719]), .Z(n2849) );
  AND U4276 ( .A(n2851), .B(n2852), .Z(o[8718]) );
  AND U4277 ( .A(p_input[28718]), .B(p_input[18718]), .Z(n2852) );
  AND U4278 ( .A(p_input[8718]), .B(p_input[38718]), .Z(n2851) );
  AND U4279 ( .A(n2853), .B(n2854), .Z(o[8717]) );
  AND U4280 ( .A(p_input[28717]), .B(p_input[18717]), .Z(n2854) );
  AND U4281 ( .A(p_input[8717]), .B(p_input[38717]), .Z(n2853) );
  AND U4282 ( .A(n2855), .B(n2856), .Z(o[8716]) );
  AND U4283 ( .A(p_input[28716]), .B(p_input[18716]), .Z(n2856) );
  AND U4284 ( .A(p_input[8716]), .B(p_input[38716]), .Z(n2855) );
  AND U4285 ( .A(n2857), .B(n2858), .Z(o[8715]) );
  AND U4286 ( .A(p_input[28715]), .B(p_input[18715]), .Z(n2858) );
  AND U4287 ( .A(p_input[8715]), .B(p_input[38715]), .Z(n2857) );
  AND U4288 ( .A(n2859), .B(n2860), .Z(o[8714]) );
  AND U4289 ( .A(p_input[28714]), .B(p_input[18714]), .Z(n2860) );
  AND U4290 ( .A(p_input[8714]), .B(p_input[38714]), .Z(n2859) );
  AND U4291 ( .A(n2861), .B(n2862), .Z(o[8713]) );
  AND U4292 ( .A(p_input[28713]), .B(p_input[18713]), .Z(n2862) );
  AND U4293 ( .A(p_input[8713]), .B(p_input[38713]), .Z(n2861) );
  AND U4294 ( .A(n2863), .B(n2864), .Z(o[8712]) );
  AND U4295 ( .A(p_input[28712]), .B(p_input[18712]), .Z(n2864) );
  AND U4296 ( .A(p_input[8712]), .B(p_input[38712]), .Z(n2863) );
  AND U4297 ( .A(n2865), .B(n2866), .Z(o[8711]) );
  AND U4298 ( .A(p_input[28711]), .B(p_input[18711]), .Z(n2866) );
  AND U4299 ( .A(p_input[8711]), .B(p_input[38711]), .Z(n2865) );
  AND U4300 ( .A(n2867), .B(n2868), .Z(o[8710]) );
  AND U4301 ( .A(p_input[28710]), .B(p_input[18710]), .Z(n2868) );
  AND U4302 ( .A(p_input[8710]), .B(p_input[38710]), .Z(n2867) );
  AND U4303 ( .A(n2869), .B(n2870), .Z(o[870]) );
  AND U4304 ( .A(p_input[20870]), .B(p_input[10870]), .Z(n2870) );
  AND U4305 ( .A(p_input[870]), .B(p_input[30870]), .Z(n2869) );
  AND U4306 ( .A(n2871), .B(n2872), .Z(o[8709]) );
  AND U4307 ( .A(p_input[28709]), .B(p_input[18709]), .Z(n2872) );
  AND U4308 ( .A(p_input[8709]), .B(p_input[38709]), .Z(n2871) );
  AND U4309 ( .A(n2873), .B(n2874), .Z(o[8708]) );
  AND U4310 ( .A(p_input[28708]), .B(p_input[18708]), .Z(n2874) );
  AND U4311 ( .A(p_input[8708]), .B(p_input[38708]), .Z(n2873) );
  AND U4312 ( .A(n2875), .B(n2876), .Z(o[8707]) );
  AND U4313 ( .A(p_input[28707]), .B(p_input[18707]), .Z(n2876) );
  AND U4314 ( .A(p_input[8707]), .B(p_input[38707]), .Z(n2875) );
  AND U4315 ( .A(n2877), .B(n2878), .Z(o[8706]) );
  AND U4316 ( .A(p_input[28706]), .B(p_input[18706]), .Z(n2878) );
  AND U4317 ( .A(p_input[8706]), .B(p_input[38706]), .Z(n2877) );
  AND U4318 ( .A(n2879), .B(n2880), .Z(o[8705]) );
  AND U4319 ( .A(p_input[28705]), .B(p_input[18705]), .Z(n2880) );
  AND U4320 ( .A(p_input[8705]), .B(p_input[38705]), .Z(n2879) );
  AND U4321 ( .A(n2881), .B(n2882), .Z(o[8704]) );
  AND U4322 ( .A(p_input[28704]), .B(p_input[18704]), .Z(n2882) );
  AND U4323 ( .A(p_input[8704]), .B(p_input[38704]), .Z(n2881) );
  AND U4324 ( .A(n2883), .B(n2884), .Z(o[8703]) );
  AND U4325 ( .A(p_input[28703]), .B(p_input[18703]), .Z(n2884) );
  AND U4326 ( .A(p_input[8703]), .B(p_input[38703]), .Z(n2883) );
  AND U4327 ( .A(n2885), .B(n2886), .Z(o[8702]) );
  AND U4328 ( .A(p_input[28702]), .B(p_input[18702]), .Z(n2886) );
  AND U4329 ( .A(p_input[8702]), .B(p_input[38702]), .Z(n2885) );
  AND U4330 ( .A(n2887), .B(n2888), .Z(o[8701]) );
  AND U4331 ( .A(p_input[28701]), .B(p_input[18701]), .Z(n2888) );
  AND U4332 ( .A(p_input[8701]), .B(p_input[38701]), .Z(n2887) );
  AND U4333 ( .A(n2889), .B(n2890), .Z(o[8700]) );
  AND U4334 ( .A(p_input[28700]), .B(p_input[18700]), .Z(n2890) );
  AND U4335 ( .A(p_input[8700]), .B(p_input[38700]), .Z(n2889) );
  AND U4336 ( .A(n2891), .B(n2892), .Z(o[86]) );
  AND U4337 ( .A(p_input[20086]), .B(p_input[10086]), .Z(n2892) );
  AND U4338 ( .A(p_input[86]), .B(p_input[30086]), .Z(n2891) );
  AND U4339 ( .A(n2893), .B(n2894), .Z(o[869]) );
  AND U4340 ( .A(p_input[20869]), .B(p_input[10869]), .Z(n2894) );
  AND U4341 ( .A(p_input[869]), .B(p_input[30869]), .Z(n2893) );
  AND U4342 ( .A(n2895), .B(n2896), .Z(o[8699]) );
  AND U4343 ( .A(p_input[28699]), .B(p_input[18699]), .Z(n2896) );
  AND U4344 ( .A(p_input[8699]), .B(p_input[38699]), .Z(n2895) );
  AND U4345 ( .A(n2897), .B(n2898), .Z(o[8698]) );
  AND U4346 ( .A(p_input[28698]), .B(p_input[18698]), .Z(n2898) );
  AND U4347 ( .A(p_input[8698]), .B(p_input[38698]), .Z(n2897) );
  AND U4348 ( .A(n2899), .B(n2900), .Z(o[8697]) );
  AND U4349 ( .A(p_input[28697]), .B(p_input[18697]), .Z(n2900) );
  AND U4350 ( .A(p_input[8697]), .B(p_input[38697]), .Z(n2899) );
  AND U4351 ( .A(n2901), .B(n2902), .Z(o[8696]) );
  AND U4352 ( .A(p_input[28696]), .B(p_input[18696]), .Z(n2902) );
  AND U4353 ( .A(p_input[8696]), .B(p_input[38696]), .Z(n2901) );
  AND U4354 ( .A(n2903), .B(n2904), .Z(o[8695]) );
  AND U4355 ( .A(p_input[28695]), .B(p_input[18695]), .Z(n2904) );
  AND U4356 ( .A(p_input[8695]), .B(p_input[38695]), .Z(n2903) );
  AND U4357 ( .A(n2905), .B(n2906), .Z(o[8694]) );
  AND U4358 ( .A(p_input[28694]), .B(p_input[18694]), .Z(n2906) );
  AND U4359 ( .A(p_input[8694]), .B(p_input[38694]), .Z(n2905) );
  AND U4360 ( .A(n2907), .B(n2908), .Z(o[8693]) );
  AND U4361 ( .A(p_input[28693]), .B(p_input[18693]), .Z(n2908) );
  AND U4362 ( .A(p_input[8693]), .B(p_input[38693]), .Z(n2907) );
  AND U4363 ( .A(n2909), .B(n2910), .Z(o[8692]) );
  AND U4364 ( .A(p_input[28692]), .B(p_input[18692]), .Z(n2910) );
  AND U4365 ( .A(p_input[8692]), .B(p_input[38692]), .Z(n2909) );
  AND U4366 ( .A(n2911), .B(n2912), .Z(o[8691]) );
  AND U4367 ( .A(p_input[28691]), .B(p_input[18691]), .Z(n2912) );
  AND U4368 ( .A(p_input[8691]), .B(p_input[38691]), .Z(n2911) );
  AND U4369 ( .A(n2913), .B(n2914), .Z(o[8690]) );
  AND U4370 ( .A(p_input[28690]), .B(p_input[18690]), .Z(n2914) );
  AND U4371 ( .A(p_input[8690]), .B(p_input[38690]), .Z(n2913) );
  AND U4372 ( .A(n2915), .B(n2916), .Z(o[868]) );
  AND U4373 ( .A(p_input[20868]), .B(p_input[10868]), .Z(n2916) );
  AND U4374 ( .A(p_input[868]), .B(p_input[30868]), .Z(n2915) );
  AND U4375 ( .A(n2917), .B(n2918), .Z(o[8689]) );
  AND U4376 ( .A(p_input[28689]), .B(p_input[18689]), .Z(n2918) );
  AND U4377 ( .A(p_input[8689]), .B(p_input[38689]), .Z(n2917) );
  AND U4378 ( .A(n2919), .B(n2920), .Z(o[8688]) );
  AND U4379 ( .A(p_input[28688]), .B(p_input[18688]), .Z(n2920) );
  AND U4380 ( .A(p_input[8688]), .B(p_input[38688]), .Z(n2919) );
  AND U4381 ( .A(n2921), .B(n2922), .Z(o[8687]) );
  AND U4382 ( .A(p_input[28687]), .B(p_input[18687]), .Z(n2922) );
  AND U4383 ( .A(p_input[8687]), .B(p_input[38687]), .Z(n2921) );
  AND U4384 ( .A(n2923), .B(n2924), .Z(o[8686]) );
  AND U4385 ( .A(p_input[28686]), .B(p_input[18686]), .Z(n2924) );
  AND U4386 ( .A(p_input[8686]), .B(p_input[38686]), .Z(n2923) );
  AND U4387 ( .A(n2925), .B(n2926), .Z(o[8685]) );
  AND U4388 ( .A(p_input[28685]), .B(p_input[18685]), .Z(n2926) );
  AND U4389 ( .A(p_input[8685]), .B(p_input[38685]), .Z(n2925) );
  AND U4390 ( .A(n2927), .B(n2928), .Z(o[8684]) );
  AND U4391 ( .A(p_input[28684]), .B(p_input[18684]), .Z(n2928) );
  AND U4392 ( .A(p_input[8684]), .B(p_input[38684]), .Z(n2927) );
  AND U4393 ( .A(n2929), .B(n2930), .Z(o[8683]) );
  AND U4394 ( .A(p_input[28683]), .B(p_input[18683]), .Z(n2930) );
  AND U4395 ( .A(p_input[8683]), .B(p_input[38683]), .Z(n2929) );
  AND U4396 ( .A(n2931), .B(n2932), .Z(o[8682]) );
  AND U4397 ( .A(p_input[28682]), .B(p_input[18682]), .Z(n2932) );
  AND U4398 ( .A(p_input[8682]), .B(p_input[38682]), .Z(n2931) );
  AND U4399 ( .A(n2933), .B(n2934), .Z(o[8681]) );
  AND U4400 ( .A(p_input[28681]), .B(p_input[18681]), .Z(n2934) );
  AND U4401 ( .A(p_input[8681]), .B(p_input[38681]), .Z(n2933) );
  AND U4402 ( .A(n2935), .B(n2936), .Z(o[8680]) );
  AND U4403 ( .A(p_input[28680]), .B(p_input[18680]), .Z(n2936) );
  AND U4404 ( .A(p_input[8680]), .B(p_input[38680]), .Z(n2935) );
  AND U4405 ( .A(n2937), .B(n2938), .Z(o[867]) );
  AND U4406 ( .A(p_input[20867]), .B(p_input[10867]), .Z(n2938) );
  AND U4407 ( .A(p_input[867]), .B(p_input[30867]), .Z(n2937) );
  AND U4408 ( .A(n2939), .B(n2940), .Z(o[8679]) );
  AND U4409 ( .A(p_input[28679]), .B(p_input[18679]), .Z(n2940) );
  AND U4410 ( .A(p_input[8679]), .B(p_input[38679]), .Z(n2939) );
  AND U4411 ( .A(n2941), .B(n2942), .Z(o[8678]) );
  AND U4412 ( .A(p_input[28678]), .B(p_input[18678]), .Z(n2942) );
  AND U4413 ( .A(p_input[8678]), .B(p_input[38678]), .Z(n2941) );
  AND U4414 ( .A(n2943), .B(n2944), .Z(o[8677]) );
  AND U4415 ( .A(p_input[28677]), .B(p_input[18677]), .Z(n2944) );
  AND U4416 ( .A(p_input[8677]), .B(p_input[38677]), .Z(n2943) );
  AND U4417 ( .A(n2945), .B(n2946), .Z(o[8676]) );
  AND U4418 ( .A(p_input[28676]), .B(p_input[18676]), .Z(n2946) );
  AND U4419 ( .A(p_input[8676]), .B(p_input[38676]), .Z(n2945) );
  AND U4420 ( .A(n2947), .B(n2948), .Z(o[8675]) );
  AND U4421 ( .A(p_input[28675]), .B(p_input[18675]), .Z(n2948) );
  AND U4422 ( .A(p_input[8675]), .B(p_input[38675]), .Z(n2947) );
  AND U4423 ( .A(n2949), .B(n2950), .Z(o[8674]) );
  AND U4424 ( .A(p_input[28674]), .B(p_input[18674]), .Z(n2950) );
  AND U4425 ( .A(p_input[8674]), .B(p_input[38674]), .Z(n2949) );
  AND U4426 ( .A(n2951), .B(n2952), .Z(o[8673]) );
  AND U4427 ( .A(p_input[28673]), .B(p_input[18673]), .Z(n2952) );
  AND U4428 ( .A(p_input[8673]), .B(p_input[38673]), .Z(n2951) );
  AND U4429 ( .A(n2953), .B(n2954), .Z(o[8672]) );
  AND U4430 ( .A(p_input[28672]), .B(p_input[18672]), .Z(n2954) );
  AND U4431 ( .A(p_input[8672]), .B(p_input[38672]), .Z(n2953) );
  AND U4432 ( .A(n2955), .B(n2956), .Z(o[8671]) );
  AND U4433 ( .A(p_input[28671]), .B(p_input[18671]), .Z(n2956) );
  AND U4434 ( .A(p_input[8671]), .B(p_input[38671]), .Z(n2955) );
  AND U4435 ( .A(n2957), .B(n2958), .Z(o[8670]) );
  AND U4436 ( .A(p_input[28670]), .B(p_input[18670]), .Z(n2958) );
  AND U4437 ( .A(p_input[8670]), .B(p_input[38670]), .Z(n2957) );
  AND U4438 ( .A(n2959), .B(n2960), .Z(o[866]) );
  AND U4439 ( .A(p_input[20866]), .B(p_input[10866]), .Z(n2960) );
  AND U4440 ( .A(p_input[866]), .B(p_input[30866]), .Z(n2959) );
  AND U4441 ( .A(n2961), .B(n2962), .Z(o[8669]) );
  AND U4442 ( .A(p_input[28669]), .B(p_input[18669]), .Z(n2962) );
  AND U4443 ( .A(p_input[8669]), .B(p_input[38669]), .Z(n2961) );
  AND U4444 ( .A(n2963), .B(n2964), .Z(o[8668]) );
  AND U4445 ( .A(p_input[28668]), .B(p_input[18668]), .Z(n2964) );
  AND U4446 ( .A(p_input[8668]), .B(p_input[38668]), .Z(n2963) );
  AND U4447 ( .A(n2965), .B(n2966), .Z(o[8667]) );
  AND U4448 ( .A(p_input[28667]), .B(p_input[18667]), .Z(n2966) );
  AND U4449 ( .A(p_input[8667]), .B(p_input[38667]), .Z(n2965) );
  AND U4450 ( .A(n2967), .B(n2968), .Z(o[8666]) );
  AND U4451 ( .A(p_input[28666]), .B(p_input[18666]), .Z(n2968) );
  AND U4452 ( .A(p_input[8666]), .B(p_input[38666]), .Z(n2967) );
  AND U4453 ( .A(n2969), .B(n2970), .Z(o[8665]) );
  AND U4454 ( .A(p_input[28665]), .B(p_input[18665]), .Z(n2970) );
  AND U4455 ( .A(p_input[8665]), .B(p_input[38665]), .Z(n2969) );
  AND U4456 ( .A(n2971), .B(n2972), .Z(o[8664]) );
  AND U4457 ( .A(p_input[28664]), .B(p_input[18664]), .Z(n2972) );
  AND U4458 ( .A(p_input[8664]), .B(p_input[38664]), .Z(n2971) );
  AND U4459 ( .A(n2973), .B(n2974), .Z(o[8663]) );
  AND U4460 ( .A(p_input[28663]), .B(p_input[18663]), .Z(n2974) );
  AND U4461 ( .A(p_input[8663]), .B(p_input[38663]), .Z(n2973) );
  AND U4462 ( .A(n2975), .B(n2976), .Z(o[8662]) );
  AND U4463 ( .A(p_input[28662]), .B(p_input[18662]), .Z(n2976) );
  AND U4464 ( .A(p_input[8662]), .B(p_input[38662]), .Z(n2975) );
  AND U4465 ( .A(n2977), .B(n2978), .Z(o[8661]) );
  AND U4466 ( .A(p_input[28661]), .B(p_input[18661]), .Z(n2978) );
  AND U4467 ( .A(p_input[8661]), .B(p_input[38661]), .Z(n2977) );
  AND U4468 ( .A(n2979), .B(n2980), .Z(o[8660]) );
  AND U4469 ( .A(p_input[28660]), .B(p_input[18660]), .Z(n2980) );
  AND U4470 ( .A(p_input[8660]), .B(p_input[38660]), .Z(n2979) );
  AND U4471 ( .A(n2981), .B(n2982), .Z(o[865]) );
  AND U4472 ( .A(p_input[20865]), .B(p_input[10865]), .Z(n2982) );
  AND U4473 ( .A(p_input[865]), .B(p_input[30865]), .Z(n2981) );
  AND U4474 ( .A(n2983), .B(n2984), .Z(o[8659]) );
  AND U4475 ( .A(p_input[28659]), .B(p_input[18659]), .Z(n2984) );
  AND U4476 ( .A(p_input[8659]), .B(p_input[38659]), .Z(n2983) );
  AND U4477 ( .A(n2985), .B(n2986), .Z(o[8658]) );
  AND U4478 ( .A(p_input[28658]), .B(p_input[18658]), .Z(n2986) );
  AND U4479 ( .A(p_input[8658]), .B(p_input[38658]), .Z(n2985) );
  AND U4480 ( .A(n2987), .B(n2988), .Z(o[8657]) );
  AND U4481 ( .A(p_input[28657]), .B(p_input[18657]), .Z(n2988) );
  AND U4482 ( .A(p_input[8657]), .B(p_input[38657]), .Z(n2987) );
  AND U4483 ( .A(n2989), .B(n2990), .Z(o[8656]) );
  AND U4484 ( .A(p_input[28656]), .B(p_input[18656]), .Z(n2990) );
  AND U4485 ( .A(p_input[8656]), .B(p_input[38656]), .Z(n2989) );
  AND U4486 ( .A(n2991), .B(n2992), .Z(o[8655]) );
  AND U4487 ( .A(p_input[28655]), .B(p_input[18655]), .Z(n2992) );
  AND U4488 ( .A(p_input[8655]), .B(p_input[38655]), .Z(n2991) );
  AND U4489 ( .A(n2993), .B(n2994), .Z(o[8654]) );
  AND U4490 ( .A(p_input[28654]), .B(p_input[18654]), .Z(n2994) );
  AND U4491 ( .A(p_input[8654]), .B(p_input[38654]), .Z(n2993) );
  AND U4492 ( .A(n2995), .B(n2996), .Z(o[8653]) );
  AND U4493 ( .A(p_input[28653]), .B(p_input[18653]), .Z(n2996) );
  AND U4494 ( .A(p_input[8653]), .B(p_input[38653]), .Z(n2995) );
  AND U4495 ( .A(n2997), .B(n2998), .Z(o[8652]) );
  AND U4496 ( .A(p_input[28652]), .B(p_input[18652]), .Z(n2998) );
  AND U4497 ( .A(p_input[8652]), .B(p_input[38652]), .Z(n2997) );
  AND U4498 ( .A(n2999), .B(n3000), .Z(o[8651]) );
  AND U4499 ( .A(p_input[28651]), .B(p_input[18651]), .Z(n3000) );
  AND U4500 ( .A(p_input[8651]), .B(p_input[38651]), .Z(n2999) );
  AND U4501 ( .A(n3001), .B(n3002), .Z(o[8650]) );
  AND U4502 ( .A(p_input[28650]), .B(p_input[18650]), .Z(n3002) );
  AND U4503 ( .A(p_input[8650]), .B(p_input[38650]), .Z(n3001) );
  AND U4504 ( .A(n3003), .B(n3004), .Z(o[864]) );
  AND U4505 ( .A(p_input[20864]), .B(p_input[10864]), .Z(n3004) );
  AND U4506 ( .A(p_input[864]), .B(p_input[30864]), .Z(n3003) );
  AND U4507 ( .A(n3005), .B(n3006), .Z(o[8649]) );
  AND U4508 ( .A(p_input[28649]), .B(p_input[18649]), .Z(n3006) );
  AND U4509 ( .A(p_input[8649]), .B(p_input[38649]), .Z(n3005) );
  AND U4510 ( .A(n3007), .B(n3008), .Z(o[8648]) );
  AND U4511 ( .A(p_input[28648]), .B(p_input[18648]), .Z(n3008) );
  AND U4512 ( .A(p_input[8648]), .B(p_input[38648]), .Z(n3007) );
  AND U4513 ( .A(n3009), .B(n3010), .Z(o[8647]) );
  AND U4514 ( .A(p_input[28647]), .B(p_input[18647]), .Z(n3010) );
  AND U4515 ( .A(p_input[8647]), .B(p_input[38647]), .Z(n3009) );
  AND U4516 ( .A(n3011), .B(n3012), .Z(o[8646]) );
  AND U4517 ( .A(p_input[28646]), .B(p_input[18646]), .Z(n3012) );
  AND U4518 ( .A(p_input[8646]), .B(p_input[38646]), .Z(n3011) );
  AND U4519 ( .A(n3013), .B(n3014), .Z(o[8645]) );
  AND U4520 ( .A(p_input[28645]), .B(p_input[18645]), .Z(n3014) );
  AND U4521 ( .A(p_input[8645]), .B(p_input[38645]), .Z(n3013) );
  AND U4522 ( .A(n3015), .B(n3016), .Z(o[8644]) );
  AND U4523 ( .A(p_input[28644]), .B(p_input[18644]), .Z(n3016) );
  AND U4524 ( .A(p_input[8644]), .B(p_input[38644]), .Z(n3015) );
  AND U4525 ( .A(n3017), .B(n3018), .Z(o[8643]) );
  AND U4526 ( .A(p_input[28643]), .B(p_input[18643]), .Z(n3018) );
  AND U4527 ( .A(p_input[8643]), .B(p_input[38643]), .Z(n3017) );
  AND U4528 ( .A(n3019), .B(n3020), .Z(o[8642]) );
  AND U4529 ( .A(p_input[28642]), .B(p_input[18642]), .Z(n3020) );
  AND U4530 ( .A(p_input[8642]), .B(p_input[38642]), .Z(n3019) );
  AND U4531 ( .A(n3021), .B(n3022), .Z(o[8641]) );
  AND U4532 ( .A(p_input[28641]), .B(p_input[18641]), .Z(n3022) );
  AND U4533 ( .A(p_input[8641]), .B(p_input[38641]), .Z(n3021) );
  AND U4534 ( .A(n3023), .B(n3024), .Z(o[8640]) );
  AND U4535 ( .A(p_input[28640]), .B(p_input[18640]), .Z(n3024) );
  AND U4536 ( .A(p_input[8640]), .B(p_input[38640]), .Z(n3023) );
  AND U4537 ( .A(n3025), .B(n3026), .Z(o[863]) );
  AND U4538 ( .A(p_input[20863]), .B(p_input[10863]), .Z(n3026) );
  AND U4539 ( .A(p_input[863]), .B(p_input[30863]), .Z(n3025) );
  AND U4540 ( .A(n3027), .B(n3028), .Z(o[8639]) );
  AND U4541 ( .A(p_input[28639]), .B(p_input[18639]), .Z(n3028) );
  AND U4542 ( .A(p_input[8639]), .B(p_input[38639]), .Z(n3027) );
  AND U4543 ( .A(n3029), .B(n3030), .Z(o[8638]) );
  AND U4544 ( .A(p_input[28638]), .B(p_input[18638]), .Z(n3030) );
  AND U4545 ( .A(p_input[8638]), .B(p_input[38638]), .Z(n3029) );
  AND U4546 ( .A(n3031), .B(n3032), .Z(o[8637]) );
  AND U4547 ( .A(p_input[28637]), .B(p_input[18637]), .Z(n3032) );
  AND U4548 ( .A(p_input[8637]), .B(p_input[38637]), .Z(n3031) );
  AND U4549 ( .A(n3033), .B(n3034), .Z(o[8636]) );
  AND U4550 ( .A(p_input[28636]), .B(p_input[18636]), .Z(n3034) );
  AND U4551 ( .A(p_input[8636]), .B(p_input[38636]), .Z(n3033) );
  AND U4552 ( .A(n3035), .B(n3036), .Z(o[8635]) );
  AND U4553 ( .A(p_input[28635]), .B(p_input[18635]), .Z(n3036) );
  AND U4554 ( .A(p_input[8635]), .B(p_input[38635]), .Z(n3035) );
  AND U4555 ( .A(n3037), .B(n3038), .Z(o[8634]) );
  AND U4556 ( .A(p_input[28634]), .B(p_input[18634]), .Z(n3038) );
  AND U4557 ( .A(p_input[8634]), .B(p_input[38634]), .Z(n3037) );
  AND U4558 ( .A(n3039), .B(n3040), .Z(o[8633]) );
  AND U4559 ( .A(p_input[28633]), .B(p_input[18633]), .Z(n3040) );
  AND U4560 ( .A(p_input[8633]), .B(p_input[38633]), .Z(n3039) );
  AND U4561 ( .A(n3041), .B(n3042), .Z(o[8632]) );
  AND U4562 ( .A(p_input[28632]), .B(p_input[18632]), .Z(n3042) );
  AND U4563 ( .A(p_input[8632]), .B(p_input[38632]), .Z(n3041) );
  AND U4564 ( .A(n3043), .B(n3044), .Z(o[8631]) );
  AND U4565 ( .A(p_input[28631]), .B(p_input[18631]), .Z(n3044) );
  AND U4566 ( .A(p_input[8631]), .B(p_input[38631]), .Z(n3043) );
  AND U4567 ( .A(n3045), .B(n3046), .Z(o[8630]) );
  AND U4568 ( .A(p_input[28630]), .B(p_input[18630]), .Z(n3046) );
  AND U4569 ( .A(p_input[8630]), .B(p_input[38630]), .Z(n3045) );
  AND U4570 ( .A(n3047), .B(n3048), .Z(o[862]) );
  AND U4571 ( .A(p_input[20862]), .B(p_input[10862]), .Z(n3048) );
  AND U4572 ( .A(p_input[862]), .B(p_input[30862]), .Z(n3047) );
  AND U4573 ( .A(n3049), .B(n3050), .Z(o[8629]) );
  AND U4574 ( .A(p_input[28629]), .B(p_input[18629]), .Z(n3050) );
  AND U4575 ( .A(p_input[8629]), .B(p_input[38629]), .Z(n3049) );
  AND U4576 ( .A(n3051), .B(n3052), .Z(o[8628]) );
  AND U4577 ( .A(p_input[28628]), .B(p_input[18628]), .Z(n3052) );
  AND U4578 ( .A(p_input[8628]), .B(p_input[38628]), .Z(n3051) );
  AND U4579 ( .A(n3053), .B(n3054), .Z(o[8627]) );
  AND U4580 ( .A(p_input[28627]), .B(p_input[18627]), .Z(n3054) );
  AND U4581 ( .A(p_input[8627]), .B(p_input[38627]), .Z(n3053) );
  AND U4582 ( .A(n3055), .B(n3056), .Z(o[8626]) );
  AND U4583 ( .A(p_input[28626]), .B(p_input[18626]), .Z(n3056) );
  AND U4584 ( .A(p_input[8626]), .B(p_input[38626]), .Z(n3055) );
  AND U4585 ( .A(n3057), .B(n3058), .Z(o[8625]) );
  AND U4586 ( .A(p_input[28625]), .B(p_input[18625]), .Z(n3058) );
  AND U4587 ( .A(p_input[8625]), .B(p_input[38625]), .Z(n3057) );
  AND U4588 ( .A(n3059), .B(n3060), .Z(o[8624]) );
  AND U4589 ( .A(p_input[28624]), .B(p_input[18624]), .Z(n3060) );
  AND U4590 ( .A(p_input[8624]), .B(p_input[38624]), .Z(n3059) );
  AND U4591 ( .A(n3061), .B(n3062), .Z(o[8623]) );
  AND U4592 ( .A(p_input[28623]), .B(p_input[18623]), .Z(n3062) );
  AND U4593 ( .A(p_input[8623]), .B(p_input[38623]), .Z(n3061) );
  AND U4594 ( .A(n3063), .B(n3064), .Z(o[8622]) );
  AND U4595 ( .A(p_input[28622]), .B(p_input[18622]), .Z(n3064) );
  AND U4596 ( .A(p_input[8622]), .B(p_input[38622]), .Z(n3063) );
  AND U4597 ( .A(n3065), .B(n3066), .Z(o[8621]) );
  AND U4598 ( .A(p_input[28621]), .B(p_input[18621]), .Z(n3066) );
  AND U4599 ( .A(p_input[8621]), .B(p_input[38621]), .Z(n3065) );
  AND U4600 ( .A(n3067), .B(n3068), .Z(o[8620]) );
  AND U4601 ( .A(p_input[28620]), .B(p_input[18620]), .Z(n3068) );
  AND U4602 ( .A(p_input[8620]), .B(p_input[38620]), .Z(n3067) );
  AND U4603 ( .A(n3069), .B(n3070), .Z(o[861]) );
  AND U4604 ( .A(p_input[20861]), .B(p_input[10861]), .Z(n3070) );
  AND U4605 ( .A(p_input[861]), .B(p_input[30861]), .Z(n3069) );
  AND U4606 ( .A(n3071), .B(n3072), .Z(o[8619]) );
  AND U4607 ( .A(p_input[28619]), .B(p_input[18619]), .Z(n3072) );
  AND U4608 ( .A(p_input[8619]), .B(p_input[38619]), .Z(n3071) );
  AND U4609 ( .A(n3073), .B(n3074), .Z(o[8618]) );
  AND U4610 ( .A(p_input[28618]), .B(p_input[18618]), .Z(n3074) );
  AND U4611 ( .A(p_input[8618]), .B(p_input[38618]), .Z(n3073) );
  AND U4612 ( .A(n3075), .B(n3076), .Z(o[8617]) );
  AND U4613 ( .A(p_input[28617]), .B(p_input[18617]), .Z(n3076) );
  AND U4614 ( .A(p_input[8617]), .B(p_input[38617]), .Z(n3075) );
  AND U4615 ( .A(n3077), .B(n3078), .Z(o[8616]) );
  AND U4616 ( .A(p_input[28616]), .B(p_input[18616]), .Z(n3078) );
  AND U4617 ( .A(p_input[8616]), .B(p_input[38616]), .Z(n3077) );
  AND U4618 ( .A(n3079), .B(n3080), .Z(o[8615]) );
  AND U4619 ( .A(p_input[28615]), .B(p_input[18615]), .Z(n3080) );
  AND U4620 ( .A(p_input[8615]), .B(p_input[38615]), .Z(n3079) );
  AND U4621 ( .A(n3081), .B(n3082), .Z(o[8614]) );
  AND U4622 ( .A(p_input[28614]), .B(p_input[18614]), .Z(n3082) );
  AND U4623 ( .A(p_input[8614]), .B(p_input[38614]), .Z(n3081) );
  AND U4624 ( .A(n3083), .B(n3084), .Z(o[8613]) );
  AND U4625 ( .A(p_input[28613]), .B(p_input[18613]), .Z(n3084) );
  AND U4626 ( .A(p_input[8613]), .B(p_input[38613]), .Z(n3083) );
  AND U4627 ( .A(n3085), .B(n3086), .Z(o[8612]) );
  AND U4628 ( .A(p_input[28612]), .B(p_input[18612]), .Z(n3086) );
  AND U4629 ( .A(p_input[8612]), .B(p_input[38612]), .Z(n3085) );
  AND U4630 ( .A(n3087), .B(n3088), .Z(o[8611]) );
  AND U4631 ( .A(p_input[28611]), .B(p_input[18611]), .Z(n3088) );
  AND U4632 ( .A(p_input[8611]), .B(p_input[38611]), .Z(n3087) );
  AND U4633 ( .A(n3089), .B(n3090), .Z(o[8610]) );
  AND U4634 ( .A(p_input[28610]), .B(p_input[18610]), .Z(n3090) );
  AND U4635 ( .A(p_input[8610]), .B(p_input[38610]), .Z(n3089) );
  AND U4636 ( .A(n3091), .B(n3092), .Z(o[860]) );
  AND U4637 ( .A(p_input[20860]), .B(p_input[10860]), .Z(n3092) );
  AND U4638 ( .A(p_input[860]), .B(p_input[30860]), .Z(n3091) );
  AND U4639 ( .A(n3093), .B(n3094), .Z(o[8609]) );
  AND U4640 ( .A(p_input[28609]), .B(p_input[18609]), .Z(n3094) );
  AND U4641 ( .A(p_input[8609]), .B(p_input[38609]), .Z(n3093) );
  AND U4642 ( .A(n3095), .B(n3096), .Z(o[8608]) );
  AND U4643 ( .A(p_input[28608]), .B(p_input[18608]), .Z(n3096) );
  AND U4644 ( .A(p_input[8608]), .B(p_input[38608]), .Z(n3095) );
  AND U4645 ( .A(n3097), .B(n3098), .Z(o[8607]) );
  AND U4646 ( .A(p_input[28607]), .B(p_input[18607]), .Z(n3098) );
  AND U4647 ( .A(p_input[8607]), .B(p_input[38607]), .Z(n3097) );
  AND U4648 ( .A(n3099), .B(n3100), .Z(o[8606]) );
  AND U4649 ( .A(p_input[28606]), .B(p_input[18606]), .Z(n3100) );
  AND U4650 ( .A(p_input[8606]), .B(p_input[38606]), .Z(n3099) );
  AND U4651 ( .A(n3101), .B(n3102), .Z(o[8605]) );
  AND U4652 ( .A(p_input[28605]), .B(p_input[18605]), .Z(n3102) );
  AND U4653 ( .A(p_input[8605]), .B(p_input[38605]), .Z(n3101) );
  AND U4654 ( .A(n3103), .B(n3104), .Z(o[8604]) );
  AND U4655 ( .A(p_input[28604]), .B(p_input[18604]), .Z(n3104) );
  AND U4656 ( .A(p_input[8604]), .B(p_input[38604]), .Z(n3103) );
  AND U4657 ( .A(n3105), .B(n3106), .Z(o[8603]) );
  AND U4658 ( .A(p_input[28603]), .B(p_input[18603]), .Z(n3106) );
  AND U4659 ( .A(p_input[8603]), .B(p_input[38603]), .Z(n3105) );
  AND U4660 ( .A(n3107), .B(n3108), .Z(o[8602]) );
  AND U4661 ( .A(p_input[28602]), .B(p_input[18602]), .Z(n3108) );
  AND U4662 ( .A(p_input[8602]), .B(p_input[38602]), .Z(n3107) );
  AND U4663 ( .A(n3109), .B(n3110), .Z(o[8601]) );
  AND U4664 ( .A(p_input[28601]), .B(p_input[18601]), .Z(n3110) );
  AND U4665 ( .A(p_input[8601]), .B(p_input[38601]), .Z(n3109) );
  AND U4666 ( .A(n3111), .B(n3112), .Z(o[8600]) );
  AND U4667 ( .A(p_input[28600]), .B(p_input[18600]), .Z(n3112) );
  AND U4668 ( .A(p_input[8600]), .B(p_input[38600]), .Z(n3111) );
  AND U4669 ( .A(n3113), .B(n3114), .Z(o[85]) );
  AND U4670 ( .A(p_input[20085]), .B(p_input[10085]), .Z(n3114) );
  AND U4671 ( .A(p_input[85]), .B(p_input[30085]), .Z(n3113) );
  AND U4672 ( .A(n3115), .B(n3116), .Z(o[859]) );
  AND U4673 ( .A(p_input[20859]), .B(p_input[10859]), .Z(n3116) );
  AND U4674 ( .A(p_input[859]), .B(p_input[30859]), .Z(n3115) );
  AND U4675 ( .A(n3117), .B(n3118), .Z(o[8599]) );
  AND U4676 ( .A(p_input[28599]), .B(p_input[18599]), .Z(n3118) );
  AND U4677 ( .A(p_input[8599]), .B(p_input[38599]), .Z(n3117) );
  AND U4678 ( .A(n3119), .B(n3120), .Z(o[8598]) );
  AND U4679 ( .A(p_input[28598]), .B(p_input[18598]), .Z(n3120) );
  AND U4680 ( .A(p_input[8598]), .B(p_input[38598]), .Z(n3119) );
  AND U4681 ( .A(n3121), .B(n3122), .Z(o[8597]) );
  AND U4682 ( .A(p_input[28597]), .B(p_input[18597]), .Z(n3122) );
  AND U4683 ( .A(p_input[8597]), .B(p_input[38597]), .Z(n3121) );
  AND U4684 ( .A(n3123), .B(n3124), .Z(o[8596]) );
  AND U4685 ( .A(p_input[28596]), .B(p_input[18596]), .Z(n3124) );
  AND U4686 ( .A(p_input[8596]), .B(p_input[38596]), .Z(n3123) );
  AND U4687 ( .A(n3125), .B(n3126), .Z(o[8595]) );
  AND U4688 ( .A(p_input[28595]), .B(p_input[18595]), .Z(n3126) );
  AND U4689 ( .A(p_input[8595]), .B(p_input[38595]), .Z(n3125) );
  AND U4690 ( .A(n3127), .B(n3128), .Z(o[8594]) );
  AND U4691 ( .A(p_input[28594]), .B(p_input[18594]), .Z(n3128) );
  AND U4692 ( .A(p_input[8594]), .B(p_input[38594]), .Z(n3127) );
  AND U4693 ( .A(n3129), .B(n3130), .Z(o[8593]) );
  AND U4694 ( .A(p_input[28593]), .B(p_input[18593]), .Z(n3130) );
  AND U4695 ( .A(p_input[8593]), .B(p_input[38593]), .Z(n3129) );
  AND U4696 ( .A(n3131), .B(n3132), .Z(o[8592]) );
  AND U4697 ( .A(p_input[28592]), .B(p_input[18592]), .Z(n3132) );
  AND U4698 ( .A(p_input[8592]), .B(p_input[38592]), .Z(n3131) );
  AND U4699 ( .A(n3133), .B(n3134), .Z(o[8591]) );
  AND U4700 ( .A(p_input[28591]), .B(p_input[18591]), .Z(n3134) );
  AND U4701 ( .A(p_input[8591]), .B(p_input[38591]), .Z(n3133) );
  AND U4702 ( .A(n3135), .B(n3136), .Z(o[8590]) );
  AND U4703 ( .A(p_input[28590]), .B(p_input[18590]), .Z(n3136) );
  AND U4704 ( .A(p_input[8590]), .B(p_input[38590]), .Z(n3135) );
  AND U4705 ( .A(n3137), .B(n3138), .Z(o[858]) );
  AND U4706 ( .A(p_input[20858]), .B(p_input[10858]), .Z(n3138) );
  AND U4707 ( .A(p_input[858]), .B(p_input[30858]), .Z(n3137) );
  AND U4708 ( .A(n3139), .B(n3140), .Z(o[8589]) );
  AND U4709 ( .A(p_input[28589]), .B(p_input[18589]), .Z(n3140) );
  AND U4710 ( .A(p_input[8589]), .B(p_input[38589]), .Z(n3139) );
  AND U4711 ( .A(n3141), .B(n3142), .Z(o[8588]) );
  AND U4712 ( .A(p_input[28588]), .B(p_input[18588]), .Z(n3142) );
  AND U4713 ( .A(p_input[8588]), .B(p_input[38588]), .Z(n3141) );
  AND U4714 ( .A(n3143), .B(n3144), .Z(o[8587]) );
  AND U4715 ( .A(p_input[28587]), .B(p_input[18587]), .Z(n3144) );
  AND U4716 ( .A(p_input[8587]), .B(p_input[38587]), .Z(n3143) );
  AND U4717 ( .A(n3145), .B(n3146), .Z(o[8586]) );
  AND U4718 ( .A(p_input[28586]), .B(p_input[18586]), .Z(n3146) );
  AND U4719 ( .A(p_input[8586]), .B(p_input[38586]), .Z(n3145) );
  AND U4720 ( .A(n3147), .B(n3148), .Z(o[8585]) );
  AND U4721 ( .A(p_input[28585]), .B(p_input[18585]), .Z(n3148) );
  AND U4722 ( .A(p_input[8585]), .B(p_input[38585]), .Z(n3147) );
  AND U4723 ( .A(n3149), .B(n3150), .Z(o[8584]) );
  AND U4724 ( .A(p_input[28584]), .B(p_input[18584]), .Z(n3150) );
  AND U4725 ( .A(p_input[8584]), .B(p_input[38584]), .Z(n3149) );
  AND U4726 ( .A(n3151), .B(n3152), .Z(o[8583]) );
  AND U4727 ( .A(p_input[28583]), .B(p_input[18583]), .Z(n3152) );
  AND U4728 ( .A(p_input[8583]), .B(p_input[38583]), .Z(n3151) );
  AND U4729 ( .A(n3153), .B(n3154), .Z(o[8582]) );
  AND U4730 ( .A(p_input[28582]), .B(p_input[18582]), .Z(n3154) );
  AND U4731 ( .A(p_input[8582]), .B(p_input[38582]), .Z(n3153) );
  AND U4732 ( .A(n3155), .B(n3156), .Z(o[8581]) );
  AND U4733 ( .A(p_input[28581]), .B(p_input[18581]), .Z(n3156) );
  AND U4734 ( .A(p_input[8581]), .B(p_input[38581]), .Z(n3155) );
  AND U4735 ( .A(n3157), .B(n3158), .Z(o[8580]) );
  AND U4736 ( .A(p_input[28580]), .B(p_input[18580]), .Z(n3158) );
  AND U4737 ( .A(p_input[8580]), .B(p_input[38580]), .Z(n3157) );
  AND U4738 ( .A(n3159), .B(n3160), .Z(o[857]) );
  AND U4739 ( .A(p_input[20857]), .B(p_input[10857]), .Z(n3160) );
  AND U4740 ( .A(p_input[857]), .B(p_input[30857]), .Z(n3159) );
  AND U4741 ( .A(n3161), .B(n3162), .Z(o[8579]) );
  AND U4742 ( .A(p_input[28579]), .B(p_input[18579]), .Z(n3162) );
  AND U4743 ( .A(p_input[8579]), .B(p_input[38579]), .Z(n3161) );
  AND U4744 ( .A(n3163), .B(n3164), .Z(o[8578]) );
  AND U4745 ( .A(p_input[28578]), .B(p_input[18578]), .Z(n3164) );
  AND U4746 ( .A(p_input[8578]), .B(p_input[38578]), .Z(n3163) );
  AND U4747 ( .A(n3165), .B(n3166), .Z(o[8577]) );
  AND U4748 ( .A(p_input[28577]), .B(p_input[18577]), .Z(n3166) );
  AND U4749 ( .A(p_input[8577]), .B(p_input[38577]), .Z(n3165) );
  AND U4750 ( .A(n3167), .B(n3168), .Z(o[8576]) );
  AND U4751 ( .A(p_input[28576]), .B(p_input[18576]), .Z(n3168) );
  AND U4752 ( .A(p_input[8576]), .B(p_input[38576]), .Z(n3167) );
  AND U4753 ( .A(n3169), .B(n3170), .Z(o[8575]) );
  AND U4754 ( .A(p_input[28575]), .B(p_input[18575]), .Z(n3170) );
  AND U4755 ( .A(p_input[8575]), .B(p_input[38575]), .Z(n3169) );
  AND U4756 ( .A(n3171), .B(n3172), .Z(o[8574]) );
  AND U4757 ( .A(p_input[28574]), .B(p_input[18574]), .Z(n3172) );
  AND U4758 ( .A(p_input[8574]), .B(p_input[38574]), .Z(n3171) );
  AND U4759 ( .A(n3173), .B(n3174), .Z(o[8573]) );
  AND U4760 ( .A(p_input[28573]), .B(p_input[18573]), .Z(n3174) );
  AND U4761 ( .A(p_input[8573]), .B(p_input[38573]), .Z(n3173) );
  AND U4762 ( .A(n3175), .B(n3176), .Z(o[8572]) );
  AND U4763 ( .A(p_input[28572]), .B(p_input[18572]), .Z(n3176) );
  AND U4764 ( .A(p_input[8572]), .B(p_input[38572]), .Z(n3175) );
  AND U4765 ( .A(n3177), .B(n3178), .Z(o[8571]) );
  AND U4766 ( .A(p_input[28571]), .B(p_input[18571]), .Z(n3178) );
  AND U4767 ( .A(p_input[8571]), .B(p_input[38571]), .Z(n3177) );
  AND U4768 ( .A(n3179), .B(n3180), .Z(o[8570]) );
  AND U4769 ( .A(p_input[28570]), .B(p_input[18570]), .Z(n3180) );
  AND U4770 ( .A(p_input[8570]), .B(p_input[38570]), .Z(n3179) );
  AND U4771 ( .A(n3181), .B(n3182), .Z(o[856]) );
  AND U4772 ( .A(p_input[20856]), .B(p_input[10856]), .Z(n3182) );
  AND U4773 ( .A(p_input[856]), .B(p_input[30856]), .Z(n3181) );
  AND U4774 ( .A(n3183), .B(n3184), .Z(o[8569]) );
  AND U4775 ( .A(p_input[28569]), .B(p_input[18569]), .Z(n3184) );
  AND U4776 ( .A(p_input[8569]), .B(p_input[38569]), .Z(n3183) );
  AND U4777 ( .A(n3185), .B(n3186), .Z(o[8568]) );
  AND U4778 ( .A(p_input[28568]), .B(p_input[18568]), .Z(n3186) );
  AND U4779 ( .A(p_input[8568]), .B(p_input[38568]), .Z(n3185) );
  AND U4780 ( .A(n3187), .B(n3188), .Z(o[8567]) );
  AND U4781 ( .A(p_input[28567]), .B(p_input[18567]), .Z(n3188) );
  AND U4782 ( .A(p_input[8567]), .B(p_input[38567]), .Z(n3187) );
  AND U4783 ( .A(n3189), .B(n3190), .Z(o[8566]) );
  AND U4784 ( .A(p_input[28566]), .B(p_input[18566]), .Z(n3190) );
  AND U4785 ( .A(p_input[8566]), .B(p_input[38566]), .Z(n3189) );
  AND U4786 ( .A(n3191), .B(n3192), .Z(o[8565]) );
  AND U4787 ( .A(p_input[28565]), .B(p_input[18565]), .Z(n3192) );
  AND U4788 ( .A(p_input[8565]), .B(p_input[38565]), .Z(n3191) );
  AND U4789 ( .A(n3193), .B(n3194), .Z(o[8564]) );
  AND U4790 ( .A(p_input[28564]), .B(p_input[18564]), .Z(n3194) );
  AND U4791 ( .A(p_input[8564]), .B(p_input[38564]), .Z(n3193) );
  AND U4792 ( .A(n3195), .B(n3196), .Z(o[8563]) );
  AND U4793 ( .A(p_input[28563]), .B(p_input[18563]), .Z(n3196) );
  AND U4794 ( .A(p_input[8563]), .B(p_input[38563]), .Z(n3195) );
  AND U4795 ( .A(n3197), .B(n3198), .Z(o[8562]) );
  AND U4796 ( .A(p_input[28562]), .B(p_input[18562]), .Z(n3198) );
  AND U4797 ( .A(p_input[8562]), .B(p_input[38562]), .Z(n3197) );
  AND U4798 ( .A(n3199), .B(n3200), .Z(o[8561]) );
  AND U4799 ( .A(p_input[28561]), .B(p_input[18561]), .Z(n3200) );
  AND U4800 ( .A(p_input[8561]), .B(p_input[38561]), .Z(n3199) );
  AND U4801 ( .A(n3201), .B(n3202), .Z(o[8560]) );
  AND U4802 ( .A(p_input[28560]), .B(p_input[18560]), .Z(n3202) );
  AND U4803 ( .A(p_input[8560]), .B(p_input[38560]), .Z(n3201) );
  AND U4804 ( .A(n3203), .B(n3204), .Z(o[855]) );
  AND U4805 ( .A(p_input[20855]), .B(p_input[10855]), .Z(n3204) );
  AND U4806 ( .A(p_input[855]), .B(p_input[30855]), .Z(n3203) );
  AND U4807 ( .A(n3205), .B(n3206), .Z(o[8559]) );
  AND U4808 ( .A(p_input[28559]), .B(p_input[18559]), .Z(n3206) );
  AND U4809 ( .A(p_input[8559]), .B(p_input[38559]), .Z(n3205) );
  AND U4810 ( .A(n3207), .B(n3208), .Z(o[8558]) );
  AND U4811 ( .A(p_input[28558]), .B(p_input[18558]), .Z(n3208) );
  AND U4812 ( .A(p_input[8558]), .B(p_input[38558]), .Z(n3207) );
  AND U4813 ( .A(n3209), .B(n3210), .Z(o[8557]) );
  AND U4814 ( .A(p_input[28557]), .B(p_input[18557]), .Z(n3210) );
  AND U4815 ( .A(p_input[8557]), .B(p_input[38557]), .Z(n3209) );
  AND U4816 ( .A(n3211), .B(n3212), .Z(o[8556]) );
  AND U4817 ( .A(p_input[28556]), .B(p_input[18556]), .Z(n3212) );
  AND U4818 ( .A(p_input[8556]), .B(p_input[38556]), .Z(n3211) );
  AND U4819 ( .A(n3213), .B(n3214), .Z(o[8555]) );
  AND U4820 ( .A(p_input[28555]), .B(p_input[18555]), .Z(n3214) );
  AND U4821 ( .A(p_input[8555]), .B(p_input[38555]), .Z(n3213) );
  AND U4822 ( .A(n3215), .B(n3216), .Z(o[8554]) );
  AND U4823 ( .A(p_input[28554]), .B(p_input[18554]), .Z(n3216) );
  AND U4824 ( .A(p_input[8554]), .B(p_input[38554]), .Z(n3215) );
  AND U4825 ( .A(n3217), .B(n3218), .Z(o[8553]) );
  AND U4826 ( .A(p_input[28553]), .B(p_input[18553]), .Z(n3218) );
  AND U4827 ( .A(p_input[8553]), .B(p_input[38553]), .Z(n3217) );
  AND U4828 ( .A(n3219), .B(n3220), .Z(o[8552]) );
  AND U4829 ( .A(p_input[28552]), .B(p_input[18552]), .Z(n3220) );
  AND U4830 ( .A(p_input[8552]), .B(p_input[38552]), .Z(n3219) );
  AND U4831 ( .A(n3221), .B(n3222), .Z(o[8551]) );
  AND U4832 ( .A(p_input[28551]), .B(p_input[18551]), .Z(n3222) );
  AND U4833 ( .A(p_input[8551]), .B(p_input[38551]), .Z(n3221) );
  AND U4834 ( .A(n3223), .B(n3224), .Z(o[8550]) );
  AND U4835 ( .A(p_input[28550]), .B(p_input[18550]), .Z(n3224) );
  AND U4836 ( .A(p_input[8550]), .B(p_input[38550]), .Z(n3223) );
  AND U4837 ( .A(n3225), .B(n3226), .Z(o[854]) );
  AND U4838 ( .A(p_input[20854]), .B(p_input[10854]), .Z(n3226) );
  AND U4839 ( .A(p_input[854]), .B(p_input[30854]), .Z(n3225) );
  AND U4840 ( .A(n3227), .B(n3228), .Z(o[8549]) );
  AND U4841 ( .A(p_input[28549]), .B(p_input[18549]), .Z(n3228) );
  AND U4842 ( .A(p_input[8549]), .B(p_input[38549]), .Z(n3227) );
  AND U4843 ( .A(n3229), .B(n3230), .Z(o[8548]) );
  AND U4844 ( .A(p_input[28548]), .B(p_input[18548]), .Z(n3230) );
  AND U4845 ( .A(p_input[8548]), .B(p_input[38548]), .Z(n3229) );
  AND U4846 ( .A(n3231), .B(n3232), .Z(o[8547]) );
  AND U4847 ( .A(p_input[28547]), .B(p_input[18547]), .Z(n3232) );
  AND U4848 ( .A(p_input[8547]), .B(p_input[38547]), .Z(n3231) );
  AND U4849 ( .A(n3233), .B(n3234), .Z(o[8546]) );
  AND U4850 ( .A(p_input[28546]), .B(p_input[18546]), .Z(n3234) );
  AND U4851 ( .A(p_input[8546]), .B(p_input[38546]), .Z(n3233) );
  AND U4852 ( .A(n3235), .B(n3236), .Z(o[8545]) );
  AND U4853 ( .A(p_input[28545]), .B(p_input[18545]), .Z(n3236) );
  AND U4854 ( .A(p_input[8545]), .B(p_input[38545]), .Z(n3235) );
  AND U4855 ( .A(n3237), .B(n3238), .Z(o[8544]) );
  AND U4856 ( .A(p_input[28544]), .B(p_input[18544]), .Z(n3238) );
  AND U4857 ( .A(p_input[8544]), .B(p_input[38544]), .Z(n3237) );
  AND U4858 ( .A(n3239), .B(n3240), .Z(o[8543]) );
  AND U4859 ( .A(p_input[28543]), .B(p_input[18543]), .Z(n3240) );
  AND U4860 ( .A(p_input[8543]), .B(p_input[38543]), .Z(n3239) );
  AND U4861 ( .A(n3241), .B(n3242), .Z(o[8542]) );
  AND U4862 ( .A(p_input[28542]), .B(p_input[18542]), .Z(n3242) );
  AND U4863 ( .A(p_input[8542]), .B(p_input[38542]), .Z(n3241) );
  AND U4864 ( .A(n3243), .B(n3244), .Z(o[8541]) );
  AND U4865 ( .A(p_input[28541]), .B(p_input[18541]), .Z(n3244) );
  AND U4866 ( .A(p_input[8541]), .B(p_input[38541]), .Z(n3243) );
  AND U4867 ( .A(n3245), .B(n3246), .Z(o[8540]) );
  AND U4868 ( .A(p_input[28540]), .B(p_input[18540]), .Z(n3246) );
  AND U4869 ( .A(p_input[8540]), .B(p_input[38540]), .Z(n3245) );
  AND U4870 ( .A(n3247), .B(n3248), .Z(o[853]) );
  AND U4871 ( .A(p_input[20853]), .B(p_input[10853]), .Z(n3248) );
  AND U4872 ( .A(p_input[853]), .B(p_input[30853]), .Z(n3247) );
  AND U4873 ( .A(n3249), .B(n3250), .Z(o[8539]) );
  AND U4874 ( .A(p_input[28539]), .B(p_input[18539]), .Z(n3250) );
  AND U4875 ( .A(p_input[8539]), .B(p_input[38539]), .Z(n3249) );
  AND U4876 ( .A(n3251), .B(n3252), .Z(o[8538]) );
  AND U4877 ( .A(p_input[28538]), .B(p_input[18538]), .Z(n3252) );
  AND U4878 ( .A(p_input[8538]), .B(p_input[38538]), .Z(n3251) );
  AND U4879 ( .A(n3253), .B(n3254), .Z(o[8537]) );
  AND U4880 ( .A(p_input[28537]), .B(p_input[18537]), .Z(n3254) );
  AND U4881 ( .A(p_input[8537]), .B(p_input[38537]), .Z(n3253) );
  AND U4882 ( .A(n3255), .B(n3256), .Z(o[8536]) );
  AND U4883 ( .A(p_input[28536]), .B(p_input[18536]), .Z(n3256) );
  AND U4884 ( .A(p_input[8536]), .B(p_input[38536]), .Z(n3255) );
  AND U4885 ( .A(n3257), .B(n3258), .Z(o[8535]) );
  AND U4886 ( .A(p_input[28535]), .B(p_input[18535]), .Z(n3258) );
  AND U4887 ( .A(p_input[8535]), .B(p_input[38535]), .Z(n3257) );
  AND U4888 ( .A(n3259), .B(n3260), .Z(o[8534]) );
  AND U4889 ( .A(p_input[28534]), .B(p_input[18534]), .Z(n3260) );
  AND U4890 ( .A(p_input[8534]), .B(p_input[38534]), .Z(n3259) );
  AND U4891 ( .A(n3261), .B(n3262), .Z(o[8533]) );
  AND U4892 ( .A(p_input[28533]), .B(p_input[18533]), .Z(n3262) );
  AND U4893 ( .A(p_input[8533]), .B(p_input[38533]), .Z(n3261) );
  AND U4894 ( .A(n3263), .B(n3264), .Z(o[8532]) );
  AND U4895 ( .A(p_input[28532]), .B(p_input[18532]), .Z(n3264) );
  AND U4896 ( .A(p_input[8532]), .B(p_input[38532]), .Z(n3263) );
  AND U4897 ( .A(n3265), .B(n3266), .Z(o[8531]) );
  AND U4898 ( .A(p_input[28531]), .B(p_input[18531]), .Z(n3266) );
  AND U4899 ( .A(p_input[8531]), .B(p_input[38531]), .Z(n3265) );
  AND U4900 ( .A(n3267), .B(n3268), .Z(o[8530]) );
  AND U4901 ( .A(p_input[28530]), .B(p_input[18530]), .Z(n3268) );
  AND U4902 ( .A(p_input[8530]), .B(p_input[38530]), .Z(n3267) );
  AND U4903 ( .A(n3269), .B(n3270), .Z(o[852]) );
  AND U4904 ( .A(p_input[20852]), .B(p_input[10852]), .Z(n3270) );
  AND U4905 ( .A(p_input[852]), .B(p_input[30852]), .Z(n3269) );
  AND U4906 ( .A(n3271), .B(n3272), .Z(o[8529]) );
  AND U4907 ( .A(p_input[28529]), .B(p_input[18529]), .Z(n3272) );
  AND U4908 ( .A(p_input[8529]), .B(p_input[38529]), .Z(n3271) );
  AND U4909 ( .A(n3273), .B(n3274), .Z(o[8528]) );
  AND U4910 ( .A(p_input[28528]), .B(p_input[18528]), .Z(n3274) );
  AND U4911 ( .A(p_input[8528]), .B(p_input[38528]), .Z(n3273) );
  AND U4912 ( .A(n3275), .B(n3276), .Z(o[8527]) );
  AND U4913 ( .A(p_input[28527]), .B(p_input[18527]), .Z(n3276) );
  AND U4914 ( .A(p_input[8527]), .B(p_input[38527]), .Z(n3275) );
  AND U4915 ( .A(n3277), .B(n3278), .Z(o[8526]) );
  AND U4916 ( .A(p_input[28526]), .B(p_input[18526]), .Z(n3278) );
  AND U4917 ( .A(p_input[8526]), .B(p_input[38526]), .Z(n3277) );
  AND U4918 ( .A(n3279), .B(n3280), .Z(o[8525]) );
  AND U4919 ( .A(p_input[28525]), .B(p_input[18525]), .Z(n3280) );
  AND U4920 ( .A(p_input[8525]), .B(p_input[38525]), .Z(n3279) );
  AND U4921 ( .A(n3281), .B(n3282), .Z(o[8524]) );
  AND U4922 ( .A(p_input[28524]), .B(p_input[18524]), .Z(n3282) );
  AND U4923 ( .A(p_input[8524]), .B(p_input[38524]), .Z(n3281) );
  AND U4924 ( .A(n3283), .B(n3284), .Z(o[8523]) );
  AND U4925 ( .A(p_input[28523]), .B(p_input[18523]), .Z(n3284) );
  AND U4926 ( .A(p_input[8523]), .B(p_input[38523]), .Z(n3283) );
  AND U4927 ( .A(n3285), .B(n3286), .Z(o[8522]) );
  AND U4928 ( .A(p_input[28522]), .B(p_input[18522]), .Z(n3286) );
  AND U4929 ( .A(p_input[8522]), .B(p_input[38522]), .Z(n3285) );
  AND U4930 ( .A(n3287), .B(n3288), .Z(o[8521]) );
  AND U4931 ( .A(p_input[28521]), .B(p_input[18521]), .Z(n3288) );
  AND U4932 ( .A(p_input[8521]), .B(p_input[38521]), .Z(n3287) );
  AND U4933 ( .A(n3289), .B(n3290), .Z(o[8520]) );
  AND U4934 ( .A(p_input[28520]), .B(p_input[18520]), .Z(n3290) );
  AND U4935 ( .A(p_input[8520]), .B(p_input[38520]), .Z(n3289) );
  AND U4936 ( .A(n3291), .B(n3292), .Z(o[851]) );
  AND U4937 ( .A(p_input[20851]), .B(p_input[10851]), .Z(n3292) );
  AND U4938 ( .A(p_input[851]), .B(p_input[30851]), .Z(n3291) );
  AND U4939 ( .A(n3293), .B(n3294), .Z(o[8519]) );
  AND U4940 ( .A(p_input[28519]), .B(p_input[18519]), .Z(n3294) );
  AND U4941 ( .A(p_input[8519]), .B(p_input[38519]), .Z(n3293) );
  AND U4942 ( .A(n3295), .B(n3296), .Z(o[8518]) );
  AND U4943 ( .A(p_input[28518]), .B(p_input[18518]), .Z(n3296) );
  AND U4944 ( .A(p_input[8518]), .B(p_input[38518]), .Z(n3295) );
  AND U4945 ( .A(n3297), .B(n3298), .Z(o[8517]) );
  AND U4946 ( .A(p_input[28517]), .B(p_input[18517]), .Z(n3298) );
  AND U4947 ( .A(p_input[8517]), .B(p_input[38517]), .Z(n3297) );
  AND U4948 ( .A(n3299), .B(n3300), .Z(o[8516]) );
  AND U4949 ( .A(p_input[28516]), .B(p_input[18516]), .Z(n3300) );
  AND U4950 ( .A(p_input[8516]), .B(p_input[38516]), .Z(n3299) );
  AND U4951 ( .A(n3301), .B(n3302), .Z(o[8515]) );
  AND U4952 ( .A(p_input[28515]), .B(p_input[18515]), .Z(n3302) );
  AND U4953 ( .A(p_input[8515]), .B(p_input[38515]), .Z(n3301) );
  AND U4954 ( .A(n3303), .B(n3304), .Z(o[8514]) );
  AND U4955 ( .A(p_input[28514]), .B(p_input[18514]), .Z(n3304) );
  AND U4956 ( .A(p_input[8514]), .B(p_input[38514]), .Z(n3303) );
  AND U4957 ( .A(n3305), .B(n3306), .Z(o[8513]) );
  AND U4958 ( .A(p_input[28513]), .B(p_input[18513]), .Z(n3306) );
  AND U4959 ( .A(p_input[8513]), .B(p_input[38513]), .Z(n3305) );
  AND U4960 ( .A(n3307), .B(n3308), .Z(o[8512]) );
  AND U4961 ( .A(p_input[28512]), .B(p_input[18512]), .Z(n3308) );
  AND U4962 ( .A(p_input[8512]), .B(p_input[38512]), .Z(n3307) );
  AND U4963 ( .A(n3309), .B(n3310), .Z(o[8511]) );
  AND U4964 ( .A(p_input[28511]), .B(p_input[18511]), .Z(n3310) );
  AND U4965 ( .A(p_input[8511]), .B(p_input[38511]), .Z(n3309) );
  AND U4966 ( .A(n3311), .B(n3312), .Z(o[8510]) );
  AND U4967 ( .A(p_input[28510]), .B(p_input[18510]), .Z(n3312) );
  AND U4968 ( .A(p_input[8510]), .B(p_input[38510]), .Z(n3311) );
  AND U4969 ( .A(n3313), .B(n3314), .Z(o[850]) );
  AND U4970 ( .A(p_input[20850]), .B(p_input[10850]), .Z(n3314) );
  AND U4971 ( .A(p_input[850]), .B(p_input[30850]), .Z(n3313) );
  AND U4972 ( .A(n3315), .B(n3316), .Z(o[8509]) );
  AND U4973 ( .A(p_input[28509]), .B(p_input[18509]), .Z(n3316) );
  AND U4974 ( .A(p_input[8509]), .B(p_input[38509]), .Z(n3315) );
  AND U4975 ( .A(n3317), .B(n3318), .Z(o[8508]) );
  AND U4976 ( .A(p_input[28508]), .B(p_input[18508]), .Z(n3318) );
  AND U4977 ( .A(p_input[8508]), .B(p_input[38508]), .Z(n3317) );
  AND U4978 ( .A(n3319), .B(n3320), .Z(o[8507]) );
  AND U4979 ( .A(p_input[28507]), .B(p_input[18507]), .Z(n3320) );
  AND U4980 ( .A(p_input[8507]), .B(p_input[38507]), .Z(n3319) );
  AND U4981 ( .A(n3321), .B(n3322), .Z(o[8506]) );
  AND U4982 ( .A(p_input[28506]), .B(p_input[18506]), .Z(n3322) );
  AND U4983 ( .A(p_input[8506]), .B(p_input[38506]), .Z(n3321) );
  AND U4984 ( .A(n3323), .B(n3324), .Z(o[8505]) );
  AND U4985 ( .A(p_input[28505]), .B(p_input[18505]), .Z(n3324) );
  AND U4986 ( .A(p_input[8505]), .B(p_input[38505]), .Z(n3323) );
  AND U4987 ( .A(n3325), .B(n3326), .Z(o[8504]) );
  AND U4988 ( .A(p_input[28504]), .B(p_input[18504]), .Z(n3326) );
  AND U4989 ( .A(p_input[8504]), .B(p_input[38504]), .Z(n3325) );
  AND U4990 ( .A(n3327), .B(n3328), .Z(o[8503]) );
  AND U4991 ( .A(p_input[28503]), .B(p_input[18503]), .Z(n3328) );
  AND U4992 ( .A(p_input[8503]), .B(p_input[38503]), .Z(n3327) );
  AND U4993 ( .A(n3329), .B(n3330), .Z(o[8502]) );
  AND U4994 ( .A(p_input[28502]), .B(p_input[18502]), .Z(n3330) );
  AND U4995 ( .A(p_input[8502]), .B(p_input[38502]), .Z(n3329) );
  AND U4996 ( .A(n3331), .B(n3332), .Z(o[8501]) );
  AND U4997 ( .A(p_input[28501]), .B(p_input[18501]), .Z(n3332) );
  AND U4998 ( .A(p_input[8501]), .B(p_input[38501]), .Z(n3331) );
  AND U4999 ( .A(n3333), .B(n3334), .Z(o[8500]) );
  AND U5000 ( .A(p_input[28500]), .B(p_input[18500]), .Z(n3334) );
  AND U5001 ( .A(p_input[8500]), .B(p_input[38500]), .Z(n3333) );
  AND U5002 ( .A(n3335), .B(n3336), .Z(o[84]) );
  AND U5003 ( .A(p_input[20084]), .B(p_input[10084]), .Z(n3336) );
  AND U5004 ( .A(p_input[84]), .B(p_input[30084]), .Z(n3335) );
  AND U5005 ( .A(n3337), .B(n3338), .Z(o[849]) );
  AND U5006 ( .A(p_input[20849]), .B(p_input[10849]), .Z(n3338) );
  AND U5007 ( .A(p_input[849]), .B(p_input[30849]), .Z(n3337) );
  AND U5008 ( .A(n3339), .B(n3340), .Z(o[8499]) );
  AND U5009 ( .A(p_input[28499]), .B(p_input[18499]), .Z(n3340) );
  AND U5010 ( .A(p_input[8499]), .B(p_input[38499]), .Z(n3339) );
  AND U5011 ( .A(n3341), .B(n3342), .Z(o[8498]) );
  AND U5012 ( .A(p_input[28498]), .B(p_input[18498]), .Z(n3342) );
  AND U5013 ( .A(p_input[8498]), .B(p_input[38498]), .Z(n3341) );
  AND U5014 ( .A(n3343), .B(n3344), .Z(o[8497]) );
  AND U5015 ( .A(p_input[28497]), .B(p_input[18497]), .Z(n3344) );
  AND U5016 ( .A(p_input[8497]), .B(p_input[38497]), .Z(n3343) );
  AND U5017 ( .A(n3345), .B(n3346), .Z(o[8496]) );
  AND U5018 ( .A(p_input[28496]), .B(p_input[18496]), .Z(n3346) );
  AND U5019 ( .A(p_input[8496]), .B(p_input[38496]), .Z(n3345) );
  AND U5020 ( .A(n3347), .B(n3348), .Z(o[8495]) );
  AND U5021 ( .A(p_input[28495]), .B(p_input[18495]), .Z(n3348) );
  AND U5022 ( .A(p_input[8495]), .B(p_input[38495]), .Z(n3347) );
  AND U5023 ( .A(n3349), .B(n3350), .Z(o[8494]) );
  AND U5024 ( .A(p_input[28494]), .B(p_input[18494]), .Z(n3350) );
  AND U5025 ( .A(p_input[8494]), .B(p_input[38494]), .Z(n3349) );
  AND U5026 ( .A(n3351), .B(n3352), .Z(o[8493]) );
  AND U5027 ( .A(p_input[28493]), .B(p_input[18493]), .Z(n3352) );
  AND U5028 ( .A(p_input[8493]), .B(p_input[38493]), .Z(n3351) );
  AND U5029 ( .A(n3353), .B(n3354), .Z(o[8492]) );
  AND U5030 ( .A(p_input[28492]), .B(p_input[18492]), .Z(n3354) );
  AND U5031 ( .A(p_input[8492]), .B(p_input[38492]), .Z(n3353) );
  AND U5032 ( .A(n3355), .B(n3356), .Z(o[8491]) );
  AND U5033 ( .A(p_input[28491]), .B(p_input[18491]), .Z(n3356) );
  AND U5034 ( .A(p_input[8491]), .B(p_input[38491]), .Z(n3355) );
  AND U5035 ( .A(n3357), .B(n3358), .Z(o[8490]) );
  AND U5036 ( .A(p_input[28490]), .B(p_input[18490]), .Z(n3358) );
  AND U5037 ( .A(p_input[8490]), .B(p_input[38490]), .Z(n3357) );
  AND U5038 ( .A(n3359), .B(n3360), .Z(o[848]) );
  AND U5039 ( .A(p_input[20848]), .B(p_input[10848]), .Z(n3360) );
  AND U5040 ( .A(p_input[848]), .B(p_input[30848]), .Z(n3359) );
  AND U5041 ( .A(n3361), .B(n3362), .Z(o[8489]) );
  AND U5042 ( .A(p_input[28489]), .B(p_input[18489]), .Z(n3362) );
  AND U5043 ( .A(p_input[8489]), .B(p_input[38489]), .Z(n3361) );
  AND U5044 ( .A(n3363), .B(n3364), .Z(o[8488]) );
  AND U5045 ( .A(p_input[28488]), .B(p_input[18488]), .Z(n3364) );
  AND U5046 ( .A(p_input[8488]), .B(p_input[38488]), .Z(n3363) );
  AND U5047 ( .A(n3365), .B(n3366), .Z(o[8487]) );
  AND U5048 ( .A(p_input[28487]), .B(p_input[18487]), .Z(n3366) );
  AND U5049 ( .A(p_input[8487]), .B(p_input[38487]), .Z(n3365) );
  AND U5050 ( .A(n3367), .B(n3368), .Z(o[8486]) );
  AND U5051 ( .A(p_input[28486]), .B(p_input[18486]), .Z(n3368) );
  AND U5052 ( .A(p_input[8486]), .B(p_input[38486]), .Z(n3367) );
  AND U5053 ( .A(n3369), .B(n3370), .Z(o[8485]) );
  AND U5054 ( .A(p_input[28485]), .B(p_input[18485]), .Z(n3370) );
  AND U5055 ( .A(p_input[8485]), .B(p_input[38485]), .Z(n3369) );
  AND U5056 ( .A(n3371), .B(n3372), .Z(o[8484]) );
  AND U5057 ( .A(p_input[28484]), .B(p_input[18484]), .Z(n3372) );
  AND U5058 ( .A(p_input[8484]), .B(p_input[38484]), .Z(n3371) );
  AND U5059 ( .A(n3373), .B(n3374), .Z(o[8483]) );
  AND U5060 ( .A(p_input[28483]), .B(p_input[18483]), .Z(n3374) );
  AND U5061 ( .A(p_input[8483]), .B(p_input[38483]), .Z(n3373) );
  AND U5062 ( .A(n3375), .B(n3376), .Z(o[8482]) );
  AND U5063 ( .A(p_input[28482]), .B(p_input[18482]), .Z(n3376) );
  AND U5064 ( .A(p_input[8482]), .B(p_input[38482]), .Z(n3375) );
  AND U5065 ( .A(n3377), .B(n3378), .Z(o[8481]) );
  AND U5066 ( .A(p_input[28481]), .B(p_input[18481]), .Z(n3378) );
  AND U5067 ( .A(p_input[8481]), .B(p_input[38481]), .Z(n3377) );
  AND U5068 ( .A(n3379), .B(n3380), .Z(o[8480]) );
  AND U5069 ( .A(p_input[28480]), .B(p_input[18480]), .Z(n3380) );
  AND U5070 ( .A(p_input[8480]), .B(p_input[38480]), .Z(n3379) );
  AND U5071 ( .A(n3381), .B(n3382), .Z(o[847]) );
  AND U5072 ( .A(p_input[20847]), .B(p_input[10847]), .Z(n3382) );
  AND U5073 ( .A(p_input[847]), .B(p_input[30847]), .Z(n3381) );
  AND U5074 ( .A(n3383), .B(n3384), .Z(o[8479]) );
  AND U5075 ( .A(p_input[28479]), .B(p_input[18479]), .Z(n3384) );
  AND U5076 ( .A(p_input[8479]), .B(p_input[38479]), .Z(n3383) );
  AND U5077 ( .A(n3385), .B(n3386), .Z(o[8478]) );
  AND U5078 ( .A(p_input[28478]), .B(p_input[18478]), .Z(n3386) );
  AND U5079 ( .A(p_input[8478]), .B(p_input[38478]), .Z(n3385) );
  AND U5080 ( .A(n3387), .B(n3388), .Z(o[8477]) );
  AND U5081 ( .A(p_input[28477]), .B(p_input[18477]), .Z(n3388) );
  AND U5082 ( .A(p_input[8477]), .B(p_input[38477]), .Z(n3387) );
  AND U5083 ( .A(n3389), .B(n3390), .Z(o[8476]) );
  AND U5084 ( .A(p_input[28476]), .B(p_input[18476]), .Z(n3390) );
  AND U5085 ( .A(p_input[8476]), .B(p_input[38476]), .Z(n3389) );
  AND U5086 ( .A(n3391), .B(n3392), .Z(o[8475]) );
  AND U5087 ( .A(p_input[28475]), .B(p_input[18475]), .Z(n3392) );
  AND U5088 ( .A(p_input[8475]), .B(p_input[38475]), .Z(n3391) );
  AND U5089 ( .A(n3393), .B(n3394), .Z(o[8474]) );
  AND U5090 ( .A(p_input[28474]), .B(p_input[18474]), .Z(n3394) );
  AND U5091 ( .A(p_input[8474]), .B(p_input[38474]), .Z(n3393) );
  AND U5092 ( .A(n3395), .B(n3396), .Z(o[8473]) );
  AND U5093 ( .A(p_input[28473]), .B(p_input[18473]), .Z(n3396) );
  AND U5094 ( .A(p_input[8473]), .B(p_input[38473]), .Z(n3395) );
  AND U5095 ( .A(n3397), .B(n3398), .Z(o[8472]) );
  AND U5096 ( .A(p_input[28472]), .B(p_input[18472]), .Z(n3398) );
  AND U5097 ( .A(p_input[8472]), .B(p_input[38472]), .Z(n3397) );
  AND U5098 ( .A(n3399), .B(n3400), .Z(o[8471]) );
  AND U5099 ( .A(p_input[28471]), .B(p_input[18471]), .Z(n3400) );
  AND U5100 ( .A(p_input[8471]), .B(p_input[38471]), .Z(n3399) );
  AND U5101 ( .A(n3401), .B(n3402), .Z(o[8470]) );
  AND U5102 ( .A(p_input[28470]), .B(p_input[18470]), .Z(n3402) );
  AND U5103 ( .A(p_input[8470]), .B(p_input[38470]), .Z(n3401) );
  AND U5104 ( .A(n3403), .B(n3404), .Z(o[846]) );
  AND U5105 ( .A(p_input[20846]), .B(p_input[10846]), .Z(n3404) );
  AND U5106 ( .A(p_input[846]), .B(p_input[30846]), .Z(n3403) );
  AND U5107 ( .A(n3405), .B(n3406), .Z(o[8469]) );
  AND U5108 ( .A(p_input[28469]), .B(p_input[18469]), .Z(n3406) );
  AND U5109 ( .A(p_input[8469]), .B(p_input[38469]), .Z(n3405) );
  AND U5110 ( .A(n3407), .B(n3408), .Z(o[8468]) );
  AND U5111 ( .A(p_input[28468]), .B(p_input[18468]), .Z(n3408) );
  AND U5112 ( .A(p_input[8468]), .B(p_input[38468]), .Z(n3407) );
  AND U5113 ( .A(n3409), .B(n3410), .Z(o[8467]) );
  AND U5114 ( .A(p_input[28467]), .B(p_input[18467]), .Z(n3410) );
  AND U5115 ( .A(p_input[8467]), .B(p_input[38467]), .Z(n3409) );
  AND U5116 ( .A(n3411), .B(n3412), .Z(o[8466]) );
  AND U5117 ( .A(p_input[28466]), .B(p_input[18466]), .Z(n3412) );
  AND U5118 ( .A(p_input[8466]), .B(p_input[38466]), .Z(n3411) );
  AND U5119 ( .A(n3413), .B(n3414), .Z(o[8465]) );
  AND U5120 ( .A(p_input[28465]), .B(p_input[18465]), .Z(n3414) );
  AND U5121 ( .A(p_input[8465]), .B(p_input[38465]), .Z(n3413) );
  AND U5122 ( .A(n3415), .B(n3416), .Z(o[8464]) );
  AND U5123 ( .A(p_input[28464]), .B(p_input[18464]), .Z(n3416) );
  AND U5124 ( .A(p_input[8464]), .B(p_input[38464]), .Z(n3415) );
  AND U5125 ( .A(n3417), .B(n3418), .Z(o[8463]) );
  AND U5126 ( .A(p_input[28463]), .B(p_input[18463]), .Z(n3418) );
  AND U5127 ( .A(p_input[8463]), .B(p_input[38463]), .Z(n3417) );
  AND U5128 ( .A(n3419), .B(n3420), .Z(o[8462]) );
  AND U5129 ( .A(p_input[28462]), .B(p_input[18462]), .Z(n3420) );
  AND U5130 ( .A(p_input[8462]), .B(p_input[38462]), .Z(n3419) );
  AND U5131 ( .A(n3421), .B(n3422), .Z(o[8461]) );
  AND U5132 ( .A(p_input[28461]), .B(p_input[18461]), .Z(n3422) );
  AND U5133 ( .A(p_input[8461]), .B(p_input[38461]), .Z(n3421) );
  AND U5134 ( .A(n3423), .B(n3424), .Z(o[8460]) );
  AND U5135 ( .A(p_input[28460]), .B(p_input[18460]), .Z(n3424) );
  AND U5136 ( .A(p_input[8460]), .B(p_input[38460]), .Z(n3423) );
  AND U5137 ( .A(n3425), .B(n3426), .Z(o[845]) );
  AND U5138 ( .A(p_input[20845]), .B(p_input[10845]), .Z(n3426) );
  AND U5139 ( .A(p_input[845]), .B(p_input[30845]), .Z(n3425) );
  AND U5140 ( .A(n3427), .B(n3428), .Z(o[8459]) );
  AND U5141 ( .A(p_input[28459]), .B(p_input[18459]), .Z(n3428) );
  AND U5142 ( .A(p_input[8459]), .B(p_input[38459]), .Z(n3427) );
  AND U5143 ( .A(n3429), .B(n3430), .Z(o[8458]) );
  AND U5144 ( .A(p_input[28458]), .B(p_input[18458]), .Z(n3430) );
  AND U5145 ( .A(p_input[8458]), .B(p_input[38458]), .Z(n3429) );
  AND U5146 ( .A(n3431), .B(n3432), .Z(o[8457]) );
  AND U5147 ( .A(p_input[28457]), .B(p_input[18457]), .Z(n3432) );
  AND U5148 ( .A(p_input[8457]), .B(p_input[38457]), .Z(n3431) );
  AND U5149 ( .A(n3433), .B(n3434), .Z(o[8456]) );
  AND U5150 ( .A(p_input[28456]), .B(p_input[18456]), .Z(n3434) );
  AND U5151 ( .A(p_input[8456]), .B(p_input[38456]), .Z(n3433) );
  AND U5152 ( .A(n3435), .B(n3436), .Z(o[8455]) );
  AND U5153 ( .A(p_input[28455]), .B(p_input[18455]), .Z(n3436) );
  AND U5154 ( .A(p_input[8455]), .B(p_input[38455]), .Z(n3435) );
  AND U5155 ( .A(n3437), .B(n3438), .Z(o[8454]) );
  AND U5156 ( .A(p_input[28454]), .B(p_input[18454]), .Z(n3438) );
  AND U5157 ( .A(p_input[8454]), .B(p_input[38454]), .Z(n3437) );
  AND U5158 ( .A(n3439), .B(n3440), .Z(o[8453]) );
  AND U5159 ( .A(p_input[28453]), .B(p_input[18453]), .Z(n3440) );
  AND U5160 ( .A(p_input[8453]), .B(p_input[38453]), .Z(n3439) );
  AND U5161 ( .A(n3441), .B(n3442), .Z(o[8452]) );
  AND U5162 ( .A(p_input[28452]), .B(p_input[18452]), .Z(n3442) );
  AND U5163 ( .A(p_input[8452]), .B(p_input[38452]), .Z(n3441) );
  AND U5164 ( .A(n3443), .B(n3444), .Z(o[8451]) );
  AND U5165 ( .A(p_input[28451]), .B(p_input[18451]), .Z(n3444) );
  AND U5166 ( .A(p_input[8451]), .B(p_input[38451]), .Z(n3443) );
  AND U5167 ( .A(n3445), .B(n3446), .Z(o[8450]) );
  AND U5168 ( .A(p_input[28450]), .B(p_input[18450]), .Z(n3446) );
  AND U5169 ( .A(p_input[8450]), .B(p_input[38450]), .Z(n3445) );
  AND U5170 ( .A(n3447), .B(n3448), .Z(o[844]) );
  AND U5171 ( .A(p_input[20844]), .B(p_input[10844]), .Z(n3448) );
  AND U5172 ( .A(p_input[844]), .B(p_input[30844]), .Z(n3447) );
  AND U5173 ( .A(n3449), .B(n3450), .Z(o[8449]) );
  AND U5174 ( .A(p_input[28449]), .B(p_input[18449]), .Z(n3450) );
  AND U5175 ( .A(p_input[8449]), .B(p_input[38449]), .Z(n3449) );
  AND U5176 ( .A(n3451), .B(n3452), .Z(o[8448]) );
  AND U5177 ( .A(p_input[28448]), .B(p_input[18448]), .Z(n3452) );
  AND U5178 ( .A(p_input[8448]), .B(p_input[38448]), .Z(n3451) );
  AND U5179 ( .A(n3453), .B(n3454), .Z(o[8447]) );
  AND U5180 ( .A(p_input[28447]), .B(p_input[18447]), .Z(n3454) );
  AND U5181 ( .A(p_input[8447]), .B(p_input[38447]), .Z(n3453) );
  AND U5182 ( .A(n3455), .B(n3456), .Z(o[8446]) );
  AND U5183 ( .A(p_input[28446]), .B(p_input[18446]), .Z(n3456) );
  AND U5184 ( .A(p_input[8446]), .B(p_input[38446]), .Z(n3455) );
  AND U5185 ( .A(n3457), .B(n3458), .Z(o[8445]) );
  AND U5186 ( .A(p_input[28445]), .B(p_input[18445]), .Z(n3458) );
  AND U5187 ( .A(p_input[8445]), .B(p_input[38445]), .Z(n3457) );
  AND U5188 ( .A(n3459), .B(n3460), .Z(o[8444]) );
  AND U5189 ( .A(p_input[28444]), .B(p_input[18444]), .Z(n3460) );
  AND U5190 ( .A(p_input[8444]), .B(p_input[38444]), .Z(n3459) );
  AND U5191 ( .A(n3461), .B(n3462), .Z(o[8443]) );
  AND U5192 ( .A(p_input[28443]), .B(p_input[18443]), .Z(n3462) );
  AND U5193 ( .A(p_input[8443]), .B(p_input[38443]), .Z(n3461) );
  AND U5194 ( .A(n3463), .B(n3464), .Z(o[8442]) );
  AND U5195 ( .A(p_input[28442]), .B(p_input[18442]), .Z(n3464) );
  AND U5196 ( .A(p_input[8442]), .B(p_input[38442]), .Z(n3463) );
  AND U5197 ( .A(n3465), .B(n3466), .Z(o[8441]) );
  AND U5198 ( .A(p_input[28441]), .B(p_input[18441]), .Z(n3466) );
  AND U5199 ( .A(p_input[8441]), .B(p_input[38441]), .Z(n3465) );
  AND U5200 ( .A(n3467), .B(n3468), .Z(o[8440]) );
  AND U5201 ( .A(p_input[28440]), .B(p_input[18440]), .Z(n3468) );
  AND U5202 ( .A(p_input[8440]), .B(p_input[38440]), .Z(n3467) );
  AND U5203 ( .A(n3469), .B(n3470), .Z(o[843]) );
  AND U5204 ( .A(p_input[20843]), .B(p_input[10843]), .Z(n3470) );
  AND U5205 ( .A(p_input[843]), .B(p_input[30843]), .Z(n3469) );
  AND U5206 ( .A(n3471), .B(n3472), .Z(o[8439]) );
  AND U5207 ( .A(p_input[28439]), .B(p_input[18439]), .Z(n3472) );
  AND U5208 ( .A(p_input[8439]), .B(p_input[38439]), .Z(n3471) );
  AND U5209 ( .A(n3473), .B(n3474), .Z(o[8438]) );
  AND U5210 ( .A(p_input[28438]), .B(p_input[18438]), .Z(n3474) );
  AND U5211 ( .A(p_input[8438]), .B(p_input[38438]), .Z(n3473) );
  AND U5212 ( .A(n3475), .B(n3476), .Z(o[8437]) );
  AND U5213 ( .A(p_input[28437]), .B(p_input[18437]), .Z(n3476) );
  AND U5214 ( .A(p_input[8437]), .B(p_input[38437]), .Z(n3475) );
  AND U5215 ( .A(n3477), .B(n3478), .Z(o[8436]) );
  AND U5216 ( .A(p_input[28436]), .B(p_input[18436]), .Z(n3478) );
  AND U5217 ( .A(p_input[8436]), .B(p_input[38436]), .Z(n3477) );
  AND U5218 ( .A(n3479), .B(n3480), .Z(o[8435]) );
  AND U5219 ( .A(p_input[28435]), .B(p_input[18435]), .Z(n3480) );
  AND U5220 ( .A(p_input[8435]), .B(p_input[38435]), .Z(n3479) );
  AND U5221 ( .A(n3481), .B(n3482), .Z(o[8434]) );
  AND U5222 ( .A(p_input[28434]), .B(p_input[18434]), .Z(n3482) );
  AND U5223 ( .A(p_input[8434]), .B(p_input[38434]), .Z(n3481) );
  AND U5224 ( .A(n3483), .B(n3484), .Z(o[8433]) );
  AND U5225 ( .A(p_input[28433]), .B(p_input[18433]), .Z(n3484) );
  AND U5226 ( .A(p_input[8433]), .B(p_input[38433]), .Z(n3483) );
  AND U5227 ( .A(n3485), .B(n3486), .Z(o[8432]) );
  AND U5228 ( .A(p_input[28432]), .B(p_input[18432]), .Z(n3486) );
  AND U5229 ( .A(p_input[8432]), .B(p_input[38432]), .Z(n3485) );
  AND U5230 ( .A(n3487), .B(n3488), .Z(o[8431]) );
  AND U5231 ( .A(p_input[28431]), .B(p_input[18431]), .Z(n3488) );
  AND U5232 ( .A(p_input[8431]), .B(p_input[38431]), .Z(n3487) );
  AND U5233 ( .A(n3489), .B(n3490), .Z(o[8430]) );
  AND U5234 ( .A(p_input[28430]), .B(p_input[18430]), .Z(n3490) );
  AND U5235 ( .A(p_input[8430]), .B(p_input[38430]), .Z(n3489) );
  AND U5236 ( .A(n3491), .B(n3492), .Z(o[842]) );
  AND U5237 ( .A(p_input[20842]), .B(p_input[10842]), .Z(n3492) );
  AND U5238 ( .A(p_input[842]), .B(p_input[30842]), .Z(n3491) );
  AND U5239 ( .A(n3493), .B(n3494), .Z(o[8429]) );
  AND U5240 ( .A(p_input[28429]), .B(p_input[18429]), .Z(n3494) );
  AND U5241 ( .A(p_input[8429]), .B(p_input[38429]), .Z(n3493) );
  AND U5242 ( .A(n3495), .B(n3496), .Z(o[8428]) );
  AND U5243 ( .A(p_input[28428]), .B(p_input[18428]), .Z(n3496) );
  AND U5244 ( .A(p_input[8428]), .B(p_input[38428]), .Z(n3495) );
  AND U5245 ( .A(n3497), .B(n3498), .Z(o[8427]) );
  AND U5246 ( .A(p_input[28427]), .B(p_input[18427]), .Z(n3498) );
  AND U5247 ( .A(p_input[8427]), .B(p_input[38427]), .Z(n3497) );
  AND U5248 ( .A(n3499), .B(n3500), .Z(o[8426]) );
  AND U5249 ( .A(p_input[28426]), .B(p_input[18426]), .Z(n3500) );
  AND U5250 ( .A(p_input[8426]), .B(p_input[38426]), .Z(n3499) );
  AND U5251 ( .A(n3501), .B(n3502), .Z(o[8425]) );
  AND U5252 ( .A(p_input[28425]), .B(p_input[18425]), .Z(n3502) );
  AND U5253 ( .A(p_input[8425]), .B(p_input[38425]), .Z(n3501) );
  AND U5254 ( .A(n3503), .B(n3504), .Z(o[8424]) );
  AND U5255 ( .A(p_input[28424]), .B(p_input[18424]), .Z(n3504) );
  AND U5256 ( .A(p_input[8424]), .B(p_input[38424]), .Z(n3503) );
  AND U5257 ( .A(n3505), .B(n3506), .Z(o[8423]) );
  AND U5258 ( .A(p_input[28423]), .B(p_input[18423]), .Z(n3506) );
  AND U5259 ( .A(p_input[8423]), .B(p_input[38423]), .Z(n3505) );
  AND U5260 ( .A(n3507), .B(n3508), .Z(o[8422]) );
  AND U5261 ( .A(p_input[28422]), .B(p_input[18422]), .Z(n3508) );
  AND U5262 ( .A(p_input[8422]), .B(p_input[38422]), .Z(n3507) );
  AND U5263 ( .A(n3509), .B(n3510), .Z(o[8421]) );
  AND U5264 ( .A(p_input[28421]), .B(p_input[18421]), .Z(n3510) );
  AND U5265 ( .A(p_input[8421]), .B(p_input[38421]), .Z(n3509) );
  AND U5266 ( .A(n3511), .B(n3512), .Z(o[8420]) );
  AND U5267 ( .A(p_input[28420]), .B(p_input[18420]), .Z(n3512) );
  AND U5268 ( .A(p_input[8420]), .B(p_input[38420]), .Z(n3511) );
  AND U5269 ( .A(n3513), .B(n3514), .Z(o[841]) );
  AND U5270 ( .A(p_input[20841]), .B(p_input[10841]), .Z(n3514) );
  AND U5271 ( .A(p_input[841]), .B(p_input[30841]), .Z(n3513) );
  AND U5272 ( .A(n3515), .B(n3516), .Z(o[8419]) );
  AND U5273 ( .A(p_input[28419]), .B(p_input[18419]), .Z(n3516) );
  AND U5274 ( .A(p_input[8419]), .B(p_input[38419]), .Z(n3515) );
  AND U5275 ( .A(n3517), .B(n3518), .Z(o[8418]) );
  AND U5276 ( .A(p_input[28418]), .B(p_input[18418]), .Z(n3518) );
  AND U5277 ( .A(p_input[8418]), .B(p_input[38418]), .Z(n3517) );
  AND U5278 ( .A(n3519), .B(n3520), .Z(o[8417]) );
  AND U5279 ( .A(p_input[28417]), .B(p_input[18417]), .Z(n3520) );
  AND U5280 ( .A(p_input[8417]), .B(p_input[38417]), .Z(n3519) );
  AND U5281 ( .A(n3521), .B(n3522), .Z(o[8416]) );
  AND U5282 ( .A(p_input[28416]), .B(p_input[18416]), .Z(n3522) );
  AND U5283 ( .A(p_input[8416]), .B(p_input[38416]), .Z(n3521) );
  AND U5284 ( .A(n3523), .B(n3524), .Z(o[8415]) );
  AND U5285 ( .A(p_input[28415]), .B(p_input[18415]), .Z(n3524) );
  AND U5286 ( .A(p_input[8415]), .B(p_input[38415]), .Z(n3523) );
  AND U5287 ( .A(n3525), .B(n3526), .Z(o[8414]) );
  AND U5288 ( .A(p_input[28414]), .B(p_input[18414]), .Z(n3526) );
  AND U5289 ( .A(p_input[8414]), .B(p_input[38414]), .Z(n3525) );
  AND U5290 ( .A(n3527), .B(n3528), .Z(o[8413]) );
  AND U5291 ( .A(p_input[28413]), .B(p_input[18413]), .Z(n3528) );
  AND U5292 ( .A(p_input[8413]), .B(p_input[38413]), .Z(n3527) );
  AND U5293 ( .A(n3529), .B(n3530), .Z(o[8412]) );
  AND U5294 ( .A(p_input[28412]), .B(p_input[18412]), .Z(n3530) );
  AND U5295 ( .A(p_input[8412]), .B(p_input[38412]), .Z(n3529) );
  AND U5296 ( .A(n3531), .B(n3532), .Z(o[8411]) );
  AND U5297 ( .A(p_input[28411]), .B(p_input[18411]), .Z(n3532) );
  AND U5298 ( .A(p_input[8411]), .B(p_input[38411]), .Z(n3531) );
  AND U5299 ( .A(n3533), .B(n3534), .Z(o[8410]) );
  AND U5300 ( .A(p_input[28410]), .B(p_input[18410]), .Z(n3534) );
  AND U5301 ( .A(p_input[8410]), .B(p_input[38410]), .Z(n3533) );
  AND U5302 ( .A(n3535), .B(n3536), .Z(o[840]) );
  AND U5303 ( .A(p_input[20840]), .B(p_input[10840]), .Z(n3536) );
  AND U5304 ( .A(p_input[840]), .B(p_input[30840]), .Z(n3535) );
  AND U5305 ( .A(n3537), .B(n3538), .Z(o[8409]) );
  AND U5306 ( .A(p_input[28409]), .B(p_input[18409]), .Z(n3538) );
  AND U5307 ( .A(p_input[8409]), .B(p_input[38409]), .Z(n3537) );
  AND U5308 ( .A(n3539), .B(n3540), .Z(o[8408]) );
  AND U5309 ( .A(p_input[28408]), .B(p_input[18408]), .Z(n3540) );
  AND U5310 ( .A(p_input[8408]), .B(p_input[38408]), .Z(n3539) );
  AND U5311 ( .A(n3541), .B(n3542), .Z(o[8407]) );
  AND U5312 ( .A(p_input[28407]), .B(p_input[18407]), .Z(n3542) );
  AND U5313 ( .A(p_input[8407]), .B(p_input[38407]), .Z(n3541) );
  AND U5314 ( .A(n3543), .B(n3544), .Z(o[8406]) );
  AND U5315 ( .A(p_input[28406]), .B(p_input[18406]), .Z(n3544) );
  AND U5316 ( .A(p_input[8406]), .B(p_input[38406]), .Z(n3543) );
  AND U5317 ( .A(n3545), .B(n3546), .Z(o[8405]) );
  AND U5318 ( .A(p_input[28405]), .B(p_input[18405]), .Z(n3546) );
  AND U5319 ( .A(p_input[8405]), .B(p_input[38405]), .Z(n3545) );
  AND U5320 ( .A(n3547), .B(n3548), .Z(o[8404]) );
  AND U5321 ( .A(p_input[28404]), .B(p_input[18404]), .Z(n3548) );
  AND U5322 ( .A(p_input[8404]), .B(p_input[38404]), .Z(n3547) );
  AND U5323 ( .A(n3549), .B(n3550), .Z(o[8403]) );
  AND U5324 ( .A(p_input[28403]), .B(p_input[18403]), .Z(n3550) );
  AND U5325 ( .A(p_input[8403]), .B(p_input[38403]), .Z(n3549) );
  AND U5326 ( .A(n3551), .B(n3552), .Z(o[8402]) );
  AND U5327 ( .A(p_input[28402]), .B(p_input[18402]), .Z(n3552) );
  AND U5328 ( .A(p_input[8402]), .B(p_input[38402]), .Z(n3551) );
  AND U5329 ( .A(n3553), .B(n3554), .Z(o[8401]) );
  AND U5330 ( .A(p_input[28401]), .B(p_input[18401]), .Z(n3554) );
  AND U5331 ( .A(p_input[8401]), .B(p_input[38401]), .Z(n3553) );
  AND U5332 ( .A(n3555), .B(n3556), .Z(o[8400]) );
  AND U5333 ( .A(p_input[28400]), .B(p_input[18400]), .Z(n3556) );
  AND U5334 ( .A(p_input[8400]), .B(p_input[38400]), .Z(n3555) );
  AND U5335 ( .A(n3557), .B(n3558), .Z(o[83]) );
  AND U5336 ( .A(p_input[20083]), .B(p_input[10083]), .Z(n3558) );
  AND U5337 ( .A(p_input[83]), .B(p_input[30083]), .Z(n3557) );
  AND U5338 ( .A(n3559), .B(n3560), .Z(o[839]) );
  AND U5339 ( .A(p_input[20839]), .B(p_input[10839]), .Z(n3560) );
  AND U5340 ( .A(p_input[839]), .B(p_input[30839]), .Z(n3559) );
  AND U5341 ( .A(n3561), .B(n3562), .Z(o[8399]) );
  AND U5342 ( .A(p_input[28399]), .B(p_input[18399]), .Z(n3562) );
  AND U5343 ( .A(p_input[8399]), .B(p_input[38399]), .Z(n3561) );
  AND U5344 ( .A(n3563), .B(n3564), .Z(o[8398]) );
  AND U5345 ( .A(p_input[28398]), .B(p_input[18398]), .Z(n3564) );
  AND U5346 ( .A(p_input[8398]), .B(p_input[38398]), .Z(n3563) );
  AND U5347 ( .A(n3565), .B(n3566), .Z(o[8397]) );
  AND U5348 ( .A(p_input[28397]), .B(p_input[18397]), .Z(n3566) );
  AND U5349 ( .A(p_input[8397]), .B(p_input[38397]), .Z(n3565) );
  AND U5350 ( .A(n3567), .B(n3568), .Z(o[8396]) );
  AND U5351 ( .A(p_input[28396]), .B(p_input[18396]), .Z(n3568) );
  AND U5352 ( .A(p_input[8396]), .B(p_input[38396]), .Z(n3567) );
  AND U5353 ( .A(n3569), .B(n3570), .Z(o[8395]) );
  AND U5354 ( .A(p_input[28395]), .B(p_input[18395]), .Z(n3570) );
  AND U5355 ( .A(p_input[8395]), .B(p_input[38395]), .Z(n3569) );
  AND U5356 ( .A(n3571), .B(n3572), .Z(o[8394]) );
  AND U5357 ( .A(p_input[28394]), .B(p_input[18394]), .Z(n3572) );
  AND U5358 ( .A(p_input[8394]), .B(p_input[38394]), .Z(n3571) );
  AND U5359 ( .A(n3573), .B(n3574), .Z(o[8393]) );
  AND U5360 ( .A(p_input[28393]), .B(p_input[18393]), .Z(n3574) );
  AND U5361 ( .A(p_input[8393]), .B(p_input[38393]), .Z(n3573) );
  AND U5362 ( .A(n3575), .B(n3576), .Z(o[8392]) );
  AND U5363 ( .A(p_input[28392]), .B(p_input[18392]), .Z(n3576) );
  AND U5364 ( .A(p_input[8392]), .B(p_input[38392]), .Z(n3575) );
  AND U5365 ( .A(n3577), .B(n3578), .Z(o[8391]) );
  AND U5366 ( .A(p_input[28391]), .B(p_input[18391]), .Z(n3578) );
  AND U5367 ( .A(p_input[8391]), .B(p_input[38391]), .Z(n3577) );
  AND U5368 ( .A(n3579), .B(n3580), .Z(o[8390]) );
  AND U5369 ( .A(p_input[28390]), .B(p_input[18390]), .Z(n3580) );
  AND U5370 ( .A(p_input[8390]), .B(p_input[38390]), .Z(n3579) );
  AND U5371 ( .A(n3581), .B(n3582), .Z(o[838]) );
  AND U5372 ( .A(p_input[20838]), .B(p_input[10838]), .Z(n3582) );
  AND U5373 ( .A(p_input[838]), .B(p_input[30838]), .Z(n3581) );
  AND U5374 ( .A(n3583), .B(n3584), .Z(o[8389]) );
  AND U5375 ( .A(p_input[28389]), .B(p_input[18389]), .Z(n3584) );
  AND U5376 ( .A(p_input[8389]), .B(p_input[38389]), .Z(n3583) );
  AND U5377 ( .A(n3585), .B(n3586), .Z(o[8388]) );
  AND U5378 ( .A(p_input[28388]), .B(p_input[18388]), .Z(n3586) );
  AND U5379 ( .A(p_input[8388]), .B(p_input[38388]), .Z(n3585) );
  AND U5380 ( .A(n3587), .B(n3588), .Z(o[8387]) );
  AND U5381 ( .A(p_input[28387]), .B(p_input[18387]), .Z(n3588) );
  AND U5382 ( .A(p_input[8387]), .B(p_input[38387]), .Z(n3587) );
  AND U5383 ( .A(n3589), .B(n3590), .Z(o[8386]) );
  AND U5384 ( .A(p_input[28386]), .B(p_input[18386]), .Z(n3590) );
  AND U5385 ( .A(p_input[8386]), .B(p_input[38386]), .Z(n3589) );
  AND U5386 ( .A(n3591), .B(n3592), .Z(o[8385]) );
  AND U5387 ( .A(p_input[28385]), .B(p_input[18385]), .Z(n3592) );
  AND U5388 ( .A(p_input[8385]), .B(p_input[38385]), .Z(n3591) );
  AND U5389 ( .A(n3593), .B(n3594), .Z(o[8384]) );
  AND U5390 ( .A(p_input[28384]), .B(p_input[18384]), .Z(n3594) );
  AND U5391 ( .A(p_input[8384]), .B(p_input[38384]), .Z(n3593) );
  AND U5392 ( .A(n3595), .B(n3596), .Z(o[8383]) );
  AND U5393 ( .A(p_input[28383]), .B(p_input[18383]), .Z(n3596) );
  AND U5394 ( .A(p_input[8383]), .B(p_input[38383]), .Z(n3595) );
  AND U5395 ( .A(n3597), .B(n3598), .Z(o[8382]) );
  AND U5396 ( .A(p_input[28382]), .B(p_input[18382]), .Z(n3598) );
  AND U5397 ( .A(p_input[8382]), .B(p_input[38382]), .Z(n3597) );
  AND U5398 ( .A(n3599), .B(n3600), .Z(o[8381]) );
  AND U5399 ( .A(p_input[28381]), .B(p_input[18381]), .Z(n3600) );
  AND U5400 ( .A(p_input[8381]), .B(p_input[38381]), .Z(n3599) );
  AND U5401 ( .A(n3601), .B(n3602), .Z(o[8380]) );
  AND U5402 ( .A(p_input[28380]), .B(p_input[18380]), .Z(n3602) );
  AND U5403 ( .A(p_input[8380]), .B(p_input[38380]), .Z(n3601) );
  AND U5404 ( .A(n3603), .B(n3604), .Z(o[837]) );
  AND U5405 ( .A(p_input[20837]), .B(p_input[10837]), .Z(n3604) );
  AND U5406 ( .A(p_input[837]), .B(p_input[30837]), .Z(n3603) );
  AND U5407 ( .A(n3605), .B(n3606), .Z(o[8379]) );
  AND U5408 ( .A(p_input[28379]), .B(p_input[18379]), .Z(n3606) );
  AND U5409 ( .A(p_input[8379]), .B(p_input[38379]), .Z(n3605) );
  AND U5410 ( .A(n3607), .B(n3608), .Z(o[8378]) );
  AND U5411 ( .A(p_input[28378]), .B(p_input[18378]), .Z(n3608) );
  AND U5412 ( .A(p_input[8378]), .B(p_input[38378]), .Z(n3607) );
  AND U5413 ( .A(n3609), .B(n3610), .Z(o[8377]) );
  AND U5414 ( .A(p_input[28377]), .B(p_input[18377]), .Z(n3610) );
  AND U5415 ( .A(p_input[8377]), .B(p_input[38377]), .Z(n3609) );
  AND U5416 ( .A(n3611), .B(n3612), .Z(o[8376]) );
  AND U5417 ( .A(p_input[28376]), .B(p_input[18376]), .Z(n3612) );
  AND U5418 ( .A(p_input[8376]), .B(p_input[38376]), .Z(n3611) );
  AND U5419 ( .A(n3613), .B(n3614), .Z(o[8375]) );
  AND U5420 ( .A(p_input[28375]), .B(p_input[18375]), .Z(n3614) );
  AND U5421 ( .A(p_input[8375]), .B(p_input[38375]), .Z(n3613) );
  AND U5422 ( .A(n3615), .B(n3616), .Z(o[8374]) );
  AND U5423 ( .A(p_input[28374]), .B(p_input[18374]), .Z(n3616) );
  AND U5424 ( .A(p_input[8374]), .B(p_input[38374]), .Z(n3615) );
  AND U5425 ( .A(n3617), .B(n3618), .Z(o[8373]) );
  AND U5426 ( .A(p_input[28373]), .B(p_input[18373]), .Z(n3618) );
  AND U5427 ( .A(p_input[8373]), .B(p_input[38373]), .Z(n3617) );
  AND U5428 ( .A(n3619), .B(n3620), .Z(o[8372]) );
  AND U5429 ( .A(p_input[28372]), .B(p_input[18372]), .Z(n3620) );
  AND U5430 ( .A(p_input[8372]), .B(p_input[38372]), .Z(n3619) );
  AND U5431 ( .A(n3621), .B(n3622), .Z(o[8371]) );
  AND U5432 ( .A(p_input[28371]), .B(p_input[18371]), .Z(n3622) );
  AND U5433 ( .A(p_input[8371]), .B(p_input[38371]), .Z(n3621) );
  AND U5434 ( .A(n3623), .B(n3624), .Z(o[8370]) );
  AND U5435 ( .A(p_input[28370]), .B(p_input[18370]), .Z(n3624) );
  AND U5436 ( .A(p_input[8370]), .B(p_input[38370]), .Z(n3623) );
  AND U5437 ( .A(n3625), .B(n3626), .Z(o[836]) );
  AND U5438 ( .A(p_input[20836]), .B(p_input[10836]), .Z(n3626) );
  AND U5439 ( .A(p_input[836]), .B(p_input[30836]), .Z(n3625) );
  AND U5440 ( .A(n3627), .B(n3628), .Z(o[8369]) );
  AND U5441 ( .A(p_input[28369]), .B(p_input[18369]), .Z(n3628) );
  AND U5442 ( .A(p_input[8369]), .B(p_input[38369]), .Z(n3627) );
  AND U5443 ( .A(n3629), .B(n3630), .Z(o[8368]) );
  AND U5444 ( .A(p_input[28368]), .B(p_input[18368]), .Z(n3630) );
  AND U5445 ( .A(p_input[8368]), .B(p_input[38368]), .Z(n3629) );
  AND U5446 ( .A(n3631), .B(n3632), .Z(o[8367]) );
  AND U5447 ( .A(p_input[28367]), .B(p_input[18367]), .Z(n3632) );
  AND U5448 ( .A(p_input[8367]), .B(p_input[38367]), .Z(n3631) );
  AND U5449 ( .A(n3633), .B(n3634), .Z(o[8366]) );
  AND U5450 ( .A(p_input[28366]), .B(p_input[18366]), .Z(n3634) );
  AND U5451 ( .A(p_input[8366]), .B(p_input[38366]), .Z(n3633) );
  AND U5452 ( .A(n3635), .B(n3636), .Z(o[8365]) );
  AND U5453 ( .A(p_input[28365]), .B(p_input[18365]), .Z(n3636) );
  AND U5454 ( .A(p_input[8365]), .B(p_input[38365]), .Z(n3635) );
  AND U5455 ( .A(n3637), .B(n3638), .Z(o[8364]) );
  AND U5456 ( .A(p_input[28364]), .B(p_input[18364]), .Z(n3638) );
  AND U5457 ( .A(p_input[8364]), .B(p_input[38364]), .Z(n3637) );
  AND U5458 ( .A(n3639), .B(n3640), .Z(o[8363]) );
  AND U5459 ( .A(p_input[28363]), .B(p_input[18363]), .Z(n3640) );
  AND U5460 ( .A(p_input[8363]), .B(p_input[38363]), .Z(n3639) );
  AND U5461 ( .A(n3641), .B(n3642), .Z(o[8362]) );
  AND U5462 ( .A(p_input[28362]), .B(p_input[18362]), .Z(n3642) );
  AND U5463 ( .A(p_input[8362]), .B(p_input[38362]), .Z(n3641) );
  AND U5464 ( .A(n3643), .B(n3644), .Z(o[8361]) );
  AND U5465 ( .A(p_input[28361]), .B(p_input[18361]), .Z(n3644) );
  AND U5466 ( .A(p_input[8361]), .B(p_input[38361]), .Z(n3643) );
  AND U5467 ( .A(n3645), .B(n3646), .Z(o[8360]) );
  AND U5468 ( .A(p_input[28360]), .B(p_input[18360]), .Z(n3646) );
  AND U5469 ( .A(p_input[8360]), .B(p_input[38360]), .Z(n3645) );
  AND U5470 ( .A(n3647), .B(n3648), .Z(o[835]) );
  AND U5471 ( .A(p_input[20835]), .B(p_input[10835]), .Z(n3648) );
  AND U5472 ( .A(p_input[835]), .B(p_input[30835]), .Z(n3647) );
  AND U5473 ( .A(n3649), .B(n3650), .Z(o[8359]) );
  AND U5474 ( .A(p_input[28359]), .B(p_input[18359]), .Z(n3650) );
  AND U5475 ( .A(p_input[8359]), .B(p_input[38359]), .Z(n3649) );
  AND U5476 ( .A(n3651), .B(n3652), .Z(o[8358]) );
  AND U5477 ( .A(p_input[28358]), .B(p_input[18358]), .Z(n3652) );
  AND U5478 ( .A(p_input[8358]), .B(p_input[38358]), .Z(n3651) );
  AND U5479 ( .A(n3653), .B(n3654), .Z(o[8357]) );
  AND U5480 ( .A(p_input[28357]), .B(p_input[18357]), .Z(n3654) );
  AND U5481 ( .A(p_input[8357]), .B(p_input[38357]), .Z(n3653) );
  AND U5482 ( .A(n3655), .B(n3656), .Z(o[8356]) );
  AND U5483 ( .A(p_input[28356]), .B(p_input[18356]), .Z(n3656) );
  AND U5484 ( .A(p_input[8356]), .B(p_input[38356]), .Z(n3655) );
  AND U5485 ( .A(n3657), .B(n3658), .Z(o[8355]) );
  AND U5486 ( .A(p_input[28355]), .B(p_input[18355]), .Z(n3658) );
  AND U5487 ( .A(p_input[8355]), .B(p_input[38355]), .Z(n3657) );
  AND U5488 ( .A(n3659), .B(n3660), .Z(o[8354]) );
  AND U5489 ( .A(p_input[28354]), .B(p_input[18354]), .Z(n3660) );
  AND U5490 ( .A(p_input[8354]), .B(p_input[38354]), .Z(n3659) );
  AND U5491 ( .A(n3661), .B(n3662), .Z(o[8353]) );
  AND U5492 ( .A(p_input[28353]), .B(p_input[18353]), .Z(n3662) );
  AND U5493 ( .A(p_input[8353]), .B(p_input[38353]), .Z(n3661) );
  AND U5494 ( .A(n3663), .B(n3664), .Z(o[8352]) );
  AND U5495 ( .A(p_input[28352]), .B(p_input[18352]), .Z(n3664) );
  AND U5496 ( .A(p_input[8352]), .B(p_input[38352]), .Z(n3663) );
  AND U5497 ( .A(n3665), .B(n3666), .Z(o[8351]) );
  AND U5498 ( .A(p_input[28351]), .B(p_input[18351]), .Z(n3666) );
  AND U5499 ( .A(p_input[8351]), .B(p_input[38351]), .Z(n3665) );
  AND U5500 ( .A(n3667), .B(n3668), .Z(o[8350]) );
  AND U5501 ( .A(p_input[28350]), .B(p_input[18350]), .Z(n3668) );
  AND U5502 ( .A(p_input[8350]), .B(p_input[38350]), .Z(n3667) );
  AND U5503 ( .A(n3669), .B(n3670), .Z(o[834]) );
  AND U5504 ( .A(p_input[20834]), .B(p_input[10834]), .Z(n3670) );
  AND U5505 ( .A(p_input[834]), .B(p_input[30834]), .Z(n3669) );
  AND U5506 ( .A(n3671), .B(n3672), .Z(o[8349]) );
  AND U5507 ( .A(p_input[28349]), .B(p_input[18349]), .Z(n3672) );
  AND U5508 ( .A(p_input[8349]), .B(p_input[38349]), .Z(n3671) );
  AND U5509 ( .A(n3673), .B(n3674), .Z(o[8348]) );
  AND U5510 ( .A(p_input[28348]), .B(p_input[18348]), .Z(n3674) );
  AND U5511 ( .A(p_input[8348]), .B(p_input[38348]), .Z(n3673) );
  AND U5512 ( .A(n3675), .B(n3676), .Z(o[8347]) );
  AND U5513 ( .A(p_input[28347]), .B(p_input[18347]), .Z(n3676) );
  AND U5514 ( .A(p_input[8347]), .B(p_input[38347]), .Z(n3675) );
  AND U5515 ( .A(n3677), .B(n3678), .Z(o[8346]) );
  AND U5516 ( .A(p_input[28346]), .B(p_input[18346]), .Z(n3678) );
  AND U5517 ( .A(p_input[8346]), .B(p_input[38346]), .Z(n3677) );
  AND U5518 ( .A(n3679), .B(n3680), .Z(o[8345]) );
  AND U5519 ( .A(p_input[28345]), .B(p_input[18345]), .Z(n3680) );
  AND U5520 ( .A(p_input[8345]), .B(p_input[38345]), .Z(n3679) );
  AND U5521 ( .A(n3681), .B(n3682), .Z(o[8344]) );
  AND U5522 ( .A(p_input[28344]), .B(p_input[18344]), .Z(n3682) );
  AND U5523 ( .A(p_input[8344]), .B(p_input[38344]), .Z(n3681) );
  AND U5524 ( .A(n3683), .B(n3684), .Z(o[8343]) );
  AND U5525 ( .A(p_input[28343]), .B(p_input[18343]), .Z(n3684) );
  AND U5526 ( .A(p_input[8343]), .B(p_input[38343]), .Z(n3683) );
  AND U5527 ( .A(n3685), .B(n3686), .Z(o[8342]) );
  AND U5528 ( .A(p_input[28342]), .B(p_input[18342]), .Z(n3686) );
  AND U5529 ( .A(p_input[8342]), .B(p_input[38342]), .Z(n3685) );
  AND U5530 ( .A(n3687), .B(n3688), .Z(o[8341]) );
  AND U5531 ( .A(p_input[28341]), .B(p_input[18341]), .Z(n3688) );
  AND U5532 ( .A(p_input[8341]), .B(p_input[38341]), .Z(n3687) );
  AND U5533 ( .A(n3689), .B(n3690), .Z(o[8340]) );
  AND U5534 ( .A(p_input[28340]), .B(p_input[18340]), .Z(n3690) );
  AND U5535 ( .A(p_input[8340]), .B(p_input[38340]), .Z(n3689) );
  AND U5536 ( .A(n3691), .B(n3692), .Z(o[833]) );
  AND U5537 ( .A(p_input[20833]), .B(p_input[10833]), .Z(n3692) );
  AND U5538 ( .A(p_input[833]), .B(p_input[30833]), .Z(n3691) );
  AND U5539 ( .A(n3693), .B(n3694), .Z(o[8339]) );
  AND U5540 ( .A(p_input[28339]), .B(p_input[18339]), .Z(n3694) );
  AND U5541 ( .A(p_input[8339]), .B(p_input[38339]), .Z(n3693) );
  AND U5542 ( .A(n3695), .B(n3696), .Z(o[8338]) );
  AND U5543 ( .A(p_input[28338]), .B(p_input[18338]), .Z(n3696) );
  AND U5544 ( .A(p_input[8338]), .B(p_input[38338]), .Z(n3695) );
  AND U5545 ( .A(n3697), .B(n3698), .Z(o[8337]) );
  AND U5546 ( .A(p_input[28337]), .B(p_input[18337]), .Z(n3698) );
  AND U5547 ( .A(p_input[8337]), .B(p_input[38337]), .Z(n3697) );
  AND U5548 ( .A(n3699), .B(n3700), .Z(o[8336]) );
  AND U5549 ( .A(p_input[28336]), .B(p_input[18336]), .Z(n3700) );
  AND U5550 ( .A(p_input[8336]), .B(p_input[38336]), .Z(n3699) );
  AND U5551 ( .A(n3701), .B(n3702), .Z(o[8335]) );
  AND U5552 ( .A(p_input[28335]), .B(p_input[18335]), .Z(n3702) );
  AND U5553 ( .A(p_input[8335]), .B(p_input[38335]), .Z(n3701) );
  AND U5554 ( .A(n3703), .B(n3704), .Z(o[8334]) );
  AND U5555 ( .A(p_input[28334]), .B(p_input[18334]), .Z(n3704) );
  AND U5556 ( .A(p_input[8334]), .B(p_input[38334]), .Z(n3703) );
  AND U5557 ( .A(n3705), .B(n3706), .Z(o[8333]) );
  AND U5558 ( .A(p_input[28333]), .B(p_input[18333]), .Z(n3706) );
  AND U5559 ( .A(p_input[8333]), .B(p_input[38333]), .Z(n3705) );
  AND U5560 ( .A(n3707), .B(n3708), .Z(o[8332]) );
  AND U5561 ( .A(p_input[28332]), .B(p_input[18332]), .Z(n3708) );
  AND U5562 ( .A(p_input[8332]), .B(p_input[38332]), .Z(n3707) );
  AND U5563 ( .A(n3709), .B(n3710), .Z(o[8331]) );
  AND U5564 ( .A(p_input[28331]), .B(p_input[18331]), .Z(n3710) );
  AND U5565 ( .A(p_input[8331]), .B(p_input[38331]), .Z(n3709) );
  AND U5566 ( .A(n3711), .B(n3712), .Z(o[8330]) );
  AND U5567 ( .A(p_input[28330]), .B(p_input[18330]), .Z(n3712) );
  AND U5568 ( .A(p_input[8330]), .B(p_input[38330]), .Z(n3711) );
  AND U5569 ( .A(n3713), .B(n3714), .Z(o[832]) );
  AND U5570 ( .A(p_input[20832]), .B(p_input[10832]), .Z(n3714) );
  AND U5571 ( .A(p_input[832]), .B(p_input[30832]), .Z(n3713) );
  AND U5572 ( .A(n3715), .B(n3716), .Z(o[8329]) );
  AND U5573 ( .A(p_input[28329]), .B(p_input[18329]), .Z(n3716) );
  AND U5574 ( .A(p_input[8329]), .B(p_input[38329]), .Z(n3715) );
  AND U5575 ( .A(n3717), .B(n3718), .Z(o[8328]) );
  AND U5576 ( .A(p_input[28328]), .B(p_input[18328]), .Z(n3718) );
  AND U5577 ( .A(p_input[8328]), .B(p_input[38328]), .Z(n3717) );
  AND U5578 ( .A(n3719), .B(n3720), .Z(o[8327]) );
  AND U5579 ( .A(p_input[28327]), .B(p_input[18327]), .Z(n3720) );
  AND U5580 ( .A(p_input[8327]), .B(p_input[38327]), .Z(n3719) );
  AND U5581 ( .A(n3721), .B(n3722), .Z(o[8326]) );
  AND U5582 ( .A(p_input[28326]), .B(p_input[18326]), .Z(n3722) );
  AND U5583 ( .A(p_input[8326]), .B(p_input[38326]), .Z(n3721) );
  AND U5584 ( .A(n3723), .B(n3724), .Z(o[8325]) );
  AND U5585 ( .A(p_input[28325]), .B(p_input[18325]), .Z(n3724) );
  AND U5586 ( .A(p_input[8325]), .B(p_input[38325]), .Z(n3723) );
  AND U5587 ( .A(n3725), .B(n3726), .Z(o[8324]) );
  AND U5588 ( .A(p_input[28324]), .B(p_input[18324]), .Z(n3726) );
  AND U5589 ( .A(p_input[8324]), .B(p_input[38324]), .Z(n3725) );
  AND U5590 ( .A(n3727), .B(n3728), .Z(o[8323]) );
  AND U5591 ( .A(p_input[28323]), .B(p_input[18323]), .Z(n3728) );
  AND U5592 ( .A(p_input[8323]), .B(p_input[38323]), .Z(n3727) );
  AND U5593 ( .A(n3729), .B(n3730), .Z(o[8322]) );
  AND U5594 ( .A(p_input[28322]), .B(p_input[18322]), .Z(n3730) );
  AND U5595 ( .A(p_input[8322]), .B(p_input[38322]), .Z(n3729) );
  AND U5596 ( .A(n3731), .B(n3732), .Z(o[8321]) );
  AND U5597 ( .A(p_input[28321]), .B(p_input[18321]), .Z(n3732) );
  AND U5598 ( .A(p_input[8321]), .B(p_input[38321]), .Z(n3731) );
  AND U5599 ( .A(n3733), .B(n3734), .Z(o[8320]) );
  AND U5600 ( .A(p_input[28320]), .B(p_input[18320]), .Z(n3734) );
  AND U5601 ( .A(p_input[8320]), .B(p_input[38320]), .Z(n3733) );
  AND U5602 ( .A(n3735), .B(n3736), .Z(o[831]) );
  AND U5603 ( .A(p_input[20831]), .B(p_input[10831]), .Z(n3736) );
  AND U5604 ( .A(p_input[831]), .B(p_input[30831]), .Z(n3735) );
  AND U5605 ( .A(n3737), .B(n3738), .Z(o[8319]) );
  AND U5606 ( .A(p_input[28319]), .B(p_input[18319]), .Z(n3738) );
  AND U5607 ( .A(p_input[8319]), .B(p_input[38319]), .Z(n3737) );
  AND U5608 ( .A(n3739), .B(n3740), .Z(o[8318]) );
  AND U5609 ( .A(p_input[28318]), .B(p_input[18318]), .Z(n3740) );
  AND U5610 ( .A(p_input[8318]), .B(p_input[38318]), .Z(n3739) );
  AND U5611 ( .A(n3741), .B(n3742), .Z(o[8317]) );
  AND U5612 ( .A(p_input[28317]), .B(p_input[18317]), .Z(n3742) );
  AND U5613 ( .A(p_input[8317]), .B(p_input[38317]), .Z(n3741) );
  AND U5614 ( .A(n3743), .B(n3744), .Z(o[8316]) );
  AND U5615 ( .A(p_input[28316]), .B(p_input[18316]), .Z(n3744) );
  AND U5616 ( .A(p_input[8316]), .B(p_input[38316]), .Z(n3743) );
  AND U5617 ( .A(n3745), .B(n3746), .Z(o[8315]) );
  AND U5618 ( .A(p_input[28315]), .B(p_input[18315]), .Z(n3746) );
  AND U5619 ( .A(p_input[8315]), .B(p_input[38315]), .Z(n3745) );
  AND U5620 ( .A(n3747), .B(n3748), .Z(o[8314]) );
  AND U5621 ( .A(p_input[28314]), .B(p_input[18314]), .Z(n3748) );
  AND U5622 ( .A(p_input[8314]), .B(p_input[38314]), .Z(n3747) );
  AND U5623 ( .A(n3749), .B(n3750), .Z(o[8313]) );
  AND U5624 ( .A(p_input[28313]), .B(p_input[18313]), .Z(n3750) );
  AND U5625 ( .A(p_input[8313]), .B(p_input[38313]), .Z(n3749) );
  AND U5626 ( .A(n3751), .B(n3752), .Z(o[8312]) );
  AND U5627 ( .A(p_input[28312]), .B(p_input[18312]), .Z(n3752) );
  AND U5628 ( .A(p_input[8312]), .B(p_input[38312]), .Z(n3751) );
  AND U5629 ( .A(n3753), .B(n3754), .Z(o[8311]) );
  AND U5630 ( .A(p_input[28311]), .B(p_input[18311]), .Z(n3754) );
  AND U5631 ( .A(p_input[8311]), .B(p_input[38311]), .Z(n3753) );
  AND U5632 ( .A(n3755), .B(n3756), .Z(o[8310]) );
  AND U5633 ( .A(p_input[28310]), .B(p_input[18310]), .Z(n3756) );
  AND U5634 ( .A(p_input[8310]), .B(p_input[38310]), .Z(n3755) );
  AND U5635 ( .A(n3757), .B(n3758), .Z(o[830]) );
  AND U5636 ( .A(p_input[20830]), .B(p_input[10830]), .Z(n3758) );
  AND U5637 ( .A(p_input[830]), .B(p_input[30830]), .Z(n3757) );
  AND U5638 ( .A(n3759), .B(n3760), .Z(o[8309]) );
  AND U5639 ( .A(p_input[28309]), .B(p_input[18309]), .Z(n3760) );
  AND U5640 ( .A(p_input[8309]), .B(p_input[38309]), .Z(n3759) );
  AND U5641 ( .A(n3761), .B(n3762), .Z(o[8308]) );
  AND U5642 ( .A(p_input[28308]), .B(p_input[18308]), .Z(n3762) );
  AND U5643 ( .A(p_input[8308]), .B(p_input[38308]), .Z(n3761) );
  AND U5644 ( .A(n3763), .B(n3764), .Z(o[8307]) );
  AND U5645 ( .A(p_input[28307]), .B(p_input[18307]), .Z(n3764) );
  AND U5646 ( .A(p_input[8307]), .B(p_input[38307]), .Z(n3763) );
  AND U5647 ( .A(n3765), .B(n3766), .Z(o[8306]) );
  AND U5648 ( .A(p_input[28306]), .B(p_input[18306]), .Z(n3766) );
  AND U5649 ( .A(p_input[8306]), .B(p_input[38306]), .Z(n3765) );
  AND U5650 ( .A(n3767), .B(n3768), .Z(o[8305]) );
  AND U5651 ( .A(p_input[28305]), .B(p_input[18305]), .Z(n3768) );
  AND U5652 ( .A(p_input[8305]), .B(p_input[38305]), .Z(n3767) );
  AND U5653 ( .A(n3769), .B(n3770), .Z(o[8304]) );
  AND U5654 ( .A(p_input[28304]), .B(p_input[18304]), .Z(n3770) );
  AND U5655 ( .A(p_input[8304]), .B(p_input[38304]), .Z(n3769) );
  AND U5656 ( .A(n3771), .B(n3772), .Z(o[8303]) );
  AND U5657 ( .A(p_input[28303]), .B(p_input[18303]), .Z(n3772) );
  AND U5658 ( .A(p_input[8303]), .B(p_input[38303]), .Z(n3771) );
  AND U5659 ( .A(n3773), .B(n3774), .Z(o[8302]) );
  AND U5660 ( .A(p_input[28302]), .B(p_input[18302]), .Z(n3774) );
  AND U5661 ( .A(p_input[8302]), .B(p_input[38302]), .Z(n3773) );
  AND U5662 ( .A(n3775), .B(n3776), .Z(o[8301]) );
  AND U5663 ( .A(p_input[28301]), .B(p_input[18301]), .Z(n3776) );
  AND U5664 ( .A(p_input[8301]), .B(p_input[38301]), .Z(n3775) );
  AND U5665 ( .A(n3777), .B(n3778), .Z(o[8300]) );
  AND U5666 ( .A(p_input[28300]), .B(p_input[18300]), .Z(n3778) );
  AND U5667 ( .A(p_input[8300]), .B(p_input[38300]), .Z(n3777) );
  AND U5668 ( .A(n3779), .B(n3780), .Z(o[82]) );
  AND U5669 ( .A(p_input[20082]), .B(p_input[10082]), .Z(n3780) );
  AND U5670 ( .A(p_input[82]), .B(p_input[30082]), .Z(n3779) );
  AND U5671 ( .A(n3781), .B(n3782), .Z(o[829]) );
  AND U5672 ( .A(p_input[20829]), .B(p_input[10829]), .Z(n3782) );
  AND U5673 ( .A(p_input[829]), .B(p_input[30829]), .Z(n3781) );
  AND U5674 ( .A(n3783), .B(n3784), .Z(o[8299]) );
  AND U5675 ( .A(p_input[28299]), .B(p_input[18299]), .Z(n3784) );
  AND U5676 ( .A(p_input[8299]), .B(p_input[38299]), .Z(n3783) );
  AND U5677 ( .A(n3785), .B(n3786), .Z(o[8298]) );
  AND U5678 ( .A(p_input[28298]), .B(p_input[18298]), .Z(n3786) );
  AND U5679 ( .A(p_input[8298]), .B(p_input[38298]), .Z(n3785) );
  AND U5680 ( .A(n3787), .B(n3788), .Z(o[8297]) );
  AND U5681 ( .A(p_input[28297]), .B(p_input[18297]), .Z(n3788) );
  AND U5682 ( .A(p_input[8297]), .B(p_input[38297]), .Z(n3787) );
  AND U5683 ( .A(n3789), .B(n3790), .Z(o[8296]) );
  AND U5684 ( .A(p_input[28296]), .B(p_input[18296]), .Z(n3790) );
  AND U5685 ( .A(p_input[8296]), .B(p_input[38296]), .Z(n3789) );
  AND U5686 ( .A(n3791), .B(n3792), .Z(o[8295]) );
  AND U5687 ( .A(p_input[28295]), .B(p_input[18295]), .Z(n3792) );
  AND U5688 ( .A(p_input[8295]), .B(p_input[38295]), .Z(n3791) );
  AND U5689 ( .A(n3793), .B(n3794), .Z(o[8294]) );
  AND U5690 ( .A(p_input[28294]), .B(p_input[18294]), .Z(n3794) );
  AND U5691 ( .A(p_input[8294]), .B(p_input[38294]), .Z(n3793) );
  AND U5692 ( .A(n3795), .B(n3796), .Z(o[8293]) );
  AND U5693 ( .A(p_input[28293]), .B(p_input[18293]), .Z(n3796) );
  AND U5694 ( .A(p_input[8293]), .B(p_input[38293]), .Z(n3795) );
  AND U5695 ( .A(n3797), .B(n3798), .Z(o[8292]) );
  AND U5696 ( .A(p_input[28292]), .B(p_input[18292]), .Z(n3798) );
  AND U5697 ( .A(p_input[8292]), .B(p_input[38292]), .Z(n3797) );
  AND U5698 ( .A(n3799), .B(n3800), .Z(o[8291]) );
  AND U5699 ( .A(p_input[28291]), .B(p_input[18291]), .Z(n3800) );
  AND U5700 ( .A(p_input[8291]), .B(p_input[38291]), .Z(n3799) );
  AND U5701 ( .A(n3801), .B(n3802), .Z(o[8290]) );
  AND U5702 ( .A(p_input[28290]), .B(p_input[18290]), .Z(n3802) );
  AND U5703 ( .A(p_input[8290]), .B(p_input[38290]), .Z(n3801) );
  AND U5704 ( .A(n3803), .B(n3804), .Z(o[828]) );
  AND U5705 ( .A(p_input[20828]), .B(p_input[10828]), .Z(n3804) );
  AND U5706 ( .A(p_input[828]), .B(p_input[30828]), .Z(n3803) );
  AND U5707 ( .A(n3805), .B(n3806), .Z(o[8289]) );
  AND U5708 ( .A(p_input[28289]), .B(p_input[18289]), .Z(n3806) );
  AND U5709 ( .A(p_input[8289]), .B(p_input[38289]), .Z(n3805) );
  AND U5710 ( .A(n3807), .B(n3808), .Z(o[8288]) );
  AND U5711 ( .A(p_input[28288]), .B(p_input[18288]), .Z(n3808) );
  AND U5712 ( .A(p_input[8288]), .B(p_input[38288]), .Z(n3807) );
  AND U5713 ( .A(n3809), .B(n3810), .Z(o[8287]) );
  AND U5714 ( .A(p_input[28287]), .B(p_input[18287]), .Z(n3810) );
  AND U5715 ( .A(p_input[8287]), .B(p_input[38287]), .Z(n3809) );
  AND U5716 ( .A(n3811), .B(n3812), .Z(o[8286]) );
  AND U5717 ( .A(p_input[28286]), .B(p_input[18286]), .Z(n3812) );
  AND U5718 ( .A(p_input[8286]), .B(p_input[38286]), .Z(n3811) );
  AND U5719 ( .A(n3813), .B(n3814), .Z(o[8285]) );
  AND U5720 ( .A(p_input[28285]), .B(p_input[18285]), .Z(n3814) );
  AND U5721 ( .A(p_input[8285]), .B(p_input[38285]), .Z(n3813) );
  AND U5722 ( .A(n3815), .B(n3816), .Z(o[8284]) );
  AND U5723 ( .A(p_input[28284]), .B(p_input[18284]), .Z(n3816) );
  AND U5724 ( .A(p_input[8284]), .B(p_input[38284]), .Z(n3815) );
  AND U5725 ( .A(n3817), .B(n3818), .Z(o[8283]) );
  AND U5726 ( .A(p_input[28283]), .B(p_input[18283]), .Z(n3818) );
  AND U5727 ( .A(p_input[8283]), .B(p_input[38283]), .Z(n3817) );
  AND U5728 ( .A(n3819), .B(n3820), .Z(o[8282]) );
  AND U5729 ( .A(p_input[28282]), .B(p_input[18282]), .Z(n3820) );
  AND U5730 ( .A(p_input[8282]), .B(p_input[38282]), .Z(n3819) );
  AND U5731 ( .A(n3821), .B(n3822), .Z(o[8281]) );
  AND U5732 ( .A(p_input[28281]), .B(p_input[18281]), .Z(n3822) );
  AND U5733 ( .A(p_input[8281]), .B(p_input[38281]), .Z(n3821) );
  AND U5734 ( .A(n3823), .B(n3824), .Z(o[8280]) );
  AND U5735 ( .A(p_input[28280]), .B(p_input[18280]), .Z(n3824) );
  AND U5736 ( .A(p_input[8280]), .B(p_input[38280]), .Z(n3823) );
  AND U5737 ( .A(n3825), .B(n3826), .Z(o[827]) );
  AND U5738 ( .A(p_input[20827]), .B(p_input[10827]), .Z(n3826) );
  AND U5739 ( .A(p_input[827]), .B(p_input[30827]), .Z(n3825) );
  AND U5740 ( .A(n3827), .B(n3828), .Z(o[8279]) );
  AND U5741 ( .A(p_input[28279]), .B(p_input[18279]), .Z(n3828) );
  AND U5742 ( .A(p_input[8279]), .B(p_input[38279]), .Z(n3827) );
  AND U5743 ( .A(n3829), .B(n3830), .Z(o[8278]) );
  AND U5744 ( .A(p_input[28278]), .B(p_input[18278]), .Z(n3830) );
  AND U5745 ( .A(p_input[8278]), .B(p_input[38278]), .Z(n3829) );
  AND U5746 ( .A(n3831), .B(n3832), .Z(o[8277]) );
  AND U5747 ( .A(p_input[28277]), .B(p_input[18277]), .Z(n3832) );
  AND U5748 ( .A(p_input[8277]), .B(p_input[38277]), .Z(n3831) );
  AND U5749 ( .A(n3833), .B(n3834), .Z(o[8276]) );
  AND U5750 ( .A(p_input[28276]), .B(p_input[18276]), .Z(n3834) );
  AND U5751 ( .A(p_input[8276]), .B(p_input[38276]), .Z(n3833) );
  AND U5752 ( .A(n3835), .B(n3836), .Z(o[8275]) );
  AND U5753 ( .A(p_input[28275]), .B(p_input[18275]), .Z(n3836) );
  AND U5754 ( .A(p_input[8275]), .B(p_input[38275]), .Z(n3835) );
  AND U5755 ( .A(n3837), .B(n3838), .Z(o[8274]) );
  AND U5756 ( .A(p_input[28274]), .B(p_input[18274]), .Z(n3838) );
  AND U5757 ( .A(p_input[8274]), .B(p_input[38274]), .Z(n3837) );
  AND U5758 ( .A(n3839), .B(n3840), .Z(o[8273]) );
  AND U5759 ( .A(p_input[28273]), .B(p_input[18273]), .Z(n3840) );
  AND U5760 ( .A(p_input[8273]), .B(p_input[38273]), .Z(n3839) );
  AND U5761 ( .A(n3841), .B(n3842), .Z(o[8272]) );
  AND U5762 ( .A(p_input[28272]), .B(p_input[18272]), .Z(n3842) );
  AND U5763 ( .A(p_input[8272]), .B(p_input[38272]), .Z(n3841) );
  AND U5764 ( .A(n3843), .B(n3844), .Z(o[8271]) );
  AND U5765 ( .A(p_input[28271]), .B(p_input[18271]), .Z(n3844) );
  AND U5766 ( .A(p_input[8271]), .B(p_input[38271]), .Z(n3843) );
  AND U5767 ( .A(n3845), .B(n3846), .Z(o[8270]) );
  AND U5768 ( .A(p_input[28270]), .B(p_input[18270]), .Z(n3846) );
  AND U5769 ( .A(p_input[8270]), .B(p_input[38270]), .Z(n3845) );
  AND U5770 ( .A(n3847), .B(n3848), .Z(o[826]) );
  AND U5771 ( .A(p_input[20826]), .B(p_input[10826]), .Z(n3848) );
  AND U5772 ( .A(p_input[826]), .B(p_input[30826]), .Z(n3847) );
  AND U5773 ( .A(n3849), .B(n3850), .Z(o[8269]) );
  AND U5774 ( .A(p_input[28269]), .B(p_input[18269]), .Z(n3850) );
  AND U5775 ( .A(p_input[8269]), .B(p_input[38269]), .Z(n3849) );
  AND U5776 ( .A(n3851), .B(n3852), .Z(o[8268]) );
  AND U5777 ( .A(p_input[28268]), .B(p_input[18268]), .Z(n3852) );
  AND U5778 ( .A(p_input[8268]), .B(p_input[38268]), .Z(n3851) );
  AND U5779 ( .A(n3853), .B(n3854), .Z(o[8267]) );
  AND U5780 ( .A(p_input[28267]), .B(p_input[18267]), .Z(n3854) );
  AND U5781 ( .A(p_input[8267]), .B(p_input[38267]), .Z(n3853) );
  AND U5782 ( .A(n3855), .B(n3856), .Z(o[8266]) );
  AND U5783 ( .A(p_input[28266]), .B(p_input[18266]), .Z(n3856) );
  AND U5784 ( .A(p_input[8266]), .B(p_input[38266]), .Z(n3855) );
  AND U5785 ( .A(n3857), .B(n3858), .Z(o[8265]) );
  AND U5786 ( .A(p_input[28265]), .B(p_input[18265]), .Z(n3858) );
  AND U5787 ( .A(p_input[8265]), .B(p_input[38265]), .Z(n3857) );
  AND U5788 ( .A(n3859), .B(n3860), .Z(o[8264]) );
  AND U5789 ( .A(p_input[28264]), .B(p_input[18264]), .Z(n3860) );
  AND U5790 ( .A(p_input[8264]), .B(p_input[38264]), .Z(n3859) );
  AND U5791 ( .A(n3861), .B(n3862), .Z(o[8263]) );
  AND U5792 ( .A(p_input[28263]), .B(p_input[18263]), .Z(n3862) );
  AND U5793 ( .A(p_input[8263]), .B(p_input[38263]), .Z(n3861) );
  AND U5794 ( .A(n3863), .B(n3864), .Z(o[8262]) );
  AND U5795 ( .A(p_input[28262]), .B(p_input[18262]), .Z(n3864) );
  AND U5796 ( .A(p_input[8262]), .B(p_input[38262]), .Z(n3863) );
  AND U5797 ( .A(n3865), .B(n3866), .Z(o[8261]) );
  AND U5798 ( .A(p_input[28261]), .B(p_input[18261]), .Z(n3866) );
  AND U5799 ( .A(p_input[8261]), .B(p_input[38261]), .Z(n3865) );
  AND U5800 ( .A(n3867), .B(n3868), .Z(o[8260]) );
  AND U5801 ( .A(p_input[28260]), .B(p_input[18260]), .Z(n3868) );
  AND U5802 ( .A(p_input[8260]), .B(p_input[38260]), .Z(n3867) );
  AND U5803 ( .A(n3869), .B(n3870), .Z(o[825]) );
  AND U5804 ( .A(p_input[20825]), .B(p_input[10825]), .Z(n3870) );
  AND U5805 ( .A(p_input[825]), .B(p_input[30825]), .Z(n3869) );
  AND U5806 ( .A(n3871), .B(n3872), .Z(o[8259]) );
  AND U5807 ( .A(p_input[28259]), .B(p_input[18259]), .Z(n3872) );
  AND U5808 ( .A(p_input[8259]), .B(p_input[38259]), .Z(n3871) );
  AND U5809 ( .A(n3873), .B(n3874), .Z(o[8258]) );
  AND U5810 ( .A(p_input[28258]), .B(p_input[18258]), .Z(n3874) );
  AND U5811 ( .A(p_input[8258]), .B(p_input[38258]), .Z(n3873) );
  AND U5812 ( .A(n3875), .B(n3876), .Z(o[8257]) );
  AND U5813 ( .A(p_input[28257]), .B(p_input[18257]), .Z(n3876) );
  AND U5814 ( .A(p_input[8257]), .B(p_input[38257]), .Z(n3875) );
  AND U5815 ( .A(n3877), .B(n3878), .Z(o[8256]) );
  AND U5816 ( .A(p_input[28256]), .B(p_input[18256]), .Z(n3878) );
  AND U5817 ( .A(p_input[8256]), .B(p_input[38256]), .Z(n3877) );
  AND U5818 ( .A(n3879), .B(n3880), .Z(o[8255]) );
  AND U5819 ( .A(p_input[28255]), .B(p_input[18255]), .Z(n3880) );
  AND U5820 ( .A(p_input[8255]), .B(p_input[38255]), .Z(n3879) );
  AND U5821 ( .A(n3881), .B(n3882), .Z(o[8254]) );
  AND U5822 ( .A(p_input[28254]), .B(p_input[18254]), .Z(n3882) );
  AND U5823 ( .A(p_input[8254]), .B(p_input[38254]), .Z(n3881) );
  AND U5824 ( .A(n3883), .B(n3884), .Z(o[8253]) );
  AND U5825 ( .A(p_input[28253]), .B(p_input[18253]), .Z(n3884) );
  AND U5826 ( .A(p_input[8253]), .B(p_input[38253]), .Z(n3883) );
  AND U5827 ( .A(n3885), .B(n3886), .Z(o[8252]) );
  AND U5828 ( .A(p_input[28252]), .B(p_input[18252]), .Z(n3886) );
  AND U5829 ( .A(p_input[8252]), .B(p_input[38252]), .Z(n3885) );
  AND U5830 ( .A(n3887), .B(n3888), .Z(o[8251]) );
  AND U5831 ( .A(p_input[28251]), .B(p_input[18251]), .Z(n3888) );
  AND U5832 ( .A(p_input[8251]), .B(p_input[38251]), .Z(n3887) );
  AND U5833 ( .A(n3889), .B(n3890), .Z(o[8250]) );
  AND U5834 ( .A(p_input[28250]), .B(p_input[18250]), .Z(n3890) );
  AND U5835 ( .A(p_input[8250]), .B(p_input[38250]), .Z(n3889) );
  AND U5836 ( .A(n3891), .B(n3892), .Z(o[824]) );
  AND U5837 ( .A(p_input[20824]), .B(p_input[10824]), .Z(n3892) );
  AND U5838 ( .A(p_input[824]), .B(p_input[30824]), .Z(n3891) );
  AND U5839 ( .A(n3893), .B(n3894), .Z(o[8249]) );
  AND U5840 ( .A(p_input[28249]), .B(p_input[18249]), .Z(n3894) );
  AND U5841 ( .A(p_input[8249]), .B(p_input[38249]), .Z(n3893) );
  AND U5842 ( .A(n3895), .B(n3896), .Z(o[8248]) );
  AND U5843 ( .A(p_input[28248]), .B(p_input[18248]), .Z(n3896) );
  AND U5844 ( .A(p_input[8248]), .B(p_input[38248]), .Z(n3895) );
  AND U5845 ( .A(n3897), .B(n3898), .Z(o[8247]) );
  AND U5846 ( .A(p_input[28247]), .B(p_input[18247]), .Z(n3898) );
  AND U5847 ( .A(p_input[8247]), .B(p_input[38247]), .Z(n3897) );
  AND U5848 ( .A(n3899), .B(n3900), .Z(o[8246]) );
  AND U5849 ( .A(p_input[28246]), .B(p_input[18246]), .Z(n3900) );
  AND U5850 ( .A(p_input[8246]), .B(p_input[38246]), .Z(n3899) );
  AND U5851 ( .A(n3901), .B(n3902), .Z(o[8245]) );
  AND U5852 ( .A(p_input[28245]), .B(p_input[18245]), .Z(n3902) );
  AND U5853 ( .A(p_input[8245]), .B(p_input[38245]), .Z(n3901) );
  AND U5854 ( .A(n3903), .B(n3904), .Z(o[8244]) );
  AND U5855 ( .A(p_input[28244]), .B(p_input[18244]), .Z(n3904) );
  AND U5856 ( .A(p_input[8244]), .B(p_input[38244]), .Z(n3903) );
  AND U5857 ( .A(n3905), .B(n3906), .Z(o[8243]) );
  AND U5858 ( .A(p_input[28243]), .B(p_input[18243]), .Z(n3906) );
  AND U5859 ( .A(p_input[8243]), .B(p_input[38243]), .Z(n3905) );
  AND U5860 ( .A(n3907), .B(n3908), .Z(o[8242]) );
  AND U5861 ( .A(p_input[28242]), .B(p_input[18242]), .Z(n3908) );
  AND U5862 ( .A(p_input[8242]), .B(p_input[38242]), .Z(n3907) );
  AND U5863 ( .A(n3909), .B(n3910), .Z(o[8241]) );
  AND U5864 ( .A(p_input[28241]), .B(p_input[18241]), .Z(n3910) );
  AND U5865 ( .A(p_input[8241]), .B(p_input[38241]), .Z(n3909) );
  AND U5866 ( .A(n3911), .B(n3912), .Z(o[8240]) );
  AND U5867 ( .A(p_input[28240]), .B(p_input[18240]), .Z(n3912) );
  AND U5868 ( .A(p_input[8240]), .B(p_input[38240]), .Z(n3911) );
  AND U5869 ( .A(n3913), .B(n3914), .Z(o[823]) );
  AND U5870 ( .A(p_input[20823]), .B(p_input[10823]), .Z(n3914) );
  AND U5871 ( .A(p_input[823]), .B(p_input[30823]), .Z(n3913) );
  AND U5872 ( .A(n3915), .B(n3916), .Z(o[8239]) );
  AND U5873 ( .A(p_input[28239]), .B(p_input[18239]), .Z(n3916) );
  AND U5874 ( .A(p_input[8239]), .B(p_input[38239]), .Z(n3915) );
  AND U5875 ( .A(n3917), .B(n3918), .Z(o[8238]) );
  AND U5876 ( .A(p_input[28238]), .B(p_input[18238]), .Z(n3918) );
  AND U5877 ( .A(p_input[8238]), .B(p_input[38238]), .Z(n3917) );
  AND U5878 ( .A(n3919), .B(n3920), .Z(o[8237]) );
  AND U5879 ( .A(p_input[28237]), .B(p_input[18237]), .Z(n3920) );
  AND U5880 ( .A(p_input[8237]), .B(p_input[38237]), .Z(n3919) );
  AND U5881 ( .A(n3921), .B(n3922), .Z(o[8236]) );
  AND U5882 ( .A(p_input[28236]), .B(p_input[18236]), .Z(n3922) );
  AND U5883 ( .A(p_input[8236]), .B(p_input[38236]), .Z(n3921) );
  AND U5884 ( .A(n3923), .B(n3924), .Z(o[8235]) );
  AND U5885 ( .A(p_input[28235]), .B(p_input[18235]), .Z(n3924) );
  AND U5886 ( .A(p_input[8235]), .B(p_input[38235]), .Z(n3923) );
  AND U5887 ( .A(n3925), .B(n3926), .Z(o[8234]) );
  AND U5888 ( .A(p_input[28234]), .B(p_input[18234]), .Z(n3926) );
  AND U5889 ( .A(p_input[8234]), .B(p_input[38234]), .Z(n3925) );
  AND U5890 ( .A(n3927), .B(n3928), .Z(o[8233]) );
  AND U5891 ( .A(p_input[28233]), .B(p_input[18233]), .Z(n3928) );
  AND U5892 ( .A(p_input[8233]), .B(p_input[38233]), .Z(n3927) );
  AND U5893 ( .A(n3929), .B(n3930), .Z(o[8232]) );
  AND U5894 ( .A(p_input[28232]), .B(p_input[18232]), .Z(n3930) );
  AND U5895 ( .A(p_input[8232]), .B(p_input[38232]), .Z(n3929) );
  AND U5896 ( .A(n3931), .B(n3932), .Z(o[8231]) );
  AND U5897 ( .A(p_input[28231]), .B(p_input[18231]), .Z(n3932) );
  AND U5898 ( .A(p_input[8231]), .B(p_input[38231]), .Z(n3931) );
  AND U5899 ( .A(n3933), .B(n3934), .Z(o[8230]) );
  AND U5900 ( .A(p_input[28230]), .B(p_input[18230]), .Z(n3934) );
  AND U5901 ( .A(p_input[8230]), .B(p_input[38230]), .Z(n3933) );
  AND U5902 ( .A(n3935), .B(n3936), .Z(o[822]) );
  AND U5903 ( .A(p_input[20822]), .B(p_input[10822]), .Z(n3936) );
  AND U5904 ( .A(p_input[822]), .B(p_input[30822]), .Z(n3935) );
  AND U5905 ( .A(n3937), .B(n3938), .Z(o[8229]) );
  AND U5906 ( .A(p_input[28229]), .B(p_input[18229]), .Z(n3938) );
  AND U5907 ( .A(p_input[8229]), .B(p_input[38229]), .Z(n3937) );
  AND U5908 ( .A(n3939), .B(n3940), .Z(o[8228]) );
  AND U5909 ( .A(p_input[28228]), .B(p_input[18228]), .Z(n3940) );
  AND U5910 ( .A(p_input[8228]), .B(p_input[38228]), .Z(n3939) );
  AND U5911 ( .A(n3941), .B(n3942), .Z(o[8227]) );
  AND U5912 ( .A(p_input[28227]), .B(p_input[18227]), .Z(n3942) );
  AND U5913 ( .A(p_input[8227]), .B(p_input[38227]), .Z(n3941) );
  AND U5914 ( .A(n3943), .B(n3944), .Z(o[8226]) );
  AND U5915 ( .A(p_input[28226]), .B(p_input[18226]), .Z(n3944) );
  AND U5916 ( .A(p_input[8226]), .B(p_input[38226]), .Z(n3943) );
  AND U5917 ( .A(n3945), .B(n3946), .Z(o[8225]) );
  AND U5918 ( .A(p_input[28225]), .B(p_input[18225]), .Z(n3946) );
  AND U5919 ( .A(p_input[8225]), .B(p_input[38225]), .Z(n3945) );
  AND U5920 ( .A(n3947), .B(n3948), .Z(o[8224]) );
  AND U5921 ( .A(p_input[28224]), .B(p_input[18224]), .Z(n3948) );
  AND U5922 ( .A(p_input[8224]), .B(p_input[38224]), .Z(n3947) );
  AND U5923 ( .A(n3949), .B(n3950), .Z(o[8223]) );
  AND U5924 ( .A(p_input[28223]), .B(p_input[18223]), .Z(n3950) );
  AND U5925 ( .A(p_input[8223]), .B(p_input[38223]), .Z(n3949) );
  AND U5926 ( .A(n3951), .B(n3952), .Z(o[8222]) );
  AND U5927 ( .A(p_input[28222]), .B(p_input[18222]), .Z(n3952) );
  AND U5928 ( .A(p_input[8222]), .B(p_input[38222]), .Z(n3951) );
  AND U5929 ( .A(n3953), .B(n3954), .Z(o[8221]) );
  AND U5930 ( .A(p_input[28221]), .B(p_input[18221]), .Z(n3954) );
  AND U5931 ( .A(p_input[8221]), .B(p_input[38221]), .Z(n3953) );
  AND U5932 ( .A(n3955), .B(n3956), .Z(o[8220]) );
  AND U5933 ( .A(p_input[28220]), .B(p_input[18220]), .Z(n3956) );
  AND U5934 ( .A(p_input[8220]), .B(p_input[38220]), .Z(n3955) );
  AND U5935 ( .A(n3957), .B(n3958), .Z(o[821]) );
  AND U5936 ( .A(p_input[20821]), .B(p_input[10821]), .Z(n3958) );
  AND U5937 ( .A(p_input[821]), .B(p_input[30821]), .Z(n3957) );
  AND U5938 ( .A(n3959), .B(n3960), .Z(o[8219]) );
  AND U5939 ( .A(p_input[28219]), .B(p_input[18219]), .Z(n3960) );
  AND U5940 ( .A(p_input[8219]), .B(p_input[38219]), .Z(n3959) );
  AND U5941 ( .A(n3961), .B(n3962), .Z(o[8218]) );
  AND U5942 ( .A(p_input[28218]), .B(p_input[18218]), .Z(n3962) );
  AND U5943 ( .A(p_input[8218]), .B(p_input[38218]), .Z(n3961) );
  AND U5944 ( .A(n3963), .B(n3964), .Z(o[8217]) );
  AND U5945 ( .A(p_input[28217]), .B(p_input[18217]), .Z(n3964) );
  AND U5946 ( .A(p_input[8217]), .B(p_input[38217]), .Z(n3963) );
  AND U5947 ( .A(n3965), .B(n3966), .Z(o[8216]) );
  AND U5948 ( .A(p_input[28216]), .B(p_input[18216]), .Z(n3966) );
  AND U5949 ( .A(p_input[8216]), .B(p_input[38216]), .Z(n3965) );
  AND U5950 ( .A(n3967), .B(n3968), .Z(o[8215]) );
  AND U5951 ( .A(p_input[28215]), .B(p_input[18215]), .Z(n3968) );
  AND U5952 ( .A(p_input[8215]), .B(p_input[38215]), .Z(n3967) );
  AND U5953 ( .A(n3969), .B(n3970), .Z(o[8214]) );
  AND U5954 ( .A(p_input[28214]), .B(p_input[18214]), .Z(n3970) );
  AND U5955 ( .A(p_input[8214]), .B(p_input[38214]), .Z(n3969) );
  AND U5956 ( .A(n3971), .B(n3972), .Z(o[8213]) );
  AND U5957 ( .A(p_input[28213]), .B(p_input[18213]), .Z(n3972) );
  AND U5958 ( .A(p_input[8213]), .B(p_input[38213]), .Z(n3971) );
  AND U5959 ( .A(n3973), .B(n3974), .Z(o[8212]) );
  AND U5960 ( .A(p_input[28212]), .B(p_input[18212]), .Z(n3974) );
  AND U5961 ( .A(p_input[8212]), .B(p_input[38212]), .Z(n3973) );
  AND U5962 ( .A(n3975), .B(n3976), .Z(o[8211]) );
  AND U5963 ( .A(p_input[28211]), .B(p_input[18211]), .Z(n3976) );
  AND U5964 ( .A(p_input[8211]), .B(p_input[38211]), .Z(n3975) );
  AND U5965 ( .A(n3977), .B(n3978), .Z(o[8210]) );
  AND U5966 ( .A(p_input[28210]), .B(p_input[18210]), .Z(n3978) );
  AND U5967 ( .A(p_input[8210]), .B(p_input[38210]), .Z(n3977) );
  AND U5968 ( .A(n3979), .B(n3980), .Z(o[820]) );
  AND U5969 ( .A(p_input[20820]), .B(p_input[10820]), .Z(n3980) );
  AND U5970 ( .A(p_input[820]), .B(p_input[30820]), .Z(n3979) );
  AND U5971 ( .A(n3981), .B(n3982), .Z(o[8209]) );
  AND U5972 ( .A(p_input[28209]), .B(p_input[18209]), .Z(n3982) );
  AND U5973 ( .A(p_input[8209]), .B(p_input[38209]), .Z(n3981) );
  AND U5974 ( .A(n3983), .B(n3984), .Z(o[8208]) );
  AND U5975 ( .A(p_input[28208]), .B(p_input[18208]), .Z(n3984) );
  AND U5976 ( .A(p_input[8208]), .B(p_input[38208]), .Z(n3983) );
  AND U5977 ( .A(n3985), .B(n3986), .Z(o[8207]) );
  AND U5978 ( .A(p_input[28207]), .B(p_input[18207]), .Z(n3986) );
  AND U5979 ( .A(p_input[8207]), .B(p_input[38207]), .Z(n3985) );
  AND U5980 ( .A(n3987), .B(n3988), .Z(o[8206]) );
  AND U5981 ( .A(p_input[28206]), .B(p_input[18206]), .Z(n3988) );
  AND U5982 ( .A(p_input[8206]), .B(p_input[38206]), .Z(n3987) );
  AND U5983 ( .A(n3989), .B(n3990), .Z(o[8205]) );
  AND U5984 ( .A(p_input[28205]), .B(p_input[18205]), .Z(n3990) );
  AND U5985 ( .A(p_input[8205]), .B(p_input[38205]), .Z(n3989) );
  AND U5986 ( .A(n3991), .B(n3992), .Z(o[8204]) );
  AND U5987 ( .A(p_input[28204]), .B(p_input[18204]), .Z(n3992) );
  AND U5988 ( .A(p_input[8204]), .B(p_input[38204]), .Z(n3991) );
  AND U5989 ( .A(n3993), .B(n3994), .Z(o[8203]) );
  AND U5990 ( .A(p_input[28203]), .B(p_input[18203]), .Z(n3994) );
  AND U5991 ( .A(p_input[8203]), .B(p_input[38203]), .Z(n3993) );
  AND U5992 ( .A(n3995), .B(n3996), .Z(o[8202]) );
  AND U5993 ( .A(p_input[28202]), .B(p_input[18202]), .Z(n3996) );
  AND U5994 ( .A(p_input[8202]), .B(p_input[38202]), .Z(n3995) );
  AND U5995 ( .A(n3997), .B(n3998), .Z(o[8201]) );
  AND U5996 ( .A(p_input[28201]), .B(p_input[18201]), .Z(n3998) );
  AND U5997 ( .A(p_input[8201]), .B(p_input[38201]), .Z(n3997) );
  AND U5998 ( .A(n3999), .B(n4000), .Z(o[8200]) );
  AND U5999 ( .A(p_input[28200]), .B(p_input[18200]), .Z(n4000) );
  AND U6000 ( .A(p_input[8200]), .B(p_input[38200]), .Z(n3999) );
  AND U6001 ( .A(n4001), .B(n4002), .Z(o[81]) );
  AND U6002 ( .A(p_input[20081]), .B(p_input[10081]), .Z(n4002) );
  AND U6003 ( .A(p_input[81]), .B(p_input[30081]), .Z(n4001) );
  AND U6004 ( .A(n4003), .B(n4004), .Z(o[819]) );
  AND U6005 ( .A(p_input[20819]), .B(p_input[10819]), .Z(n4004) );
  AND U6006 ( .A(p_input[819]), .B(p_input[30819]), .Z(n4003) );
  AND U6007 ( .A(n4005), .B(n4006), .Z(o[8199]) );
  AND U6008 ( .A(p_input[28199]), .B(p_input[18199]), .Z(n4006) );
  AND U6009 ( .A(p_input[8199]), .B(p_input[38199]), .Z(n4005) );
  AND U6010 ( .A(n4007), .B(n4008), .Z(o[8198]) );
  AND U6011 ( .A(p_input[28198]), .B(p_input[18198]), .Z(n4008) );
  AND U6012 ( .A(p_input[8198]), .B(p_input[38198]), .Z(n4007) );
  AND U6013 ( .A(n4009), .B(n4010), .Z(o[8197]) );
  AND U6014 ( .A(p_input[28197]), .B(p_input[18197]), .Z(n4010) );
  AND U6015 ( .A(p_input[8197]), .B(p_input[38197]), .Z(n4009) );
  AND U6016 ( .A(n4011), .B(n4012), .Z(o[8196]) );
  AND U6017 ( .A(p_input[28196]), .B(p_input[18196]), .Z(n4012) );
  AND U6018 ( .A(p_input[8196]), .B(p_input[38196]), .Z(n4011) );
  AND U6019 ( .A(n4013), .B(n4014), .Z(o[8195]) );
  AND U6020 ( .A(p_input[28195]), .B(p_input[18195]), .Z(n4014) );
  AND U6021 ( .A(p_input[8195]), .B(p_input[38195]), .Z(n4013) );
  AND U6022 ( .A(n4015), .B(n4016), .Z(o[8194]) );
  AND U6023 ( .A(p_input[28194]), .B(p_input[18194]), .Z(n4016) );
  AND U6024 ( .A(p_input[8194]), .B(p_input[38194]), .Z(n4015) );
  AND U6025 ( .A(n4017), .B(n4018), .Z(o[8193]) );
  AND U6026 ( .A(p_input[28193]), .B(p_input[18193]), .Z(n4018) );
  AND U6027 ( .A(p_input[8193]), .B(p_input[38193]), .Z(n4017) );
  AND U6028 ( .A(n4019), .B(n4020), .Z(o[8192]) );
  AND U6029 ( .A(p_input[28192]), .B(p_input[18192]), .Z(n4020) );
  AND U6030 ( .A(p_input[8192]), .B(p_input[38192]), .Z(n4019) );
  AND U6031 ( .A(n4021), .B(n4022), .Z(o[8191]) );
  AND U6032 ( .A(p_input[28191]), .B(p_input[18191]), .Z(n4022) );
  AND U6033 ( .A(p_input[8191]), .B(p_input[38191]), .Z(n4021) );
  AND U6034 ( .A(n4023), .B(n4024), .Z(o[8190]) );
  AND U6035 ( .A(p_input[28190]), .B(p_input[18190]), .Z(n4024) );
  AND U6036 ( .A(p_input[8190]), .B(p_input[38190]), .Z(n4023) );
  AND U6037 ( .A(n4025), .B(n4026), .Z(o[818]) );
  AND U6038 ( .A(p_input[20818]), .B(p_input[10818]), .Z(n4026) );
  AND U6039 ( .A(p_input[818]), .B(p_input[30818]), .Z(n4025) );
  AND U6040 ( .A(n4027), .B(n4028), .Z(o[8189]) );
  AND U6041 ( .A(p_input[28189]), .B(p_input[18189]), .Z(n4028) );
  AND U6042 ( .A(p_input[8189]), .B(p_input[38189]), .Z(n4027) );
  AND U6043 ( .A(n4029), .B(n4030), .Z(o[8188]) );
  AND U6044 ( .A(p_input[28188]), .B(p_input[18188]), .Z(n4030) );
  AND U6045 ( .A(p_input[8188]), .B(p_input[38188]), .Z(n4029) );
  AND U6046 ( .A(n4031), .B(n4032), .Z(o[8187]) );
  AND U6047 ( .A(p_input[28187]), .B(p_input[18187]), .Z(n4032) );
  AND U6048 ( .A(p_input[8187]), .B(p_input[38187]), .Z(n4031) );
  AND U6049 ( .A(n4033), .B(n4034), .Z(o[8186]) );
  AND U6050 ( .A(p_input[28186]), .B(p_input[18186]), .Z(n4034) );
  AND U6051 ( .A(p_input[8186]), .B(p_input[38186]), .Z(n4033) );
  AND U6052 ( .A(n4035), .B(n4036), .Z(o[8185]) );
  AND U6053 ( .A(p_input[28185]), .B(p_input[18185]), .Z(n4036) );
  AND U6054 ( .A(p_input[8185]), .B(p_input[38185]), .Z(n4035) );
  AND U6055 ( .A(n4037), .B(n4038), .Z(o[8184]) );
  AND U6056 ( .A(p_input[28184]), .B(p_input[18184]), .Z(n4038) );
  AND U6057 ( .A(p_input[8184]), .B(p_input[38184]), .Z(n4037) );
  AND U6058 ( .A(n4039), .B(n4040), .Z(o[8183]) );
  AND U6059 ( .A(p_input[28183]), .B(p_input[18183]), .Z(n4040) );
  AND U6060 ( .A(p_input[8183]), .B(p_input[38183]), .Z(n4039) );
  AND U6061 ( .A(n4041), .B(n4042), .Z(o[8182]) );
  AND U6062 ( .A(p_input[28182]), .B(p_input[18182]), .Z(n4042) );
  AND U6063 ( .A(p_input[8182]), .B(p_input[38182]), .Z(n4041) );
  AND U6064 ( .A(n4043), .B(n4044), .Z(o[8181]) );
  AND U6065 ( .A(p_input[28181]), .B(p_input[18181]), .Z(n4044) );
  AND U6066 ( .A(p_input[8181]), .B(p_input[38181]), .Z(n4043) );
  AND U6067 ( .A(n4045), .B(n4046), .Z(o[8180]) );
  AND U6068 ( .A(p_input[28180]), .B(p_input[18180]), .Z(n4046) );
  AND U6069 ( .A(p_input[8180]), .B(p_input[38180]), .Z(n4045) );
  AND U6070 ( .A(n4047), .B(n4048), .Z(o[817]) );
  AND U6071 ( .A(p_input[20817]), .B(p_input[10817]), .Z(n4048) );
  AND U6072 ( .A(p_input[817]), .B(p_input[30817]), .Z(n4047) );
  AND U6073 ( .A(n4049), .B(n4050), .Z(o[8179]) );
  AND U6074 ( .A(p_input[28179]), .B(p_input[18179]), .Z(n4050) );
  AND U6075 ( .A(p_input[8179]), .B(p_input[38179]), .Z(n4049) );
  AND U6076 ( .A(n4051), .B(n4052), .Z(o[8178]) );
  AND U6077 ( .A(p_input[28178]), .B(p_input[18178]), .Z(n4052) );
  AND U6078 ( .A(p_input[8178]), .B(p_input[38178]), .Z(n4051) );
  AND U6079 ( .A(n4053), .B(n4054), .Z(o[8177]) );
  AND U6080 ( .A(p_input[28177]), .B(p_input[18177]), .Z(n4054) );
  AND U6081 ( .A(p_input[8177]), .B(p_input[38177]), .Z(n4053) );
  AND U6082 ( .A(n4055), .B(n4056), .Z(o[8176]) );
  AND U6083 ( .A(p_input[28176]), .B(p_input[18176]), .Z(n4056) );
  AND U6084 ( .A(p_input[8176]), .B(p_input[38176]), .Z(n4055) );
  AND U6085 ( .A(n4057), .B(n4058), .Z(o[8175]) );
  AND U6086 ( .A(p_input[28175]), .B(p_input[18175]), .Z(n4058) );
  AND U6087 ( .A(p_input[8175]), .B(p_input[38175]), .Z(n4057) );
  AND U6088 ( .A(n4059), .B(n4060), .Z(o[8174]) );
  AND U6089 ( .A(p_input[28174]), .B(p_input[18174]), .Z(n4060) );
  AND U6090 ( .A(p_input[8174]), .B(p_input[38174]), .Z(n4059) );
  AND U6091 ( .A(n4061), .B(n4062), .Z(o[8173]) );
  AND U6092 ( .A(p_input[28173]), .B(p_input[18173]), .Z(n4062) );
  AND U6093 ( .A(p_input[8173]), .B(p_input[38173]), .Z(n4061) );
  AND U6094 ( .A(n4063), .B(n4064), .Z(o[8172]) );
  AND U6095 ( .A(p_input[28172]), .B(p_input[18172]), .Z(n4064) );
  AND U6096 ( .A(p_input[8172]), .B(p_input[38172]), .Z(n4063) );
  AND U6097 ( .A(n4065), .B(n4066), .Z(o[8171]) );
  AND U6098 ( .A(p_input[28171]), .B(p_input[18171]), .Z(n4066) );
  AND U6099 ( .A(p_input[8171]), .B(p_input[38171]), .Z(n4065) );
  AND U6100 ( .A(n4067), .B(n4068), .Z(o[8170]) );
  AND U6101 ( .A(p_input[28170]), .B(p_input[18170]), .Z(n4068) );
  AND U6102 ( .A(p_input[8170]), .B(p_input[38170]), .Z(n4067) );
  AND U6103 ( .A(n4069), .B(n4070), .Z(o[816]) );
  AND U6104 ( .A(p_input[20816]), .B(p_input[10816]), .Z(n4070) );
  AND U6105 ( .A(p_input[816]), .B(p_input[30816]), .Z(n4069) );
  AND U6106 ( .A(n4071), .B(n4072), .Z(o[8169]) );
  AND U6107 ( .A(p_input[28169]), .B(p_input[18169]), .Z(n4072) );
  AND U6108 ( .A(p_input[8169]), .B(p_input[38169]), .Z(n4071) );
  AND U6109 ( .A(n4073), .B(n4074), .Z(o[8168]) );
  AND U6110 ( .A(p_input[28168]), .B(p_input[18168]), .Z(n4074) );
  AND U6111 ( .A(p_input[8168]), .B(p_input[38168]), .Z(n4073) );
  AND U6112 ( .A(n4075), .B(n4076), .Z(o[8167]) );
  AND U6113 ( .A(p_input[28167]), .B(p_input[18167]), .Z(n4076) );
  AND U6114 ( .A(p_input[8167]), .B(p_input[38167]), .Z(n4075) );
  AND U6115 ( .A(n4077), .B(n4078), .Z(o[8166]) );
  AND U6116 ( .A(p_input[28166]), .B(p_input[18166]), .Z(n4078) );
  AND U6117 ( .A(p_input[8166]), .B(p_input[38166]), .Z(n4077) );
  AND U6118 ( .A(n4079), .B(n4080), .Z(o[8165]) );
  AND U6119 ( .A(p_input[28165]), .B(p_input[18165]), .Z(n4080) );
  AND U6120 ( .A(p_input[8165]), .B(p_input[38165]), .Z(n4079) );
  AND U6121 ( .A(n4081), .B(n4082), .Z(o[8164]) );
  AND U6122 ( .A(p_input[28164]), .B(p_input[18164]), .Z(n4082) );
  AND U6123 ( .A(p_input[8164]), .B(p_input[38164]), .Z(n4081) );
  AND U6124 ( .A(n4083), .B(n4084), .Z(o[8163]) );
  AND U6125 ( .A(p_input[28163]), .B(p_input[18163]), .Z(n4084) );
  AND U6126 ( .A(p_input[8163]), .B(p_input[38163]), .Z(n4083) );
  AND U6127 ( .A(n4085), .B(n4086), .Z(o[8162]) );
  AND U6128 ( .A(p_input[28162]), .B(p_input[18162]), .Z(n4086) );
  AND U6129 ( .A(p_input[8162]), .B(p_input[38162]), .Z(n4085) );
  AND U6130 ( .A(n4087), .B(n4088), .Z(o[8161]) );
  AND U6131 ( .A(p_input[28161]), .B(p_input[18161]), .Z(n4088) );
  AND U6132 ( .A(p_input[8161]), .B(p_input[38161]), .Z(n4087) );
  AND U6133 ( .A(n4089), .B(n4090), .Z(o[8160]) );
  AND U6134 ( .A(p_input[28160]), .B(p_input[18160]), .Z(n4090) );
  AND U6135 ( .A(p_input[8160]), .B(p_input[38160]), .Z(n4089) );
  AND U6136 ( .A(n4091), .B(n4092), .Z(o[815]) );
  AND U6137 ( .A(p_input[20815]), .B(p_input[10815]), .Z(n4092) );
  AND U6138 ( .A(p_input[815]), .B(p_input[30815]), .Z(n4091) );
  AND U6139 ( .A(n4093), .B(n4094), .Z(o[8159]) );
  AND U6140 ( .A(p_input[28159]), .B(p_input[18159]), .Z(n4094) );
  AND U6141 ( .A(p_input[8159]), .B(p_input[38159]), .Z(n4093) );
  AND U6142 ( .A(n4095), .B(n4096), .Z(o[8158]) );
  AND U6143 ( .A(p_input[28158]), .B(p_input[18158]), .Z(n4096) );
  AND U6144 ( .A(p_input[8158]), .B(p_input[38158]), .Z(n4095) );
  AND U6145 ( .A(n4097), .B(n4098), .Z(o[8157]) );
  AND U6146 ( .A(p_input[28157]), .B(p_input[18157]), .Z(n4098) );
  AND U6147 ( .A(p_input[8157]), .B(p_input[38157]), .Z(n4097) );
  AND U6148 ( .A(n4099), .B(n4100), .Z(o[8156]) );
  AND U6149 ( .A(p_input[28156]), .B(p_input[18156]), .Z(n4100) );
  AND U6150 ( .A(p_input[8156]), .B(p_input[38156]), .Z(n4099) );
  AND U6151 ( .A(n4101), .B(n4102), .Z(o[8155]) );
  AND U6152 ( .A(p_input[28155]), .B(p_input[18155]), .Z(n4102) );
  AND U6153 ( .A(p_input[8155]), .B(p_input[38155]), .Z(n4101) );
  AND U6154 ( .A(n4103), .B(n4104), .Z(o[8154]) );
  AND U6155 ( .A(p_input[28154]), .B(p_input[18154]), .Z(n4104) );
  AND U6156 ( .A(p_input[8154]), .B(p_input[38154]), .Z(n4103) );
  AND U6157 ( .A(n4105), .B(n4106), .Z(o[8153]) );
  AND U6158 ( .A(p_input[28153]), .B(p_input[18153]), .Z(n4106) );
  AND U6159 ( .A(p_input[8153]), .B(p_input[38153]), .Z(n4105) );
  AND U6160 ( .A(n4107), .B(n4108), .Z(o[8152]) );
  AND U6161 ( .A(p_input[28152]), .B(p_input[18152]), .Z(n4108) );
  AND U6162 ( .A(p_input[8152]), .B(p_input[38152]), .Z(n4107) );
  AND U6163 ( .A(n4109), .B(n4110), .Z(o[8151]) );
  AND U6164 ( .A(p_input[28151]), .B(p_input[18151]), .Z(n4110) );
  AND U6165 ( .A(p_input[8151]), .B(p_input[38151]), .Z(n4109) );
  AND U6166 ( .A(n4111), .B(n4112), .Z(o[8150]) );
  AND U6167 ( .A(p_input[28150]), .B(p_input[18150]), .Z(n4112) );
  AND U6168 ( .A(p_input[8150]), .B(p_input[38150]), .Z(n4111) );
  AND U6169 ( .A(n4113), .B(n4114), .Z(o[814]) );
  AND U6170 ( .A(p_input[20814]), .B(p_input[10814]), .Z(n4114) );
  AND U6171 ( .A(p_input[814]), .B(p_input[30814]), .Z(n4113) );
  AND U6172 ( .A(n4115), .B(n4116), .Z(o[8149]) );
  AND U6173 ( .A(p_input[28149]), .B(p_input[18149]), .Z(n4116) );
  AND U6174 ( .A(p_input[8149]), .B(p_input[38149]), .Z(n4115) );
  AND U6175 ( .A(n4117), .B(n4118), .Z(o[8148]) );
  AND U6176 ( .A(p_input[28148]), .B(p_input[18148]), .Z(n4118) );
  AND U6177 ( .A(p_input[8148]), .B(p_input[38148]), .Z(n4117) );
  AND U6178 ( .A(n4119), .B(n4120), .Z(o[8147]) );
  AND U6179 ( .A(p_input[28147]), .B(p_input[18147]), .Z(n4120) );
  AND U6180 ( .A(p_input[8147]), .B(p_input[38147]), .Z(n4119) );
  AND U6181 ( .A(n4121), .B(n4122), .Z(o[8146]) );
  AND U6182 ( .A(p_input[28146]), .B(p_input[18146]), .Z(n4122) );
  AND U6183 ( .A(p_input[8146]), .B(p_input[38146]), .Z(n4121) );
  AND U6184 ( .A(n4123), .B(n4124), .Z(o[8145]) );
  AND U6185 ( .A(p_input[28145]), .B(p_input[18145]), .Z(n4124) );
  AND U6186 ( .A(p_input[8145]), .B(p_input[38145]), .Z(n4123) );
  AND U6187 ( .A(n4125), .B(n4126), .Z(o[8144]) );
  AND U6188 ( .A(p_input[28144]), .B(p_input[18144]), .Z(n4126) );
  AND U6189 ( .A(p_input[8144]), .B(p_input[38144]), .Z(n4125) );
  AND U6190 ( .A(n4127), .B(n4128), .Z(o[8143]) );
  AND U6191 ( .A(p_input[28143]), .B(p_input[18143]), .Z(n4128) );
  AND U6192 ( .A(p_input[8143]), .B(p_input[38143]), .Z(n4127) );
  AND U6193 ( .A(n4129), .B(n4130), .Z(o[8142]) );
  AND U6194 ( .A(p_input[28142]), .B(p_input[18142]), .Z(n4130) );
  AND U6195 ( .A(p_input[8142]), .B(p_input[38142]), .Z(n4129) );
  AND U6196 ( .A(n4131), .B(n4132), .Z(o[8141]) );
  AND U6197 ( .A(p_input[28141]), .B(p_input[18141]), .Z(n4132) );
  AND U6198 ( .A(p_input[8141]), .B(p_input[38141]), .Z(n4131) );
  AND U6199 ( .A(n4133), .B(n4134), .Z(o[8140]) );
  AND U6200 ( .A(p_input[28140]), .B(p_input[18140]), .Z(n4134) );
  AND U6201 ( .A(p_input[8140]), .B(p_input[38140]), .Z(n4133) );
  AND U6202 ( .A(n4135), .B(n4136), .Z(o[813]) );
  AND U6203 ( .A(p_input[20813]), .B(p_input[10813]), .Z(n4136) );
  AND U6204 ( .A(p_input[813]), .B(p_input[30813]), .Z(n4135) );
  AND U6205 ( .A(n4137), .B(n4138), .Z(o[8139]) );
  AND U6206 ( .A(p_input[28139]), .B(p_input[18139]), .Z(n4138) );
  AND U6207 ( .A(p_input[8139]), .B(p_input[38139]), .Z(n4137) );
  AND U6208 ( .A(n4139), .B(n4140), .Z(o[8138]) );
  AND U6209 ( .A(p_input[28138]), .B(p_input[18138]), .Z(n4140) );
  AND U6210 ( .A(p_input[8138]), .B(p_input[38138]), .Z(n4139) );
  AND U6211 ( .A(n4141), .B(n4142), .Z(o[8137]) );
  AND U6212 ( .A(p_input[28137]), .B(p_input[18137]), .Z(n4142) );
  AND U6213 ( .A(p_input[8137]), .B(p_input[38137]), .Z(n4141) );
  AND U6214 ( .A(n4143), .B(n4144), .Z(o[8136]) );
  AND U6215 ( .A(p_input[28136]), .B(p_input[18136]), .Z(n4144) );
  AND U6216 ( .A(p_input[8136]), .B(p_input[38136]), .Z(n4143) );
  AND U6217 ( .A(n4145), .B(n4146), .Z(o[8135]) );
  AND U6218 ( .A(p_input[28135]), .B(p_input[18135]), .Z(n4146) );
  AND U6219 ( .A(p_input[8135]), .B(p_input[38135]), .Z(n4145) );
  AND U6220 ( .A(n4147), .B(n4148), .Z(o[8134]) );
  AND U6221 ( .A(p_input[28134]), .B(p_input[18134]), .Z(n4148) );
  AND U6222 ( .A(p_input[8134]), .B(p_input[38134]), .Z(n4147) );
  AND U6223 ( .A(n4149), .B(n4150), .Z(o[8133]) );
  AND U6224 ( .A(p_input[28133]), .B(p_input[18133]), .Z(n4150) );
  AND U6225 ( .A(p_input[8133]), .B(p_input[38133]), .Z(n4149) );
  AND U6226 ( .A(n4151), .B(n4152), .Z(o[8132]) );
  AND U6227 ( .A(p_input[28132]), .B(p_input[18132]), .Z(n4152) );
  AND U6228 ( .A(p_input[8132]), .B(p_input[38132]), .Z(n4151) );
  AND U6229 ( .A(n4153), .B(n4154), .Z(o[8131]) );
  AND U6230 ( .A(p_input[28131]), .B(p_input[18131]), .Z(n4154) );
  AND U6231 ( .A(p_input[8131]), .B(p_input[38131]), .Z(n4153) );
  AND U6232 ( .A(n4155), .B(n4156), .Z(o[8130]) );
  AND U6233 ( .A(p_input[28130]), .B(p_input[18130]), .Z(n4156) );
  AND U6234 ( .A(p_input[8130]), .B(p_input[38130]), .Z(n4155) );
  AND U6235 ( .A(n4157), .B(n4158), .Z(o[812]) );
  AND U6236 ( .A(p_input[20812]), .B(p_input[10812]), .Z(n4158) );
  AND U6237 ( .A(p_input[812]), .B(p_input[30812]), .Z(n4157) );
  AND U6238 ( .A(n4159), .B(n4160), .Z(o[8129]) );
  AND U6239 ( .A(p_input[28129]), .B(p_input[18129]), .Z(n4160) );
  AND U6240 ( .A(p_input[8129]), .B(p_input[38129]), .Z(n4159) );
  AND U6241 ( .A(n4161), .B(n4162), .Z(o[8128]) );
  AND U6242 ( .A(p_input[28128]), .B(p_input[18128]), .Z(n4162) );
  AND U6243 ( .A(p_input[8128]), .B(p_input[38128]), .Z(n4161) );
  AND U6244 ( .A(n4163), .B(n4164), .Z(o[8127]) );
  AND U6245 ( .A(p_input[28127]), .B(p_input[18127]), .Z(n4164) );
  AND U6246 ( .A(p_input[8127]), .B(p_input[38127]), .Z(n4163) );
  AND U6247 ( .A(n4165), .B(n4166), .Z(o[8126]) );
  AND U6248 ( .A(p_input[28126]), .B(p_input[18126]), .Z(n4166) );
  AND U6249 ( .A(p_input[8126]), .B(p_input[38126]), .Z(n4165) );
  AND U6250 ( .A(n4167), .B(n4168), .Z(o[8125]) );
  AND U6251 ( .A(p_input[28125]), .B(p_input[18125]), .Z(n4168) );
  AND U6252 ( .A(p_input[8125]), .B(p_input[38125]), .Z(n4167) );
  AND U6253 ( .A(n4169), .B(n4170), .Z(o[8124]) );
  AND U6254 ( .A(p_input[28124]), .B(p_input[18124]), .Z(n4170) );
  AND U6255 ( .A(p_input[8124]), .B(p_input[38124]), .Z(n4169) );
  AND U6256 ( .A(n4171), .B(n4172), .Z(o[8123]) );
  AND U6257 ( .A(p_input[28123]), .B(p_input[18123]), .Z(n4172) );
  AND U6258 ( .A(p_input[8123]), .B(p_input[38123]), .Z(n4171) );
  AND U6259 ( .A(n4173), .B(n4174), .Z(o[8122]) );
  AND U6260 ( .A(p_input[28122]), .B(p_input[18122]), .Z(n4174) );
  AND U6261 ( .A(p_input[8122]), .B(p_input[38122]), .Z(n4173) );
  AND U6262 ( .A(n4175), .B(n4176), .Z(o[8121]) );
  AND U6263 ( .A(p_input[28121]), .B(p_input[18121]), .Z(n4176) );
  AND U6264 ( .A(p_input[8121]), .B(p_input[38121]), .Z(n4175) );
  AND U6265 ( .A(n4177), .B(n4178), .Z(o[8120]) );
  AND U6266 ( .A(p_input[28120]), .B(p_input[18120]), .Z(n4178) );
  AND U6267 ( .A(p_input[8120]), .B(p_input[38120]), .Z(n4177) );
  AND U6268 ( .A(n4179), .B(n4180), .Z(o[811]) );
  AND U6269 ( .A(p_input[20811]), .B(p_input[10811]), .Z(n4180) );
  AND U6270 ( .A(p_input[811]), .B(p_input[30811]), .Z(n4179) );
  AND U6271 ( .A(n4181), .B(n4182), .Z(o[8119]) );
  AND U6272 ( .A(p_input[28119]), .B(p_input[18119]), .Z(n4182) );
  AND U6273 ( .A(p_input[8119]), .B(p_input[38119]), .Z(n4181) );
  AND U6274 ( .A(n4183), .B(n4184), .Z(o[8118]) );
  AND U6275 ( .A(p_input[28118]), .B(p_input[18118]), .Z(n4184) );
  AND U6276 ( .A(p_input[8118]), .B(p_input[38118]), .Z(n4183) );
  AND U6277 ( .A(n4185), .B(n4186), .Z(o[8117]) );
  AND U6278 ( .A(p_input[28117]), .B(p_input[18117]), .Z(n4186) );
  AND U6279 ( .A(p_input[8117]), .B(p_input[38117]), .Z(n4185) );
  AND U6280 ( .A(n4187), .B(n4188), .Z(o[8116]) );
  AND U6281 ( .A(p_input[28116]), .B(p_input[18116]), .Z(n4188) );
  AND U6282 ( .A(p_input[8116]), .B(p_input[38116]), .Z(n4187) );
  AND U6283 ( .A(n4189), .B(n4190), .Z(o[8115]) );
  AND U6284 ( .A(p_input[28115]), .B(p_input[18115]), .Z(n4190) );
  AND U6285 ( .A(p_input[8115]), .B(p_input[38115]), .Z(n4189) );
  AND U6286 ( .A(n4191), .B(n4192), .Z(o[8114]) );
  AND U6287 ( .A(p_input[28114]), .B(p_input[18114]), .Z(n4192) );
  AND U6288 ( .A(p_input[8114]), .B(p_input[38114]), .Z(n4191) );
  AND U6289 ( .A(n4193), .B(n4194), .Z(o[8113]) );
  AND U6290 ( .A(p_input[28113]), .B(p_input[18113]), .Z(n4194) );
  AND U6291 ( .A(p_input[8113]), .B(p_input[38113]), .Z(n4193) );
  AND U6292 ( .A(n4195), .B(n4196), .Z(o[8112]) );
  AND U6293 ( .A(p_input[28112]), .B(p_input[18112]), .Z(n4196) );
  AND U6294 ( .A(p_input[8112]), .B(p_input[38112]), .Z(n4195) );
  AND U6295 ( .A(n4197), .B(n4198), .Z(o[8111]) );
  AND U6296 ( .A(p_input[28111]), .B(p_input[18111]), .Z(n4198) );
  AND U6297 ( .A(p_input[8111]), .B(p_input[38111]), .Z(n4197) );
  AND U6298 ( .A(n4199), .B(n4200), .Z(o[8110]) );
  AND U6299 ( .A(p_input[28110]), .B(p_input[18110]), .Z(n4200) );
  AND U6300 ( .A(p_input[8110]), .B(p_input[38110]), .Z(n4199) );
  AND U6301 ( .A(n4201), .B(n4202), .Z(o[810]) );
  AND U6302 ( .A(p_input[20810]), .B(p_input[10810]), .Z(n4202) );
  AND U6303 ( .A(p_input[810]), .B(p_input[30810]), .Z(n4201) );
  AND U6304 ( .A(n4203), .B(n4204), .Z(o[8109]) );
  AND U6305 ( .A(p_input[28109]), .B(p_input[18109]), .Z(n4204) );
  AND U6306 ( .A(p_input[8109]), .B(p_input[38109]), .Z(n4203) );
  AND U6307 ( .A(n4205), .B(n4206), .Z(o[8108]) );
  AND U6308 ( .A(p_input[28108]), .B(p_input[18108]), .Z(n4206) );
  AND U6309 ( .A(p_input[8108]), .B(p_input[38108]), .Z(n4205) );
  AND U6310 ( .A(n4207), .B(n4208), .Z(o[8107]) );
  AND U6311 ( .A(p_input[28107]), .B(p_input[18107]), .Z(n4208) );
  AND U6312 ( .A(p_input[8107]), .B(p_input[38107]), .Z(n4207) );
  AND U6313 ( .A(n4209), .B(n4210), .Z(o[8106]) );
  AND U6314 ( .A(p_input[28106]), .B(p_input[18106]), .Z(n4210) );
  AND U6315 ( .A(p_input[8106]), .B(p_input[38106]), .Z(n4209) );
  AND U6316 ( .A(n4211), .B(n4212), .Z(o[8105]) );
  AND U6317 ( .A(p_input[28105]), .B(p_input[18105]), .Z(n4212) );
  AND U6318 ( .A(p_input[8105]), .B(p_input[38105]), .Z(n4211) );
  AND U6319 ( .A(n4213), .B(n4214), .Z(o[8104]) );
  AND U6320 ( .A(p_input[28104]), .B(p_input[18104]), .Z(n4214) );
  AND U6321 ( .A(p_input[8104]), .B(p_input[38104]), .Z(n4213) );
  AND U6322 ( .A(n4215), .B(n4216), .Z(o[8103]) );
  AND U6323 ( .A(p_input[28103]), .B(p_input[18103]), .Z(n4216) );
  AND U6324 ( .A(p_input[8103]), .B(p_input[38103]), .Z(n4215) );
  AND U6325 ( .A(n4217), .B(n4218), .Z(o[8102]) );
  AND U6326 ( .A(p_input[28102]), .B(p_input[18102]), .Z(n4218) );
  AND U6327 ( .A(p_input[8102]), .B(p_input[38102]), .Z(n4217) );
  AND U6328 ( .A(n4219), .B(n4220), .Z(o[8101]) );
  AND U6329 ( .A(p_input[28101]), .B(p_input[18101]), .Z(n4220) );
  AND U6330 ( .A(p_input[8101]), .B(p_input[38101]), .Z(n4219) );
  AND U6331 ( .A(n4221), .B(n4222), .Z(o[8100]) );
  AND U6332 ( .A(p_input[28100]), .B(p_input[18100]), .Z(n4222) );
  AND U6333 ( .A(p_input[8100]), .B(p_input[38100]), .Z(n4221) );
  AND U6334 ( .A(n4223), .B(n4224), .Z(o[80]) );
  AND U6335 ( .A(p_input[20080]), .B(p_input[10080]), .Z(n4224) );
  AND U6336 ( .A(p_input[80]), .B(p_input[30080]), .Z(n4223) );
  AND U6337 ( .A(n4225), .B(n4226), .Z(o[809]) );
  AND U6338 ( .A(p_input[20809]), .B(p_input[10809]), .Z(n4226) );
  AND U6339 ( .A(p_input[809]), .B(p_input[30809]), .Z(n4225) );
  AND U6340 ( .A(n4227), .B(n4228), .Z(o[8099]) );
  AND U6341 ( .A(p_input[28099]), .B(p_input[18099]), .Z(n4228) );
  AND U6342 ( .A(p_input[8099]), .B(p_input[38099]), .Z(n4227) );
  AND U6343 ( .A(n4229), .B(n4230), .Z(o[8098]) );
  AND U6344 ( .A(p_input[28098]), .B(p_input[18098]), .Z(n4230) );
  AND U6345 ( .A(p_input[8098]), .B(p_input[38098]), .Z(n4229) );
  AND U6346 ( .A(n4231), .B(n4232), .Z(o[8097]) );
  AND U6347 ( .A(p_input[28097]), .B(p_input[18097]), .Z(n4232) );
  AND U6348 ( .A(p_input[8097]), .B(p_input[38097]), .Z(n4231) );
  AND U6349 ( .A(n4233), .B(n4234), .Z(o[8096]) );
  AND U6350 ( .A(p_input[28096]), .B(p_input[18096]), .Z(n4234) );
  AND U6351 ( .A(p_input[8096]), .B(p_input[38096]), .Z(n4233) );
  AND U6352 ( .A(n4235), .B(n4236), .Z(o[8095]) );
  AND U6353 ( .A(p_input[28095]), .B(p_input[18095]), .Z(n4236) );
  AND U6354 ( .A(p_input[8095]), .B(p_input[38095]), .Z(n4235) );
  AND U6355 ( .A(n4237), .B(n4238), .Z(o[8094]) );
  AND U6356 ( .A(p_input[28094]), .B(p_input[18094]), .Z(n4238) );
  AND U6357 ( .A(p_input[8094]), .B(p_input[38094]), .Z(n4237) );
  AND U6358 ( .A(n4239), .B(n4240), .Z(o[8093]) );
  AND U6359 ( .A(p_input[28093]), .B(p_input[18093]), .Z(n4240) );
  AND U6360 ( .A(p_input[8093]), .B(p_input[38093]), .Z(n4239) );
  AND U6361 ( .A(n4241), .B(n4242), .Z(o[8092]) );
  AND U6362 ( .A(p_input[28092]), .B(p_input[18092]), .Z(n4242) );
  AND U6363 ( .A(p_input[8092]), .B(p_input[38092]), .Z(n4241) );
  AND U6364 ( .A(n4243), .B(n4244), .Z(o[8091]) );
  AND U6365 ( .A(p_input[28091]), .B(p_input[18091]), .Z(n4244) );
  AND U6366 ( .A(p_input[8091]), .B(p_input[38091]), .Z(n4243) );
  AND U6367 ( .A(n4245), .B(n4246), .Z(o[8090]) );
  AND U6368 ( .A(p_input[28090]), .B(p_input[18090]), .Z(n4246) );
  AND U6369 ( .A(p_input[8090]), .B(p_input[38090]), .Z(n4245) );
  AND U6370 ( .A(n4247), .B(n4248), .Z(o[808]) );
  AND U6371 ( .A(p_input[20808]), .B(p_input[10808]), .Z(n4248) );
  AND U6372 ( .A(p_input[808]), .B(p_input[30808]), .Z(n4247) );
  AND U6373 ( .A(n4249), .B(n4250), .Z(o[8089]) );
  AND U6374 ( .A(p_input[28089]), .B(p_input[18089]), .Z(n4250) );
  AND U6375 ( .A(p_input[8089]), .B(p_input[38089]), .Z(n4249) );
  AND U6376 ( .A(n4251), .B(n4252), .Z(o[8088]) );
  AND U6377 ( .A(p_input[28088]), .B(p_input[18088]), .Z(n4252) );
  AND U6378 ( .A(p_input[8088]), .B(p_input[38088]), .Z(n4251) );
  AND U6379 ( .A(n4253), .B(n4254), .Z(o[8087]) );
  AND U6380 ( .A(p_input[28087]), .B(p_input[18087]), .Z(n4254) );
  AND U6381 ( .A(p_input[8087]), .B(p_input[38087]), .Z(n4253) );
  AND U6382 ( .A(n4255), .B(n4256), .Z(o[8086]) );
  AND U6383 ( .A(p_input[28086]), .B(p_input[18086]), .Z(n4256) );
  AND U6384 ( .A(p_input[8086]), .B(p_input[38086]), .Z(n4255) );
  AND U6385 ( .A(n4257), .B(n4258), .Z(o[8085]) );
  AND U6386 ( .A(p_input[28085]), .B(p_input[18085]), .Z(n4258) );
  AND U6387 ( .A(p_input[8085]), .B(p_input[38085]), .Z(n4257) );
  AND U6388 ( .A(n4259), .B(n4260), .Z(o[8084]) );
  AND U6389 ( .A(p_input[28084]), .B(p_input[18084]), .Z(n4260) );
  AND U6390 ( .A(p_input[8084]), .B(p_input[38084]), .Z(n4259) );
  AND U6391 ( .A(n4261), .B(n4262), .Z(o[8083]) );
  AND U6392 ( .A(p_input[28083]), .B(p_input[18083]), .Z(n4262) );
  AND U6393 ( .A(p_input[8083]), .B(p_input[38083]), .Z(n4261) );
  AND U6394 ( .A(n4263), .B(n4264), .Z(o[8082]) );
  AND U6395 ( .A(p_input[28082]), .B(p_input[18082]), .Z(n4264) );
  AND U6396 ( .A(p_input[8082]), .B(p_input[38082]), .Z(n4263) );
  AND U6397 ( .A(n4265), .B(n4266), .Z(o[8081]) );
  AND U6398 ( .A(p_input[28081]), .B(p_input[18081]), .Z(n4266) );
  AND U6399 ( .A(p_input[8081]), .B(p_input[38081]), .Z(n4265) );
  AND U6400 ( .A(n4267), .B(n4268), .Z(o[8080]) );
  AND U6401 ( .A(p_input[28080]), .B(p_input[18080]), .Z(n4268) );
  AND U6402 ( .A(p_input[8080]), .B(p_input[38080]), .Z(n4267) );
  AND U6403 ( .A(n4269), .B(n4270), .Z(o[807]) );
  AND U6404 ( .A(p_input[20807]), .B(p_input[10807]), .Z(n4270) );
  AND U6405 ( .A(p_input[807]), .B(p_input[30807]), .Z(n4269) );
  AND U6406 ( .A(n4271), .B(n4272), .Z(o[8079]) );
  AND U6407 ( .A(p_input[28079]), .B(p_input[18079]), .Z(n4272) );
  AND U6408 ( .A(p_input[8079]), .B(p_input[38079]), .Z(n4271) );
  AND U6409 ( .A(n4273), .B(n4274), .Z(o[8078]) );
  AND U6410 ( .A(p_input[28078]), .B(p_input[18078]), .Z(n4274) );
  AND U6411 ( .A(p_input[8078]), .B(p_input[38078]), .Z(n4273) );
  AND U6412 ( .A(n4275), .B(n4276), .Z(o[8077]) );
  AND U6413 ( .A(p_input[28077]), .B(p_input[18077]), .Z(n4276) );
  AND U6414 ( .A(p_input[8077]), .B(p_input[38077]), .Z(n4275) );
  AND U6415 ( .A(n4277), .B(n4278), .Z(o[8076]) );
  AND U6416 ( .A(p_input[28076]), .B(p_input[18076]), .Z(n4278) );
  AND U6417 ( .A(p_input[8076]), .B(p_input[38076]), .Z(n4277) );
  AND U6418 ( .A(n4279), .B(n4280), .Z(o[8075]) );
  AND U6419 ( .A(p_input[28075]), .B(p_input[18075]), .Z(n4280) );
  AND U6420 ( .A(p_input[8075]), .B(p_input[38075]), .Z(n4279) );
  AND U6421 ( .A(n4281), .B(n4282), .Z(o[8074]) );
  AND U6422 ( .A(p_input[28074]), .B(p_input[18074]), .Z(n4282) );
  AND U6423 ( .A(p_input[8074]), .B(p_input[38074]), .Z(n4281) );
  AND U6424 ( .A(n4283), .B(n4284), .Z(o[8073]) );
  AND U6425 ( .A(p_input[28073]), .B(p_input[18073]), .Z(n4284) );
  AND U6426 ( .A(p_input[8073]), .B(p_input[38073]), .Z(n4283) );
  AND U6427 ( .A(n4285), .B(n4286), .Z(o[8072]) );
  AND U6428 ( .A(p_input[28072]), .B(p_input[18072]), .Z(n4286) );
  AND U6429 ( .A(p_input[8072]), .B(p_input[38072]), .Z(n4285) );
  AND U6430 ( .A(n4287), .B(n4288), .Z(o[8071]) );
  AND U6431 ( .A(p_input[28071]), .B(p_input[18071]), .Z(n4288) );
  AND U6432 ( .A(p_input[8071]), .B(p_input[38071]), .Z(n4287) );
  AND U6433 ( .A(n4289), .B(n4290), .Z(o[8070]) );
  AND U6434 ( .A(p_input[28070]), .B(p_input[18070]), .Z(n4290) );
  AND U6435 ( .A(p_input[8070]), .B(p_input[38070]), .Z(n4289) );
  AND U6436 ( .A(n4291), .B(n4292), .Z(o[806]) );
  AND U6437 ( .A(p_input[20806]), .B(p_input[10806]), .Z(n4292) );
  AND U6438 ( .A(p_input[806]), .B(p_input[30806]), .Z(n4291) );
  AND U6439 ( .A(n4293), .B(n4294), .Z(o[8069]) );
  AND U6440 ( .A(p_input[28069]), .B(p_input[18069]), .Z(n4294) );
  AND U6441 ( .A(p_input[8069]), .B(p_input[38069]), .Z(n4293) );
  AND U6442 ( .A(n4295), .B(n4296), .Z(o[8068]) );
  AND U6443 ( .A(p_input[28068]), .B(p_input[18068]), .Z(n4296) );
  AND U6444 ( .A(p_input[8068]), .B(p_input[38068]), .Z(n4295) );
  AND U6445 ( .A(n4297), .B(n4298), .Z(o[8067]) );
  AND U6446 ( .A(p_input[28067]), .B(p_input[18067]), .Z(n4298) );
  AND U6447 ( .A(p_input[8067]), .B(p_input[38067]), .Z(n4297) );
  AND U6448 ( .A(n4299), .B(n4300), .Z(o[8066]) );
  AND U6449 ( .A(p_input[28066]), .B(p_input[18066]), .Z(n4300) );
  AND U6450 ( .A(p_input[8066]), .B(p_input[38066]), .Z(n4299) );
  AND U6451 ( .A(n4301), .B(n4302), .Z(o[8065]) );
  AND U6452 ( .A(p_input[28065]), .B(p_input[18065]), .Z(n4302) );
  AND U6453 ( .A(p_input[8065]), .B(p_input[38065]), .Z(n4301) );
  AND U6454 ( .A(n4303), .B(n4304), .Z(o[8064]) );
  AND U6455 ( .A(p_input[28064]), .B(p_input[18064]), .Z(n4304) );
  AND U6456 ( .A(p_input[8064]), .B(p_input[38064]), .Z(n4303) );
  AND U6457 ( .A(n4305), .B(n4306), .Z(o[8063]) );
  AND U6458 ( .A(p_input[28063]), .B(p_input[18063]), .Z(n4306) );
  AND U6459 ( .A(p_input[8063]), .B(p_input[38063]), .Z(n4305) );
  AND U6460 ( .A(n4307), .B(n4308), .Z(o[8062]) );
  AND U6461 ( .A(p_input[28062]), .B(p_input[18062]), .Z(n4308) );
  AND U6462 ( .A(p_input[8062]), .B(p_input[38062]), .Z(n4307) );
  AND U6463 ( .A(n4309), .B(n4310), .Z(o[8061]) );
  AND U6464 ( .A(p_input[28061]), .B(p_input[18061]), .Z(n4310) );
  AND U6465 ( .A(p_input[8061]), .B(p_input[38061]), .Z(n4309) );
  AND U6466 ( .A(n4311), .B(n4312), .Z(o[8060]) );
  AND U6467 ( .A(p_input[28060]), .B(p_input[18060]), .Z(n4312) );
  AND U6468 ( .A(p_input[8060]), .B(p_input[38060]), .Z(n4311) );
  AND U6469 ( .A(n4313), .B(n4314), .Z(o[805]) );
  AND U6470 ( .A(p_input[20805]), .B(p_input[10805]), .Z(n4314) );
  AND U6471 ( .A(p_input[805]), .B(p_input[30805]), .Z(n4313) );
  AND U6472 ( .A(n4315), .B(n4316), .Z(o[8059]) );
  AND U6473 ( .A(p_input[28059]), .B(p_input[18059]), .Z(n4316) );
  AND U6474 ( .A(p_input[8059]), .B(p_input[38059]), .Z(n4315) );
  AND U6475 ( .A(n4317), .B(n4318), .Z(o[8058]) );
  AND U6476 ( .A(p_input[28058]), .B(p_input[18058]), .Z(n4318) );
  AND U6477 ( .A(p_input[8058]), .B(p_input[38058]), .Z(n4317) );
  AND U6478 ( .A(n4319), .B(n4320), .Z(o[8057]) );
  AND U6479 ( .A(p_input[28057]), .B(p_input[18057]), .Z(n4320) );
  AND U6480 ( .A(p_input[8057]), .B(p_input[38057]), .Z(n4319) );
  AND U6481 ( .A(n4321), .B(n4322), .Z(o[8056]) );
  AND U6482 ( .A(p_input[28056]), .B(p_input[18056]), .Z(n4322) );
  AND U6483 ( .A(p_input[8056]), .B(p_input[38056]), .Z(n4321) );
  AND U6484 ( .A(n4323), .B(n4324), .Z(o[8055]) );
  AND U6485 ( .A(p_input[28055]), .B(p_input[18055]), .Z(n4324) );
  AND U6486 ( .A(p_input[8055]), .B(p_input[38055]), .Z(n4323) );
  AND U6487 ( .A(n4325), .B(n4326), .Z(o[8054]) );
  AND U6488 ( .A(p_input[28054]), .B(p_input[18054]), .Z(n4326) );
  AND U6489 ( .A(p_input[8054]), .B(p_input[38054]), .Z(n4325) );
  AND U6490 ( .A(n4327), .B(n4328), .Z(o[8053]) );
  AND U6491 ( .A(p_input[28053]), .B(p_input[18053]), .Z(n4328) );
  AND U6492 ( .A(p_input[8053]), .B(p_input[38053]), .Z(n4327) );
  AND U6493 ( .A(n4329), .B(n4330), .Z(o[8052]) );
  AND U6494 ( .A(p_input[28052]), .B(p_input[18052]), .Z(n4330) );
  AND U6495 ( .A(p_input[8052]), .B(p_input[38052]), .Z(n4329) );
  AND U6496 ( .A(n4331), .B(n4332), .Z(o[8051]) );
  AND U6497 ( .A(p_input[28051]), .B(p_input[18051]), .Z(n4332) );
  AND U6498 ( .A(p_input[8051]), .B(p_input[38051]), .Z(n4331) );
  AND U6499 ( .A(n4333), .B(n4334), .Z(o[8050]) );
  AND U6500 ( .A(p_input[28050]), .B(p_input[18050]), .Z(n4334) );
  AND U6501 ( .A(p_input[8050]), .B(p_input[38050]), .Z(n4333) );
  AND U6502 ( .A(n4335), .B(n4336), .Z(o[804]) );
  AND U6503 ( .A(p_input[20804]), .B(p_input[10804]), .Z(n4336) );
  AND U6504 ( .A(p_input[804]), .B(p_input[30804]), .Z(n4335) );
  AND U6505 ( .A(n4337), .B(n4338), .Z(o[8049]) );
  AND U6506 ( .A(p_input[28049]), .B(p_input[18049]), .Z(n4338) );
  AND U6507 ( .A(p_input[8049]), .B(p_input[38049]), .Z(n4337) );
  AND U6508 ( .A(n4339), .B(n4340), .Z(o[8048]) );
  AND U6509 ( .A(p_input[28048]), .B(p_input[18048]), .Z(n4340) );
  AND U6510 ( .A(p_input[8048]), .B(p_input[38048]), .Z(n4339) );
  AND U6511 ( .A(n4341), .B(n4342), .Z(o[8047]) );
  AND U6512 ( .A(p_input[28047]), .B(p_input[18047]), .Z(n4342) );
  AND U6513 ( .A(p_input[8047]), .B(p_input[38047]), .Z(n4341) );
  AND U6514 ( .A(n4343), .B(n4344), .Z(o[8046]) );
  AND U6515 ( .A(p_input[28046]), .B(p_input[18046]), .Z(n4344) );
  AND U6516 ( .A(p_input[8046]), .B(p_input[38046]), .Z(n4343) );
  AND U6517 ( .A(n4345), .B(n4346), .Z(o[8045]) );
  AND U6518 ( .A(p_input[28045]), .B(p_input[18045]), .Z(n4346) );
  AND U6519 ( .A(p_input[8045]), .B(p_input[38045]), .Z(n4345) );
  AND U6520 ( .A(n4347), .B(n4348), .Z(o[8044]) );
  AND U6521 ( .A(p_input[28044]), .B(p_input[18044]), .Z(n4348) );
  AND U6522 ( .A(p_input[8044]), .B(p_input[38044]), .Z(n4347) );
  AND U6523 ( .A(n4349), .B(n4350), .Z(o[8043]) );
  AND U6524 ( .A(p_input[28043]), .B(p_input[18043]), .Z(n4350) );
  AND U6525 ( .A(p_input[8043]), .B(p_input[38043]), .Z(n4349) );
  AND U6526 ( .A(n4351), .B(n4352), .Z(o[8042]) );
  AND U6527 ( .A(p_input[28042]), .B(p_input[18042]), .Z(n4352) );
  AND U6528 ( .A(p_input[8042]), .B(p_input[38042]), .Z(n4351) );
  AND U6529 ( .A(n4353), .B(n4354), .Z(o[8041]) );
  AND U6530 ( .A(p_input[28041]), .B(p_input[18041]), .Z(n4354) );
  AND U6531 ( .A(p_input[8041]), .B(p_input[38041]), .Z(n4353) );
  AND U6532 ( .A(n4355), .B(n4356), .Z(o[8040]) );
  AND U6533 ( .A(p_input[28040]), .B(p_input[18040]), .Z(n4356) );
  AND U6534 ( .A(p_input[8040]), .B(p_input[38040]), .Z(n4355) );
  AND U6535 ( .A(n4357), .B(n4358), .Z(o[803]) );
  AND U6536 ( .A(p_input[20803]), .B(p_input[10803]), .Z(n4358) );
  AND U6537 ( .A(p_input[803]), .B(p_input[30803]), .Z(n4357) );
  AND U6538 ( .A(n4359), .B(n4360), .Z(o[8039]) );
  AND U6539 ( .A(p_input[28039]), .B(p_input[18039]), .Z(n4360) );
  AND U6540 ( .A(p_input[8039]), .B(p_input[38039]), .Z(n4359) );
  AND U6541 ( .A(n4361), .B(n4362), .Z(o[8038]) );
  AND U6542 ( .A(p_input[28038]), .B(p_input[18038]), .Z(n4362) );
  AND U6543 ( .A(p_input[8038]), .B(p_input[38038]), .Z(n4361) );
  AND U6544 ( .A(n4363), .B(n4364), .Z(o[8037]) );
  AND U6545 ( .A(p_input[28037]), .B(p_input[18037]), .Z(n4364) );
  AND U6546 ( .A(p_input[8037]), .B(p_input[38037]), .Z(n4363) );
  AND U6547 ( .A(n4365), .B(n4366), .Z(o[8036]) );
  AND U6548 ( .A(p_input[28036]), .B(p_input[18036]), .Z(n4366) );
  AND U6549 ( .A(p_input[8036]), .B(p_input[38036]), .Z(n4365) );
  AND U6550 ( .A(n4367), .B(n4368), .Z(o[8035]) );
  AND U6551 ( .A(p_input[28035]), .B(p_input[18035]), .Z(n4368) );
  AND U6552 ( .A(p_input[8035]), .B(p_input[38035]), .Z(n4367) );
  AND U6553 ( .A(n4369), .B(n4370), .Z(o[8034]) );
  AND U6554 ( .A(p_input[28034]), .B(p_input[18034]), .Z(n4370) );
  AND U6555 ( .A(p_input[8034]), .B(p_input[38034]), .Z(n4369) );
  AND U6556 ( .A(n4371), .B(n4372), .Z(o[8033]) );
  AND U6557 ( .A(p_input[28033]), .B(p_input[18033]), .Z(n4372) );
  AND U6558 ( .A(p_input[8033]), .B(p_input[38033]), .Z(n4371) );
  AND U6559 ( .A(n4373), .B(n4374), .Z(o[8032]) );
  AND U6560 ( .A(p_input[28032]), .B(p_input[18032]), .Z(n4374) );
  AND U6561 ( .A(p_input[8032]), .B(p_input[38032]), .Z(n4373) );
  AND U6562 ( .A(n4375), .B(n4376), .Z(o[8031]) );
  AND U6563 ( .A(p_input[28031]), .B(p_input[18031]), .Z(n4376) );
  AND U6564 ( .A(p_input[8031]), .B(p_input[38031]), .Z(n4375) );
  AND U6565 ( .A(n4377), .B(n4378), .Z(o[8030]) );
  AND U6566 ( .A(p_input[28030]), .B(p_input[18030]), .Z(n4378) );
  AND U6567 ( .A(p_input[8030]), .B(p_input[38030]), .Z(n4377) );
  AND U6568 ( .A(n4379), .B(n4380), .Z(o[802]) );
  AND U6569 ( .A(p_input[20802]), .B(p_input[10802]), .Z(n4380) );
  AND U6570 ( .A(p_input[802]), .B(p_input[30802]), .Z(n4379) );
  AND U6571 ( .A(n4381), .B(n4382), .Z(o[8029]) );
  AND U6572 ( .A(p_input[28029]), .B(p_input[18029]), .Z(n4382) );
  AND U6573 ( .A(p_input[8029]), .B(p_input[38029]), .Z(n4381) );
  AND U6574 ( .A(n4383), .B(n4384), .Z(o[8028]) );
  AND U6575 ( .A(p_input[28028]), .B(p_input[18028]), .Z(n4384) );
  AND U6576 ( .A(p_input[8028]), .B(p_input[38028]), .Z(n4383) );
  AND U6577 ( .A(n4385), .B(n4386), .Z(o[8027]) );
  AND U6578 ( .A(p_input[28027]), .B(p_input[18027]), .Z(n4386) );
  AND U6579 ( .A(p_input[8027]), .B(p_input[38027]), .Z(n4385) );
  AND U6580 ( .A(n4387), .B(n4388), .Z(o[8026]) );
  AND U6581 ( .A(p_input[28026]), .B(p_input[18026]), .Z(n4388) );
  AND U6582 ( .A(p_input[8026]), .B(p_input[38026]), .Z(n4387) );
  AND U6583 ( .A(n4389), .B(n4390), .Z(o[8025]) );
  AND U6584 ( .A(p_input[28025]), .B(p_input[18025]), .Z(n4390) );
  AND U6585 ( .A(p_input[8025]), .B(p_input[38025]), .Z(n4389) );
  AND U6586 ( .A(n4391), .B(n4392), .Z(o[8024]) );
  AND U6587 ( .A(p_input[28024]), .B(p_input[18024]), .Z(n4392) );
  AND U6588 ( .A(p_input[8024]), .B(p_input[38024]), .Z(n4391) );
  AND U6589 ( .A(n4393), .B(n4394), .Z(o[8023]) );
  AND U6590 ( .A(p_input[28023]), .B(p_input[18023]), .Z(n4394) );
  AND U6591 ( .A(p_input[8023]), .B(p_input[38023]), .Z(n4393) );
  AND U6592 ( .A(n4395), .B(n4396), .Z(o[8022]) );
  AND U6593 ( .A(p_input[28022]), .B(p_input[18022]), .Z(n4396) );
  AND U6594 ( .A(p_input[8022]), .B(p_input[38022]), .Z(n4395) );
  AND U6595 ( .A(n4397), .B(n4398), .Z(o[8021]) );
  AND U6596 ( .A(p_input[28021]), .B(p_input[18021]), .Z(n4398) );
  AND U6597 ( .A(p_input[8021]), .B(p_input[38021]), .Z(n4397) );
  AND U6598 ( .A(n4399), .B(n4400), .Z(o[8020]) );
  AND U6599 ( .A(p_input[28020]), .B(p_input[18020]), .Z(n4400) );
  AND U6600 ( .A(p_input[8020]), .B(p_input[38020]), .Z(n4399) );
  AND U6601 ( .A(n4401), .B(n4402), .Z(o[801]) );
  AND U6602 ( .A(p_input[20801]), .B(p_input[10801]), .Z(n4402) );
  AND U6603 ( .A(p_input[801]), .B(p_input[30801]), .Z(n4401) );
  AND U6604 ( .A(n4403), .B(n4404), .Z(o[8019]) );
  AND U6605 ( .A(p_input[28019]), .B(p_input[18019]), .Z(n4404) );
  AND U6606 ( .A(p_input[8019]), .B(p_input[38019]), .Z(n4403) );
  AND U6607 ( .A(n4405), .B(n4406), .Z(o[8018]) );
  AND U6608 ( .A(p_input[28018]), .B(p_input[18018]), .Z(n4406) );
  AND U6609 ( .A(p_input[8018]), .B(p_input[38018]), .Z(n4405) );
  AND U6610 ( .A(n4407), .B(n4408), .Z(o[8017]) );
  AND U6611 ( .A(p_input[28017]), .B(p_input[18017]), .Z(n4408) );
  AND U6612 ( .A(p_input[8017]), .B(p_input[38017]), .Z(n4407) );
  AND U6613 ( .A(n4409), .B(n4410), .Z(o[8016]) );
  AND U6614 ( .A(p_input[28016]), .B(p_input[18016]), .Z(n4410) );
  AND U6615 ( .A(p_input[8016]), .B(p_input[38016]), .Z(n4409) );
  AND U6616 ( .A(n4411), .B(n4412), .Z(o[8015]) );
  AND U6617 ( .A(p_input[28015]), .B(p_input[18015]), .Z(n4412) );
  AND U6618 ( .A(p_input[8015]), .B(p_input[38015]), .Z(n4411) );
  AND U6619 ( .A(n4413), .B(n4414), .Z(o[8014]) );
  AND U6620 ( .A(p_input[28014]), .B(p_input[18014]), .Z(n4414) );
  AND U6621 ( .A(p_input[8014]), .B(p_input[38014]), .Z(n4413) );
  AND U6622 ( .A(n4415), .B(n4416), .Z(o[8013]) );
  AND U6623 ( .A(p_input[28013]), .B(p_input[18013]), .Z(n4416) );
  AND U6624 ( .A(p_input[8013]), .B(p_input[38013]), .Z(n4415) );
  AND U6625 ( .A(n4417), .B(n4418), .Z(o[8012]) );
  AND U6626 ( .A(p_input[28012]), .B(p_input[18012]), .Z(n4418) );
  AND U6627 ( .A(p_input[8012]), .B(p_input[38012]), .Z(n4417) );
  AND U6628 ( .A(n4419), .B(n4420), .Z(o[8011]) );
  AND U6629 ( .A(p_input[28011]), .B(p_input[18011]), .Z(n4420) );
  AND U6630 ( .A(p_input[8011]), .B(p_input[38011]), .Z(n4419) );
  AND U6631 ( .A(n4421), .B(n4422), .Z(o[8010]) );
  AND U6632 ( .A(p_input[28010]), .B(p_input[18010]), .Z(n4422) );
  AND U6633 ( .A(p_input[8010]), .B(p_input[38010]), .Z(n4421) );
  AND U6634 ( .A(n4423), .B(n4424), .Z(o[800]) );
  AND U6635 ( .A(p_input[20800]), .B(p_input[10800]), .Z(n4424) );
  AND U6636 ( .A(p_input[800]), .B(p_input[30800]), .Z(n4423) );
  AND U6637 ( .A(n4425), .B(n4426), .Z(o[8009]) );
  AND U6638 ( .A(p_input[28009]), .B(p_input[18009]), .Z(n4426) );
  AND U6639 ( .A(p_input[8009]), .B(p_input[38009]), .Z(n4425) );
  AND U6640 ( .A(n4427), .B(n4428), .Z(o[8008]) );
  AND U6641 ( .A(p_input[28008]), .B(p_input[18008]), .Z(n4428) );
  AND U6642 ( .A(p_input[8008]), .B(p_input[38008]), .Z(n4427) );
  AND U6643 ( .A(n4429), .B(n4430), .Z(o[8007]) );
  AND U6644 ( .A(p_input[28007]), .B(p_input[18007]), .Z(n4430) );
  AND U6645 ( .A(p_input[8007]), .B(p_input[38007]), .Z(n4429) );
  AND U6646 ( .A(n4431), .B(n4432), .Z(o[8006]) );
  AND U6647 ( .A(p_input[28006]), .B(p_input[18006]), .Z(n4432) );
  AND U6648 ( .A(p_input[8006]), .B(p_input[38006]), .Z(n4431) );
  AND U6649 ( .A(n4433), .B(n4434), .Z(o[8005]) );
  AND U6650 ( .A(p_input[28005]), .B(p_input[18005]), .Z(n4434) );
  AND U6651 ( .A(p_input[8005]), .B(p_input[38005]), .Z(n4433) );
  AND U6652 ( .A(n4435), .B(n4436), .Z(o[8004]) );
  AND U6653 ( .A(p_input[28004]), .B(p_input[18004]), .Z(n4436) );
  AND U6654 ( .A(p_input[8004]), .B(p_input[38004]), .Z(n4435) );
  AND U6655 ( .A(n4437), .B(n4438), .Z(o[8003]) );
  AND U6656 ( .A(p_input[28003]), .B(p_input[18003]), .Z(n4438) );
  AND U6657 ( .A(p_input[8003]), .B(p_input[38003]), .Z(n4437) );
  AND U6658 ( .A(n4439), .B(n4440), .Z(o[8002]) );
  AND U6659 ( .A(p_input[28002]), .B(p_input[18002]), .Z(n4440) );
  AND U6660 ( .A(p_input[8002]), .B(p_input[38002]), .Z(n4439) );
  AND U6661 ( .A(n4441), .B(n4442), .Z(o[8001]) );
  AND U6662 ( .A(p_input[28001]), .B(p_input[18001]), .Z(n4442) );
  AND U6663 ( .A(p_input[8001]), .B(p_input[38001]), .Z(n4441) );
  AND U6664 ( .A(n4443), .B(n4444), .Z(o[8000]) );
  AND U6665 ( .A(p_input[28000]), .B(p_input[18000]), .Z(n4444) );
  AND U6666 ( .A(p_input[8000]), .B(p_input[38000]), .Z(n4443) );
  AND U6667 ( .A(n4445), .B(n4446), .Z(o[7]) );
  AND U6668 ( .A(p_input[20007]), .B(p_input[10007]), .Z(n4446) );
  AND U6669 ( .A(p_input[7]), .B(p_input[30007]), .Z(n4445) );
  AND U6670 ( .A(n4447), .B(n4448), .Z(o[79]) );
  AND U6671 ( .A(p_input[20079]), .B(p_input[10079]), .Z(n4448) );
  AND U6672 ( .A(p_input[79]), .B(p_input[30079]), .Z(n4447) );
  AND U6673 ( .A(n4449), .B(n4450), .Z(o[799]) );
  AND U6674 ( .A(p_input[20799]), .B(p_input[10799]), .Z(n4450) );
  AND U6675 ( .A(p_input[799]), .B(p_input[30799]), .Z(n4449) );
  AND U6676 ( .A(n4451), .B(n4452), .Z(o[7999]) );
  AND U6677 ( .A(p_input[27999]), .B(p_input[17999]), .Z(n4452) );
  AND U6678 ( .A(p_input[7999]), .B(p_input[37999]), .Z(n4451) );
  AND U6679 ( .A(n4453), .B(n4454), .Z(o[7998]) );
  AND U6680 ( .A(p_input[27998]), .B(p_input[17998]), .Z(n4454) );
  AND U6681 ( .A(p_input[7998]), .B(p_input[37998]), .Z(n4453) );
  AND U6682 ( .A(n4455), .B(n4456), .Z(o[7997]) );
  AND U6683 ( .A(p_input[27997]), .B(p_input[17997]), .Z(n4456) );
  AND U6684 ( .A(p_input[7997]), .B(p_input[37997]), .Z(n4455) );
  AND U6685 ( .A(n4457), .B(n4458), .Z(o[7996]) );
  AND U6686 ( .A(p_input[27996]), .B(p_input[17996]), .Z(n4458) );
  AND U6687 ( .A(p_input[7996]), .B(p_input[37996]), .Z(n4457) );
  AND U6688 ( .A(n4459), .B(n4460), .Z(o[7995]) );
  AND U6689 ( .A(p_input[27995]), .B(p_input[17995]), .Z(n4460) );
  AND U6690 ( .A(p_input[7995]), .B(p_input[37995]), .Z(n4459) );
  AND U6691 ( .A(n4461), .B(n4462), .Z(o[7994]) );
  AND U6692 ( .A(p_input[27994]), .B(p_input[17994]), .Z(n4462) );
  AND U6693 ( .A(p_input[7994]), .B(p_input[37994]), .Z(n4461) );
  AND U6694 ( .A(n4463), .B(n4464), .Z(o[7993]) );
  AND U6695 ( .A(p_input[27993]), .B(p_input[17993]), .Z(n4464) );
  AND U6696 ( .A(p_input[7993]), .B(p_input[37993]), .Z(n4463) );
  AND U6697 ( .A(n4465), .B(n4466), .Z(o[7992]) );
  AND U6698 ( .A(p_input[27992]), .B(p_input[17992]), .Z(n4466) );
  AND U6699 ( .A(p_input[7992]), .B(p_input[37992]), .Z(n4465) );
  AND U6700 ( .A(n4467), .B(n4468), .Z(o[7991]) );
  AND U6701 ( .A(p_input[27991]), .B(p_input[17991]), .Z(n4468) );
  AND U6702 ( .A(p_input[7991]), .B(p_input[37991]), .Z(n4467) );
  AND U6703 ( .A(n4469), .B(n4470), .Z(o[7990]) );
  AND U6704 ( .A(p_input[27990]), .B(p_input[17990]), .Z(n4470) );
  AND U6705 ( .A(p_input[7990]), .B(p_input[37990]), .Z(n4469) );
  AND U6706 ( .A(n4471), .B(n4472), .Z(o[798]) );
  AND U6707 ( .A(p_input[20798]), .B(p_input[10798]), .Z(n4472) );
  AND U6708 ( .A(p_input[798]), .B(p_input[30798]), .Z(n4471) );
  AND U6709 ( .A(n4473), .B(n4474), .Z(o[7989]) );
  AND U6710 ( .A(p_input[27989]), .B(p_input[17989]), .Z(n4474) );
  AND U6711 ( .A(p_input[7989]), .B(p_input[37989]), .Z(n4473) );
  AND U6712 ( .A(n4475), .B(n4476), .Z(o[7988]) );
  AND U6713 ( .A(p_input[27988]), .B(p_input[17988]), .Z(n4476) );
  AND U6714 ( .A(p_input[7988]), .B(p_input[37988]), .Z(n4475) );
  AND U6715 ( .A(n4477), .B(n4478), .Z(o[7987]) );
  AND U6716 ( .A(p_input[27987]), .B(p_input[17987]), .Z(n4478) );
  AND U6717 ( .A(p_input[7987]), .B(p_input[37987]), .Z(n4477) );
  AND U6718 ( .A(n4479), .B(n4480), .Z(o[7986]) );
  AND U6719 ( .A(p_input[27986]), .B(p_input[17986]), .Z(n4480) );
  AND U6720 ( .A(p_input[7986]), .B(p_input[37986]), .Z(n4479) );
  AND U6721 ( .A(n4481), .B(n4482), .Z(o[7985]) );
  AND U6722 ( .A(p_input[27985]), .B(p_input[17985]), .Z(n4482) );
  AND U6723 ( .A(p_input[7985]), .B(p_input[37985]), .Z(n4481) );
  AND U6724 ( .A(n4483), .B(n4484), .Z(o[7984]) );
  AND U6725 ( .A(p_input[27984]), .B(p_input[17984]), .Z(n4484) );
  AND U6726 ( .A(p_input[7984]), .B(p_input[37984]), .Z(n4483) );
  AND U6727 ( .A(n4485), .B(n4486), .Z(o[7983]) );
  AND U6728 ( .A(p_input[27983]), .B(p_input[17983]), .Z(n4486) );
  AND U6729 ( .A(p_input[7983]), .B(p_input[37983]), .Z(n4485) );
  AND U6730 ( .A(n4487), .B(n4488), .Z(o[7982]) );
  AND U6731 ( .A(p_input[27982]), .B(p_input[17982]), .Z(n4488) );
  AND U6732 ( .A(p_input[7982]), .B(p_input[37982]), .Z(n4487) );
  AND U6733 ( .A(n4489), .B(n4490), .Z(o[7981]) );
  AND U6734 ( .A(p_input[27981]), .B(p_input[17981]), .Z(n4490) );
  AND U6735 ( .A(p_input[7981]), .B(p_input[37981]), .Z(n4489) );
  AND U6736 ( .A(n4491), .B(n4492), .Z(o[7980]) );
  AND U6737 ( .A(p_input[27980]), .B(p_input[17980]), .Z(n4492) );
  AND U6738 ( .A(p_input[7980]), .B(p_input[37980]), .Z(n4491) );
  AND U6739 ( .A(n4493), .B(n4494), .Z(o[797]) );
  AND U6740 ( .A(p_input[20797]), .B(p_input[10797]), .Z(n4494) );
  AND U6741 ( .A(p_input[797]), .B(p_input[30797]), .Z(n4493) );
  AND U6742 ( .A(n4495), .B(n4496), .Z(o[7979]) );
  AND U6743 ( .A(p_input[27979]), .B(p_input[17979]), .Z(n4496) );
  AND U6744 ( .A(p_input[7979]), .B(p_input[37979]), .Z(n4495) );
  AND U6745 ( .A(n4497), .B(n4498), .Z(o[7978]) );
  AND U6746 ( .A(p_input[27978]), .B(p_input[17978]), .Z(n4498) );
  AND U6747 ( .A(p_input[7978]), .B(p_input[37978]), .Z(n4497) );
  AND U6748 ( .A(n4499), .B(n4500), .Z(o[7977]) );
  AND U6749 ( .A(p_input[27977]), .B(p_input[17977]), .Z(n4500) );
  AND U6750 ( .A(p_input[7977]), .B(p_input[37977]), .Z(n4499) );
  AND U6751 ( .A(n4501), .B(n4502), .Z(o[7976]) );
  AND U6752 ( .A(p_input[27976]), .B(p_input[17976]), .Z(n4502) );
  AND U6753 ( .A(p_input[7976]), .B(p_input[37976]), .Z(n4501) );
  AND U6754 ( .A(n4503), .B(n4504), .Z(o[7975]) );
  AND U6755 ( .A(p_input[27975]), .B(p_input[17975]), .Z(n4504) );
  AND U6756 ( .A(p_input[7975]), .B(p_input[37975]), .Z(n4503) );
  AND U6757 ( .A(n4505), .B(n4506), .Z(o[7974]) );
  AND U6758 ( .A(p_input[27974]), .B(p_input[17974]), .Z(n4506) );
  AND U6759 ( .A(p_input[7974]), .B(p_input[37974]), .Z(n4505) );
  AND U6760 ( .A(n4507), .B(n4508), .Z(o[7973]) );
  AND U6761 ( .A(p_input[27973]), .B(p_input[17973]), .Z(n4508) );
  AND U6762 ( .A(p_input[7973]), .B(p_input[37973]), .Z(n4507) );
  AND U6763 ( .A(n4509), .B(n4510), .Z(o[7972]) );
  AND U6764 ( .A(p_input[27972]), .B(p_input[17972]), .Z(n4510) );
  AND U6765 ( .A(p_input[7972]), .B(p_input[37972]), .Z(n4509) );
  AND U6766 ( .A(n4511), .B(n4512), .Z(o[7971]) );
  AND U6767 ( .A(p_input[27971]), .B(p_input[17971]), .Z(n4512) );
  AND U6768 ( .A(p_input[7971]), .B(p_input[37971]), .Z(n4511) );
  AND U6769 ( .A(n4513), .B(n4514), .Z(o[7970]) );
  AND U6770 ( .A(p_input[27970]), .B(p_input[17970]), .Z(n4514) );
  AND U6771 ( .A(p_input[7970]), .B(p_input[37970]), .Z(n4513) );
  AND U6772 ( .A(n4515), .B(n4516), .Z(o[796]) );
  AND U6773 ( .A(p_input[20796]), .B(p_input[10796]), .Z(n4516) );
  AND U6774 ( .A(p_input[796]), .B(p_input[30796]), .Z(n4515) );
  AND U6775 ( .A(n4517), .B(n4518), .Z(o[7969]) );
  AND U6776 ( .A(p_input[27969]), .B(p_input[17969]), .Z(n4518) );
  AND U6777 ( .A(p_input[7969]), .B(p_input[37969]), .Z(n4517) );
  AND U6778 ( .A(n4519), .B(n4520), .Z(o[7968]) );
  AND U6779 ( .A(p_input[27968]), .B(p_input[17968]), .Z(n4520) );
  AND U6780 ( .A(p_input[7968]), .B(p_input[37968]), .Z(n4519) );
  AND U6781 ( .A(n4521), .B(n4522), .Z(o[7967]) );
  AND U6782 ( .A(p_input[27967]), .B(p_input[17967]), .Z(n4522) );
  AND U6783 ( .A(p_input[7967]), .B(p_input[37967]), .Z(n4521) );
  AND U6784 ( .A(n4523), .B(n4524), .Z(o[7966]) );
  AND U6785 ( .A(p_input[27966]), .B(p_input[17966]), .Z(n4524) );
  AND U6786 ( .A(p_input[7966]), .B(p_input[37966]), .Z(n4523) );
  AND U6787 ( .A(n4525), .B(n4526), .Z(o[7965]) );
  AND U6788 ( .A(p_input[27965]), .B(p_input[17965]), .Z(n4526) );
  AND U6789 ( .A(p_input[7965]), .B(p_input[37965]), .Z(n4525) );
  AND U6790 ( .A(n4527), .B(n4528), .Z(o[7964]) );
  AND U6791 ( .A(p_input[27964]), .B(p_input[17964]), .Z(n4528) );
  AND U6792 ( .A(p_input[7964]), .B(p_input[37964]), .Z(n4527) );
  AND U6793 ( .A(n4529), .B(n4530), .Z(o[7963]) );
  AND U6794 ( .A(p_input[27963]), .B(p_input[17963]), .Z(n4530) );
  AND U6795 ( .A(p_input[7963]), .B(p_input[37963]), .Z(n4529) );
  AND U6796 ( .A(n4531), .B(n4532), .Z(o[7962]) );
  AND U6797 ( .A(p_input[27962]), .B(p_input[17962]), .Z(n4532) );
  AND U6798 ( .A(p_input[7962]), .B(p_input[37962]), .Z(n4531) );
  AND U6799 ( .A(n4533), .B(n4534), .Z(o[7961]) );
  AND U6800 ( .A(p_input[27961]), .B(p_input[17961]), .Z(n4534) );
  AND U6801 ( .A(p_input[7961]), .B(p_input[37961]), .Z(n4533) );
  AND U6802 ( .A(n4535), .B(n4536), .Z(o[7960]) );
  AND U6803 ( .A(p_input[27960]), .B(p_input[17960]), .Z(n4536) );
  AND U6804 ( .A(p_input[7960]), .B(p_input[37960]), .Z(n4535) );
  AND U6805 ( .A(n4537), .B(n4538), .Z(o[795]) );
  AND U6806 ( .A(p_input[20795]), .B(p_input[10795]), .Z(n4538) );
  AND U6807 ( .A(p_input[795]), .B(p_input[30795]), .Z(n4537) );
  AND U6808 ( .A(n4539), .B(n4540), .Z(o[7959]) );
  AND U6809 ( .A(p_input[27959]), .B(p_input[17959]), .Z(n4540) );
  AND U6810 ( .A(p_input[7959]), .B(p_input[37959]), .Z(n4539) );
  AND U6811 ( .A(n4541), .B(n4542), .Z(o[7958]) );
  AND U6812 ( .A(p_input[27958]), .B(p_input[17958]), .Z(n4542) );
  AND U6813 ( .A(p_input[7958]), .B(p_input[37958]), .Z(n4541) );
  AND U6814 ( .A(n4543), .B(n4544), .Z(o[7957]) );
  AND U6815 ( .A(p_input[27957]), .B(p_input[17957]), .Z(n4544) );
  AND U6816 ( .A(p_input[7957]), .B(p_input[37957]), .Z(n4543) );
  AND U6817 ( .A(n4545), .B(n4546), .Z(o[7956]) );
  AND U6818 ( .A(p_input[27956]), .B(p_input[17956]), .Z(n4546) );
  AND U6819 ( .A(p_input[7956]), .B(p_input[37956]), .Z(n4545) );
  AND U6820 ( .A(n4547), .B(n4548), .Z(o[7955]) );
  AND U6821 ( .A(p_input[27955]), .B(p_input[17955]), .Z(n4548) );
  AND U6822 ( .A(p_input[7955]), .B(p_input[37955]), .Z(n4547) );
  AND U6823 ( .A(n4549), .B(n4550), .Z(o[7954]) );
  AND U6824 ( .A(p_input[27954]), .B(p_input[17954]), .Z(n4550) );
  AND U6825 ( .A(p_input[7954]), .B(p_input[37954]), .Z(n4549) );
  AND U6826 ( .A(n4551), .B(n4552), .Z(o[7953]) );
  AND U6827 ( .A(p_input[27953]), .B(p_input[17953]), .Z(n4552) );
  AND U6828 ( .A(p_input[7953]), .B(p_input[37953]), .Z(n4551) );
  AND U6829 ( .A(n4553), .B(n4554), .Z(o[7952]) );
  AND U6830 ( .A(p_input[27952]), .B(p_input[17952]), .Z(n4554) );
  AND U6831 ( .A(p_input[7952]), .B(p_input[37952]), .Z(n4553) );
  AND U6832 ( .A(n4555), .B(n4556), .Z(o[7951]) );
  AND U6833 ( .A(p_input[27951]), .B(p_input[17951]), .Z(n4556) );
  AND U6834 ( .A(p_input[7951]), .B(p_input[37951]), .Z(n4555) );
  AND U6835 ( .A(n4557), .B(n4558), .Z(o[7950]) );
  AND U6836 ( .A(p_input[27950]), .B(p_input[17950]), .Z(n4558) );
  AND U6837 ( .A(p_input[7950]), .B(p_input[37950]), .Z(n4557) );
  AND U6838 ( .A(n4559), .B(n4560), .Z(o[794]) );
  AND U6839 ( .A(p_input[20794]), .B(p_input[10794]), .Z(n4560) );
  AND U6840 ( .A(p_input[794]), .B(p_input[30794]), .Z(n4559) );
  AND U6841 ( .A(n4561), .B(n4562), .Z(o[7949]) );
  AND U6842 ( .A(p_input[27949]), .B(p_input[17949]), .Z(n4562) );
  AND U6843 ( .A(p_input[7949]), .B(p_input[37949]), .Z(n4561) );
  AND U6844 ( .A(n4563), .B(n4564), .Z(o[7948]) );
  AND U6845 ( .A(p_input[27948]), .B(p_input[17948]), .Z(n4564) );
  AND U6846 ( .A(p_input[7948]), .B(p_input[37948]), .Z(n4563) );
  AND U6847 ( .A(n4565), .B(n4566), .Z(o[7947]) );
  AND U6848 ( .A(p_input[27947]), .B(p_input[17947]), .Z(n4566) );
  AND U6849 ( .A(p_input[7947]), .B(p_input[37947]), .Z(n4565) );
  AND U6850 ( .A(n4567), .B(n4568), .Z(o[7946]) );
  AND U6851 ( .A(p_input[27946]), .B(p_input[17946]), .Z(n4568) );
  AND U6852 ( .A(p_input[7946]), .B(p_input[37946]), .Z(n4567) );
  AND U6853 ( .A(n4569), .B(n4570), .Z(o[7945]) );
  AND U6854 ( .A(p_input[27945]), .B(p_input[17945]), .Z(n4570) );
  AND U6855 ( .A(p_input[7945]), .B(p_input[37945]), .Z(n4569) );
  AND U6856 ( .A(n4571), .B(n4572), .Z(o[7944]) );
  AND U6857 ( .A(p_input[27944]), .B(p_input[17944]), .Z(n4572) );
  AND U6858 ( .A(p_input[7944]), .B(p_input[37944]), .Z(n4571) );
  AND U6859 ( .A(n4573), .B(n4574), .Z(o[7943]) );
  AND U6860 ( .A(p_input[27943]), .B(p_input[17943]), .Z(n4574) );
  AND U6861 ( .A(p_input[7943]), .B(p_input[37943]), .Z(n4573) );
  AND U6862 ( .A(n4575), .B(n4576), .Z(o[7942]) );
  AND U6863 ( .A(p_input[27942]), .B(p_input[17942]), .Z(n4576) );
  AND U6864 ( .A(p_input[7942]), .B(p_input[37942]), .Z(n4575) );
  AND U6865 ( .A(n4577), .B(n4578), .Z(o[7941]) );
  AND U6866 ( .A(p_input[27941]), .B(p_input[17941]), .Z(n4578) );
  AND U6867 ( .A(p_input[7941]), .B(p_input[37941]), .Z(n4577) );
  AND U6868 ( .A(n4579), .B(n4580), .Z(o[7940]) );
  AND U6869 ( .A(p_input[27940]), .B(p_input[17940]), .Z(n4580) );
  AND U6870 ( .A(p_input[7940]), .B(p_input[37940]), .Z(n4579) );
  AND U6871 ( .A(n4581), .B(n4582), .Z(o[793]) );
  AND U6872 ( .A(p_input[20793]), .B(p_input[10793]), .Z(n4582) );
  AND U6873 ( .A(p_input[793]), .B(p_input[30793]), .Z(n4581) );
  AND U6874 ( .A(n4583), .B(n4584), .Z(o[7939]) );
  AND U6875 ( .A(p_input[27939]), .B(p_input[17939]), .Z(n4584) );
  AND U6876 ( .A(p_input[7939]), .B(p_input[37939]), .Z(n4583) );
  AND U6877 ( .A(n4585), .B(n4586), .Z(o[7938]) );
  AND U6878 ( .A(p_input[27938]), .B(p_input[17938]), .Z(n4586) );
  AND U6879 ( .A(p_input[7938]), .B(p_input[37938]), .Z(n4585) );
  AND U6880 ( .A(n4587), .B(n4588), .Z(o[7937]) );
  AND U6881 ( .A(p_input[27937]), .B(p_input[17937]), .Z(n4588) );
  AND U6882 ( .A(p_input[7937]), .B(p_input[37937]), .Z(n4587) );
  AND U6883 ( .A(n4589), .B(n4590), .Z(o[7936]) );
  AND U6884 ( .A(p_input[27936]), .B(p_input[17936]), .Z(n4590) );
  AND U6885 ( .A(p_input[7936]), .B(p_input[37936]), .Z(n4589) );
  AND U6886 ( .A(n4591), .B(n4592), .Z(o[7935]) );
  AND U6887 ( .A(p_input[27935]), .B(p_input[17935]), .Z(n4592) );
  AND U6888 ( .A(p_input[7935]), .B(p_input[37935]), .Z(n4591) );
  AND U6889 ( .A(n4593), .B(n4594), .Z(o[7934]) );
  AND U6890 ( .A(p_input[27934]), .B(p_input[17934]), .Z(n4594) );
  AND U6891 ( .A(p_input[7934]), .B(p_input[37934]), .Z(n4593) );
  AND U6892 ( .A(n4595), .B(n4596), .Z(o[7933]) );
  AND U6893 ( .A(p_input[27933]), .B(p_input[17933]), .Z(n4596) );
  AND U6894 ( .A(p_input[7933]), .B(p_input[37933]), .Z(n4595) );
  AND U6895 ( .A(n4597), .B(n4598), .Z(o[7932]) );
  AND U6896 ( .A(p_input[27932]), .B(p_input[17932]), .Z(n4598) );
  AND U6897 ( .A(p_input[7932]), .B(p_input[37932]), .Z(n4597) );
  AND U6898 ( .A(n4599), .B(n4600), .Z(o[7931]) );
  AND U6899 ( .A(p_input[27931]), .B(p_input[17931]), .Z(n4600) );
  AND U6900 ( .A(p_input[7931]), .B(p_input[37931]), .Z(n4599) );
  AND U6901 ( .A(n4601), .B(n4602), .Z(o[7930]) );
  AND U6902 ( .A(p_input[27930]), .B(p_input[17930]), .Z(n4602) );
  AND U6903 ( .A(p_input[7930]), .B(p_input[37930]), .Z(n4601) );
  AND U6904 ( .A(n4603), .B(n4604), .Z(o[792]) );
  AND U6905 ( .A(p_input[20792]), .B(p_input[10792]), .Z(n4604) );
  AND U6906 ( .A(p_input[792]), .B(p_input[30792]), .Z(n4603) );
  AND U6907 ( .A(n4605), .B(n4606), .Z(o[7929]) );
  AND U6908 ( .A(p_input[27929]), .B(p_input[17929]), .Z(n4606) );
  AND U6909 ( .A(p_input[7929]), .B(p_input[37929]), .Z(n4605) );
  AND U6910 ( .A(n4607), .B(n4608), .Z(o[7928]) );
  AND U6911 ( .A(p_input[27928]), .B(p_input[17928]), .Z(n4608) );
  AND U6912 ( .A(p_input[7928]), .B(p_input[37928]), .Z(n4607) );
  AND U6913 ( .A(n4609), .B(n4610), .Z(o[7927]) );
  AND U6914 ( .A(p_input[27927]), .B(p_input[17927]), .Z(n4610) );
  AND U6915 ( .A(p_input[7927]), .B(p_input[37927]), .Z(n4609) );
  AND U6916 ( .A(n4611), .B(n4612), .Z(o[7926]) );
  AND U6917 ( .A(p_input[27926]), .B(p_input[17926]), .Z(n4612) );
  AND U6918 ( .A(p_input[7926]), .B(p_input[37926]), .Z(n4611) );
  AND U6919 ( .A(n4613), .B(n4614), .Z(o[7925]) );
  AND U6920 ( .A(p_input[27925]), .B(p_input[17925]), .Z(n4614) );
  AND U6921 ( .A(p_input[7925]), .B(p_input[37925]), .Z(n4613) );
  AND U6922 ( .A(n4615), .B(n4616), .Z(o[7924]) );
  AND U6923 ( .A(p_input[27924]), .B(p_input[17924]), .Z(n4616) );
  AND U6924 ( .A(p_input[7924]), .B(p_input[37924]), .Z(n4615) );
  AND U6925 ( .A(n4617), .B(n4618), .Z(o[7923]) );
  AND U6926 ( .A(p_input[27923]), .B(p_input[17923]), .Z(n4618) );
  AND U6927 ( .A(p_input[7923]), .B(p_input[37923]), .Z(n4617) );
  AND U6928 ( .A(n4619), .B(n4620), .Z(o[7922]) );
  AND U6929 ( .A(p_input[27922]), .B(p_input[17922]), .Z(n4620) );
  AND U6930 ( .A(p_input[7922]), .B(p_input[37922]), .Z(n4619) );
  AND U6931 ( .A(n4621), .B(n4622), .Z(o[7921]) );
  AND U6932 ( .A(p_input[27921]), .B(p_input[17921]), .Z(n4622) );
  AND U6933 ( .A(p_input[7921]), .B(p_input[37921]), .Z(n4621) );
  AND U6934 ( .A(n4623), .B(n4624), .Z(o[7920]) );
  AND U6935 ( .A(p_input[27920]), .B(p_input[17920]), .Z(n4624) );
  AND U6936 ( .A(p_input[7920]), .B(p_input[37920]), .Z(n4623) );
  AND U6937 ( .A(n4625), .B(n4626), .Z(o[791]) );
  AND U6938 ( .A(p_input[20791]), .B(p_input[10791]), .Z(n4626) );
  AND U6939 ( .A(p_input[791]), .B(p_input[30791]), .Z(n4625) );
  AND U6940 ( .A(n4627), .B(n4628), .Z(o[7919]) );
  AND U6941 ( .A(p_input[27919]), .B(p_input[17919]), .Z(n4628) );
  AND U6942 ( .A(p_input[7919]), .B(p_input[37919]), .Z(n4627) );
  AND U6943 ( .A(n4629), .B(n4630), .Z(o[7918]) );
  AND U6944 ( .A(p_input[27918]), .B(p_input[17918]), .Z(n4630) );
  AND U6945 ( .A(p_input[7918]), .B(p_input[37918]), .Z(n4629) );
  AND U6946 ( .A(n4631), .B(n4632), .Z(o[7917]) );
  AND U6947 ( .A(p_input[27917]), .B(p_input[17917]), .Z(n4632) );
  AND U6948 ( .A(p_input[7917]), .B(p_input[37917]), .Z(n4631) );
  AND U6949 ( .A(n4633), .B(n4634), .Z(o[7916]) );
  AND U6950 ( .A(p_input[27916]), .B(p_input[17916]), .Z(n4634) );
  AND U6951 ( .A(p_input[7916]), .B(p_input[37916]), .Z(n4633) );
  AND U6952 ( .A(n4635), .B(n4636), .Z(o[7915]) );
  AND U6953 ( .A(p_input[27915]), .B(p_input[17915]), .Z(n4636) );
  AND U6954 ( .A(p_input[7915]), .B(p_input[37915]), .Z(n4635) );
  AND U6955 ( .A(n4637), .B(n4638), .Z(o[7914]) );
  AND U6956 ( .A(p_input[27914]), .B(p_input[17914]), .Z(n4638) );
  AND U6957 ( .A(p_input[7914]), .B(p_input[37914]), .Z(n4637) );
  AND U6958 ( .A(n4639), .B(n4640), .Z(o[7913]) );
  AND U6959 ( .A(p_input[27913]), .B(p_input[17913]), .Z(n4640) );
  AND U6960 ( .A(p_input[7913]), .B(p_input[37913]), .Z(n4639) );
  AND U6961 ( .A(n4641), .B(n4642), .Z(o[7912]) );
  AND U6962 ( .A(p_input[27912]), .B(p_input[17912]), .Z(n4642) );
  AND U6963 ( .A(p_input[7912]), .B(p_input[37912]), .Z(n4641) );
  AND U6964 ( .A(n4643), .B(n4644), .Z(o[7911]) );
  AND U6965 ( .A(p_input[27911]), .B(p_input[17911]), .Z(n4644) );
  AND U6966 ( .A(p_input[7911]), .B(p_input[37911]), .Z(n4643) );
  AND U6967 ( .A(n4645), .B(n4646), .Z(o[7910]) );
  AND U6968 ( .A(p_input[27910]), .B(p_input[17910]), .Z(n4646) );
  AND U6969 ( .A(p_input[7910]), .B(p_input[37910]), .Z(n4645) );
  AND U6970 ( .A(n4647), .B(n4648), .Z(o[790]) );
  AND U6971 ( .A(p_input[20790]), .B(p_input[10790]), .Z(n4648) );
  AND U6972 ( .A(p_input[790]), .B(p_input[30790]), .Z(n4647) );
  AND U6973 ( .A(n4649), .B(n4650), .Z(o[7909]) );
  AND U6974 ( .A(p_input[27909]), .B(p_input[17909]), .Z(n4650) );
  AND U6975 ( .A(p_input[7909]), .B(p_input[37909]), .Z(n4649) );
  AND U6976 ( .A(n4651), .B(n4652), .Z(o[7908]) );
  AND U6977 ( .A(p_input[27908]), .B(p_input[17908]), .Z(n4652) );
  AND U6978 ( .A(p_input[7908]), .B(p_input[37908]), .Z(n4651) );
  AND U6979 ( .A(n4653), .B(n4654), .Z(o[7907]) );
  AND U6980 ( .A(p_input[27907]), .B(p_input[17907]), .Z(n4654) );
  AND U6981 ( .A(p_input[7907]), .B(p_input[37907]), .Z(n4653) );
  AND U6982 ( .A(n4655), .B(n4656), .Z(o[7906]) );
  AND U6983 ( .A(p_input[27906]), .B(p_input[17906]), .Z(n4656) );
  AND U6984 ( .A(p_input[7906]), .B(p_input[37906]), .Z(n4655) );
  AND U6985 ( .A(n4657), .B(n4658), .Z(o[7905]) );
  AND U6986 ( .A(p_input[27905]), .B(p_input[17905]), .Z(n4658) );
  AND U6987 ( .A(p_input[7905]), .B(p_input[37905]), .Z(n4657) );
  AND U6988 ( .A(n4659), .B(n4660), .Z(o[7904]) );
  AND U6989 ( .A(p_input[27904]), .B(p_input[17904]), .Z(n4660) );
  AND U6990 ( .A(p_input[7904]), .B(p_input[37904]), .Z(n4659) );
  AND U6991 ( .A(n4661), .B(n4662), .Z(o[7903]) );
  AND U6992 ( .A(p_input[27903]), .B(p_input[17903]), .Z(n4662) );
  AND U6993 ( .A(p_input[7903]), .B(p_input[37903]), .Z(n4661) );
  AND U6994 ( .A(n4663), .B(n4664), .Z(o[7902]) );
  AND U6995 ( .A(p_input[27902]), .B(p_input[17902]), .Z(n4664) );
  AND U6996 ( .A(p_input[7902]), .B(p_input[37902]), .Z(n4663) );
  AND U6997 ( .A(n4665), .B(n4666), .Z(o[7901]) );
  AND U6998 ( .A(p_input[27901]), .B(p_input[17901]), .Z(n4666) );
  AND U6999 ( .A(p_input[7901]), .B(p_input[37901]), .Z(n4665) );
  AND U7000 ( .A(n4667), .B(n4668), .Z(o[7900]) );
  AND U7001 ( .A(p_input[27900]), .B(p_input[17900]), .Z(n4668) );
  AND U7002 ( .A(p_input[7900]), .B(p_input[37900]), .Z(n4667) );
  AND U7003 ( .A(n4669), .B(n4670), .Z(o[78]) );
  AND U7004 ( .A(p_input[20078]), .B(p_input[10078]), .Z(n4670) );
  AND U7005 ( .A(p_input[78]), .B(p_input[30078]), .Z(n4669) );
  AND U7006 ( .A(n4671), .B(n4672), .Z(o[789]) );
  AND U7007 ( .A(p_input[20789]), .B(p_input[10789]), .Z(n4672) );
  AND U7008 ( .A(p_input[789]), .B(p_input[30789]), .Z(n4671) );
  AND U7009 ( .A(n4673), .B(n4674), .Z(o[7899]) );
  AND U7010 ( .A(p_input[27899]), .B(p_input[17899]), .Z(n4674) );
  AND U7011 ( .A(p_input[7899]), .B(p_input[37899]), .Z(n4673) );
  AND U7012 ( .A(n4675), .B(n4676), .Z(o[7898]) );
  AND U7013 ( .A(p_input[27898]), .B(p_input[17898]), .Z(n4676) );
  AND U7014 ( .A(p_input[7898]), .B(p_input[37898]), .Z(n4675) );
  AND U7015 ( .A(n4677), .B(n4678), .Z(o[7897]) );
  AND U7016 ( .A(p_input[27897]), .B(p_input[17897]), .Z(n4678) );
  AND U7017 ( .A(p_input[7897]), .B(p_input[37897]), .Z(n4677) );
  AND U7018 ( .A(n4679), .B(n4680), .Z(o[7896]) );
  AND U7019 ( .A(p_input[27896]), .B(p_input[17896]), .Z(n4680) );
  AND U7020 ( .A(p_input[7896]), .B(p_input[37896]), .Z(n4679) );
  AND U7021 ( .A(n4681), .B(n4682), .Z(o[7895]) );
  AND U7022 ( .A(p_input[27895]), .B(p_input[17895]), .Z(n4682) );
  AND U7023 ( .A(p_input[7895]), .B(p_input[37895]), .Z(n4681) );
  AND U7024 ( .A(n4683), .B(n4684), .Z(o[7894]) );
  AND U7025 ( .A(p_input[27894]), .B(p_input[17894]), .Z(n4684) );
  AND U7026 ( .A(p_input[7894]), .B(p_input[37894]), .Z(n4683) );
  AND U7027 ( .A(n4685), .B(n4686), .Z(o[7893]) );
  AND U7028 ( .A(p_input[27893]), .B(p_input[17893]), .Z(n4686) );
  AND U7029 ( .A(p_input[7893]), .B(p_input[37893]), .Z(n4685) );
  AND U7030 ( .A(n4687), .B(n4688), .Z(o[7892]) );
  AND U7031 ( .A(p_input[27892]), .B(p_input[17892]), .Z(n4688) );
  AND U7032 ( .A(p_input[7892]), .B(p_input[37892]), .Z(n4687) );
  AND U7033 ( .A(n4689), .B(n4690), .Z(o[7891]) );
  AND U7034 ( .A(p_input[27891]), .B(p_input[17891]), .Z(n4690) );
  AND U7035 ( .A(p_input[7891]), .B(p_input[37891]), .Z(n4689) );
  AND U7036 ( .A(n4691), .B(n4692), .Z(o[7890]) );
  AND U7037 ( .A(p_input[27890]), .B(p_input[17890]), .Z(n4692) );
  AND U7038 ( .A(p_input[7890]), .B(p_input[37890]), .Z(n4691) );
  AND U7039 ( .A(n4693), .B(n4694), .Z(o[788]) );
  AND U7040 ( .A(p_input[20788]), .B(p_input[10788]), .Z(n4694) );
  AND U7041 ( .A(p_input[788]), .B(p_input[30788]), .Z(n4693) );
  AND U7042 ( .A(n4695), .B(n4696), .Z(o[7889]) );
  AND U7043 ( .A(p_input[27889]), .B(p_input[17889]), .Z(n4696) );
  AND U7044 ( .A(p_input[7889]), .B(p_input[37889]), .Z(n4695) );
  AND U7045 ( .A(n4697), .B(n4698), .Z(o[7888]) );
  AND U7046 ( .A(p_input[27888]), .B(p_input[17888]), .Z(n4698) );
  AND U7047 ( .A(p_input[7888]), .B(p_input[37888]), .Z(n4697) );
  AND U7048 ( .A(n4699), .B(n4700), .Z(o[7887]) );
  AND U7049 ( .A(p_input[27887]), .B(p_input[17887]), .Z(n4700) );
  AND U7050 ( .A(p_input[7887]), .B(p_input[37887]), .Z(n4699) );
  AND U7051 ( .A(n4701), .B(n4702), .Z(o[7886]) );
  AND U7052 ( .A(p_input[27886]), .B(p_input[17886]), .Z(n4702) );
  AND U7053 ( .A(p_input[7886]), .B(p_input[37886]), .Z(n4701) );
  AND U7054 ( .A(n4703), .B(n4704), .Z(o[7885]) );
  AND U7055 ( .A(p_input[27885]), .B(p_input[17885]), .Z(n4704) );
  AND U7056 ( .A(p_input[7885]), .B(p_input[37885]), .Z(n4703) );
  AND U7057 ( .A(n4705), .B(n4706), .Z(o[7884]) );
  AND U7058 ( .A(p_input[27884]), .B(p_input[17884]), .Z(n4706) );
  AND U7059 ( .A(p_input[7884]), .B(p_input[37884]), .Z(n4705) );
  AND U7060 ( .A(n4707), .B(n4708), .Z(o[7883]) );
  AND U7061 ( .A(p_input[27883]), .B(p_input[17883]), .Z(n4708) );
  AND U7062 ( .A(p_input[7883]), .B(p_input[37883]), .Z(n4707) );
  AND U7063 ( .A(n4709), .B(n4710), .Z(o[7882]) );
  AND U7064 ( .A(p_input[27882]), .B(p_input[17882]), .Z(n4710) );
  AND U7065 ( .A(p_input[7882]), .B(p_input[37882]), .Z(n4709) );
  AND U7066 ( .A(n4711), .B(n4712), .Z(o[7881]) );
  AND U7067 ( .A(p_input[27881]), .B(p_input[17881]), .Z(n4712) );
  AND U7068 ( .A(p_input[7881]), .B(p_input[37881]), .Z(n4711) );
  AND U7069 ( .A(n4713), .B(n4714), .Z(o[7880]) );
  AND U7070 ( .A(p_input[27880]), .B(p_input[17880]), .Z(n4714) );
  AND U7071 ( .A(p_input[7880]), .B(p_input[37880]), .Z(n4713) );
  AND U7072 ( .A(n4715), .B(n4716), .Z(o[787]) );
  AND U7073 ( .A(p_input[20787]), .B(p_input[10787]), .Z(n4716) );
  AND U7074 ( .A(p_input[787]), .B(p_input[30787]), .Z(n4715) );
  AND U7075 ( .A(n4717), .B(n4718), .Z(o[7879]) );
  AND U7076 ( .A(p_input[27879]), .B(p_input[17879]), .Z(n4718) );
  AND U7077 ( .A(p_input[7879]), .B(p_input[37879]), .Z(n4717) );
  AND U7078 ( .A(n4719), .B(n4720), .Z(o[7878]) );
  AND U7079 ( .A(p_input[27878]), .B(p_input[17878]), .Z(n4720) );
  AND U7080 ( .A(p_input[7878]), .B(p_input[37878]), .Z(n4719) );
  AND U7081 ( .A(n4721), .B(n4722), .Z(o[7877]) );
  AND U7082 ( .A(p_input[27877]), .B(p_input[17877]), .Z(n4722) );
  AND U7083 ( .A(p_input[7877]), .B(p_input[37877]), .Z(n4721) );
  AND U7084 ( .A(n4723), .B(n4724), .Z(o[7876]) );
  AND U7085 ( .A(p_input[27876]), .B(p_input[17876]), .Z(n4724) );
  AND U7086 ( .A(p_input[7876]), .B(p_input[37876]), .Z(n4723) );
  AND U7087 ( .A(n4725), .B(n4726), .Z(o[7875]) );
  AND U7088 ( .A(p_input[27875]), .B(p_input[17875]), .Z(n4726) );
  AND U7089 ( .A(p_input[7875]), .B(p_input[37875]), .Z(n4725) );
  AND U7090 ( .A(n4727), .B(n4728), .Z(o[7874]) );
  AND U7091 ( .A(p_input[27874]), .B(p_input[17874]), .Z(n4728) );
  AND U7092 ( .A(p_input[7874]), .B(p_input[37874]), .Z(n4727) );
  AND U7093 ( .A(n4729), .B(n4730), .Z(o[7873]) );
  AND U7094 ( .A(p_input[27873]), .B(p_input[17873]), .Z(n4730) );
  AND U7095 ( .A(p_input[7873]), .B(p_input[37873]), .Z(n4729) );
  AND U7096 ( .A(n4731), .B(n4732), .Z(o[7872]) );
  AND U7097 ( .A(p_input[27872]), .B(p_input[17872]), .Z(n4732) );
  AND U7098 ( .A(p_input[7872]), .B(p_input[37872]), .Z(n4731) );
  AND U7099 ( .A(n4733), .B(n4734), .Z(o[7871]) );
  AND U7100 ( .A(p_input[27871]), .B(p_input[17871]), .Z(n4734) );
  AND U7101 ( .A(p_input[7871]), .B(p_input[37871]), .Z(n4733) );
  AND U7102 ( .A(n4735), .B(n4736), .Z(o[7870]) );
  AND U7103 ( .A(p_input[27870]), .B(p_input[17870]), .Z(n4736) );
  AND U7104 ( .A(p_input[7870]), .B(p_input[37870]), .Z(n4735) );
  AND U7105 ( .A(n4737), .B(n4738), .Z(o[786]) );
  AND U7106 ( .A(p_input[20786]), .B(p_input[10786]), .Z(n4738) );
  AND U7107 ( .A(p_input[786]), .B(p_input[30786]), .Z(n4737) );
  AND U7108 ( .A(n4739), .B(n4740), .Z(o[7869]) );
  AND U7109 ( .A(p_input[27869]), .B(p_input[17869]), .Z(n4740) );
  AND U7110 ( .A(p_input[7869]), .B(p_input[37869]), .Z(n4739) );
  AND U7111 ( .A(n4741), .B(n4742), .Z(o[7868]) );
  AND U7112 ( .A(p_input[27868]), .B(p_input[17868]), .Z(n4742) );
  AND U7113 ( .A(p_input[7868]), .B(p_input[37868]), .Z(n4741) );
  AND U7114 ( .A(n4743), .B(n4744), .Z(o[7867]) );
  AND U7115 ( .A(p_input[27867]), .B(p_input[17867]), .Z(n4744) );
  AND U7116 ( .A(p_input[7867]), .B(p_input[37867]), .Z(n4743) );
  AND U7117 ( .A(n4745), .B(n4746), .Z(o[7866]) );
  AND U7118 ( .A(p_input[27866]), .B(p_input[17866]), .Z(n4746) );
  AND U7119 ( .A(p_input[7866]), .B(p_input[37866]), .Z(n4745) );
  AND U7120 ( .A(n4747), .B(n4748), .Z(o[7865]) );
  AND U7121 ( .A(p_input[27865]), .B(p_input[17865]), .Z(n4748) );
  AND U7122 ( .A(p_input[7865]), .B(p_input[37865]), .Z(n4747) );
  AND U7123 ( .A(n4749), .B(n4750), .Z(o[7864]) );
  AND U7124 ( .A(p_input[27864]), .B(p_input[17864]), .Z(n4750) );
  AND U7125 ( .A(p_input[7864]), .B(p_input[37864]), .Z(n4749) );
  AND U7126 ( .A(n4751), .B(n4752), .Z(o[7863]) );
  AND U7127 ( .A(p_input[27863]), .B(p_input[17863]), .Z(n4752) );
  AND U7128 ( .A(p_input[7863]), .B(p_input[37863]), .Z(n4751) );
  AND U7129 ( .A(n4753), .B(n4754), .Z(o[7862]) );
  AND U7130 ( .A(p_input[27862]), .B(p_input[17862]), .Z(n4754) );
  AND U7131 ( .A(p_input[7862]), .B(p_input[37862]), .Z(n4753) );
  AND U7132 ( .A(n4755), .B(n4756), .Z(o[7861]) );
  AND U7133 ( .A(p_input[27861]), .B(p_input[17861]), .Z(n4756) );
  AND U7134 ( .A(p_input[7861]), .B(p_input[37861]), .Z(n4755) );
  AND U7135 ( .A(n4757), .B(n4758), .Z(o[7860]) );
  AND U7136 ( .A(p_input[27860]), .B(p_input[17860]), .Z(n4758) );
  AND U7137 ( .A(p_input[7860]), .B(p_input[37860]), .Z(n4757) );
  AND U7138 ( .A(n4759), .B(n4760), .Z(o[785]) );
  AND U7139 ( .A(p_input[20785]), .B(p_input[10785]), .Z(n4760) );
  AND U7140 ( .A(p_input[785]), .B(p_input[30785]), .Z(n4759) );
  AND U7141 ( .A(n4761), .B(n4762), .Z(o[7859]) );
  AND U7142 ( .A(p_input[27859]), .B(p_input[17859]), .Z(n4762) );
  AND U7143 ( .A(p_input[7859]), .B(p_input[37859]), .Z(n4761) );
  AND U7144 ( .A(n4763), .B(n4764), .Z(o[7858]) );
  AND U7145 ( .A(p_input[27858]), .B(p_input[17858]), .Z(n4764) );
  AND U7146 ( .A(p_input[7858]), .B(p_input[37858]), .Z(n4763) );
  AND U7147 ( .A(n4765), .B(n4766), .Z(o[7857]) );
  AND U7148 ( .A(p_input[27857]), .B(p_input[17857]), .Z(n4766) );
  AND U7149 ( .A(p_input[7857]), .B(p_input[37857]), .Z(n4765) );
  AND U7150 ( .A(n4767), .B(n4768), .Z(o[7856]) );
  AND U7151 ( .A(p_input[27856]), .B(p_input[17856]), .Z(n4768) );
  AND U7152 ( .A(p_input[7856]), .B(p_input[37856]), .Z(n4767) );
  AND U7153 ( .A(n4769), .B(n4770), .Z(o[7855]) );
  AND U7154 ( .A(p_input[27855]), .B(p_input[17855]), .Z(n4770) );
  AND U7155 ( .A(p_input[7855]), .B(p_input[37855]), .Z(n4769) );
  AND U7156 ( .A(n4771), .B(n4772), .Z(o[7854]) );
  AND U7157 ( .A(p_input[27854]), .B(p_input[17854]), .Z(n4772) );
  AND U7158 ( .A(p_input[7854]), .B(p_input[37854]), .Z(n4771) );
  AND U7159 ( .A(n4773), .B(n4774), .Z(o[7853]) );
  AND U7160 ( .A(p_input[27853]), .B(p_input[17853]), .Z(n4774) );
  AND U7161 ( .A(p_input[7853]), .B(p_input[37853]), .Z(n4773) );
  AND U7162 ( .A(n4775), .B(n4776), .Z(o[7852]) );
  AND U7163 ( .A(p_input[27852]), .B(p_input[17852]), .Z(n4776) );
  AND U7164 ( .A(p_input[7852]), .B(p_input[37852]), .Z(n4775) );
  AND U7165 ( .A(n4777), .B(n4778), .Z(o[7851]) );
  AND U7166 ( .A(p_input[27851]), .B(p_input[17851]), .Z(n4778) );
  AND U7167 ( .A(p_input[7851]), .B(p_input[37851]), .Z(n4777) );
  AND U7168 ( .A(n4779), .B(n4780), .Z(o[7850]) );
  AND U7169 ( .A(p_input[27850]), .B(p_input[17850]), .Z(n4780) );
  AND U7170 ( .A(p_input[7850]), .B(p_input[37850]), .Z(n4779) );
  AND U7171 ( .A(n4781), .B(n4782), .Z(o[784]) );
  AND U7172 ( .A(p_input[20784]), .B(p_input[10784]), .Z(n4782) );
  AND U7173 ( .A(p_input[784]), .B(p_input[30784]), .Z(n4781) );
  AND U7174 ( .A(n4783), .B(n4784), .Z(o[7849]) );
  AND U7175 ( .A(p_input[27849]), .B(p_input[17849]), .Z(n4784) );
  AND U7176 ( .A(p_input[7849]), .B(p_input[37849]), .Z(n4783) );
  AND U7177 ( .A(n4785), .B(n4786), .Z(o[7848]) );
  AND U7178 ( .A(p_input[27848]), .B(p_input[17848]), .Z(n4786) );
  AND U7179 ( .A(p_input[7848]), .B(p_input[37848]), .Z(n4785) );
  AND U7180 ( .A(n4787), .B(n4788), .Z(o[7847]) );
  AND U7181 ( .A(p_input[27847]), .B(p_input[17847]), .Z(n4788) );
  AND U7182 ( .A(p_input[7847]), .B(p_input[37847]), .Z(n4787) );
  AND U7183 ( .A(n4789), .B(n4790), .Z(o[7846]) );
  AND U7184 ( .A(p_input[27846]), .B(p_input[17846]), .Z(n4790) );
  AND U7185 ( .A(p_input[7846]), .B(p_input[37846]), .Z(n4789) );
  AND U7186 ( .A(n4791), .B(n4792), .Z(o[7845]) );
  AND U7187 ( .A(p_input[27845]), .B(p_input[17845]), .Z(n4792) );
  AND U7188 ( .A(p_input[7845]), .B(p_input[37845]), .Z(n4791) );
  AND U7189 ( .A(n4793), .B(n4794), .Z(o[7844]) );
  AND U7190 ( .A(p_input[27844]), .B(p_input[17844]), .Z(n4794) );
  AND U7191 ( .A(p_input[7844]), .B(p_input[37844]), .Z(n4793) );
  AND U7192 ( .A(n4795), .B(n4796), .Z(o[7843]) );
  AND U7193 ( .A(p_input[27843]), .B(p_input[17843]), .Z(n4796) );
  AND U7194 ( .A(p_input[7843]), .B(p_input[37843]), .Z(n4795) );
  AND U7195 ( .A(n4797), .B(n4798), .Z(o[7842]) );
  AND U7196 ( .A(p_input[27842]), .B(p_input[17842]), .Z(n4798) );
  AND U7197 ( .A(p_input[7842]), .B(p_input[37842]), .Z(n4797) );
  AND U7198 ( .A(n4799), .B(n4800), .Z(o[7841]) );
  AND U7199 ( .A(p_input[27841]), .B(p_input[17841]), .Z(n4800) );
  AND U7200 ( .A(p_input[7841]), .B(p_input[37841]), .Z(n4799) );
  AND U7201 ( .A(n4801), .B(n4802), .Z(o[7840]) );
  AND U7202 ( .A(p_input[27840]), .B(p_input[17840]), .Z(n4802) );
  AND U7203 ( .A(p_input[7840]), .B(p_input[37840]), .Z(n4801) );
  AND U7204 ( .A(n4803), .B(n4804), .Z(o[783]) );
  AND U7205 ( .A(p_input[20783]), .B(p_input[10783]), .Z(n4804) );
  AND U7206 ( .A(p_input[783]), .B(p_input[30783]), .Z(n4803) );
  AND U7207 ( .A(n4805), .B(n4806), .Z(o[7839]) );
  AND U7208 ( .A(p_input[27839]), .B(p_input[17839]), .Z(n4806) );
  AND U7209 ( .A(p_input[7839]), .B(p_input[37839]), .Z(n4805) );
  AND U7210 ( .A(n4807), .B(n4808), .Z(o[7838]) );
  AND U7211 ( .A(p_input[27838]), .B(p_input[17838]), .Z(n4808) );
  AND U7212 ( .A(p_input[7838]), .B(p_input[37838]), .Z(n4807) );
  AND U7213 ( .A(n4809), .B(n4810), .Z(o[7837]) );
  AND U7214 ( .A(p_input[27837]), .B(p_input[17837]), .Z(n4810) );
  AND U7215 ( .A(p_input[7837]), .B(p_input[37837]), .Z(n4809) );
  AND U7216 ( .A(n4811), .B(n4812), .Z(o[7836]) );
  AND U7217 ( .A(p_input[27836]), .B(p_input[17836]), .Z(n4812) );
  AND U7218 ( .A(p_input[7836]), .B(p_input[37836]), .Z(n4811) );
  AND U7219 ( .A(n4813), .B(n4814), .Z(o[7835]) );
  AND U7220 ( .A(p_input[27835]), .B(p_input[17835]), .Z(n4814) );
  AND U7221 ( .A(p_input[7835]), .B(p_input[37835]), .Z(n4813) );
  AND U7222 ( .A(n4815), .B(n4816), .Z(o[7834]) );
  AND U7223 ( .A(p_input[27834]), .B(p_input[17834]), .Z(n4816) );
  AND U7224 ( .A(p_input[7834]), .B(p_input[37834]), .Z(n4815) );
  AND U7225 ( .A(n4817), .B(n4818), .Z(o[7833]) );
  AND U7226 ( .A(p_input[27833]), .B(p_input[17833]), .Z(n4818) );
  AND U7227 ( .A(p_input[7833]), .B(p_input[37833]), .Z(n4817) );
  AND U7228 ( .A(n4819), .B(n4820), .Z(o[7832]) );
  AND U7229 ( .A(p_input[27832]), .B(p_input[17832]), .Z(n4820) );
  AND U7230 ( .A(p_input[7832]), .B(p_input[37832]), .Z(n4819) );
  AND U7231 ( .A(n4821), .B(n4822), .Z(o[7831]) );
  AND U7232 ( .A(p_input[27831]), .B(p_input[17831]), .Z(n4822) );
  AND U7233 ( .A(p_input[7831]), .B(p_input[37831]), .Z(n4821) );
  AND U7234 ( .A(n4823), .B(n4824), .Z(o[7830]) );
  AND U7235 ( .A(p_input[27830]), .B(p_input[17830]), .Z(n4824) );
  AND U7236 ( .A(p_input[7830]), .B(p_input[37830]), .Z(n4823) );
  AND U7237 ( .A(n4825), .B(n4826), .Z(o[782]) );
  AND U7238 ( .A(p_input[20782]), .B(p_input[10782]), .Z(n4826) );
  AND U7239 ( .A(p_input[782]), .B(p_input[30782]), .Z(n4825) );
  AND U7240 ( .A(n4827), .B(n4828), .Z(o[7829]) );
  AND U7241 ( .A(p_input[27829]), .B(p_input[17829]), .Z(n4828) );
  AND U7242 ( .A(p_input[7829]), .B(p_input[37829]), .Z(n4827) );
  AND U7243 ( .A(n4829), .B(n4830), .Z(o[7828]) );
  AND U7244 ( .A(p_input[27828]), .B(p_input[17828]), .Z(n4830) );
  AND U7245 ( .A(p_input[7828]), .B(p_input[37828]), .Z(n4829) );
  AND U7246 ( .A(n4831), .B(n4832), .Z(o[7827]) );
  AND U7247 ( .A(p_input[27827]), .B(p_input[17827]), .Z(n4832) );
  AND U7248 ( .A(p_input[7827]), .B(p_input[37827]), .Z(n4831) );
  AND U7249 ( .A(n4833), .B(n4834), .Z(o[7826]) );
  AND U7250 ( .A(p_input[27826]), .B(p_input[17826]), .Z(n4834) );
  AND U7251 ( .A(p_input[7826]), .B(p_input[37826]), .Z(n4833) );
  AND U7252 ( .A(n4835), .B(n4836), .Z(o[7825]) );
  AND U7253 ( .A(p_input[27825]), .B(p_input[17825]), .Z(n4836) );
  AND U7254 ( .A(p_input[7825]), .B(p_input[37825]), .Z(n4835) );
  AND U7255 ( .A(n4837), .B(n4838), .Z(o[7824]) );
  AND U7256 ( .A(p_input[27824]), .B(p_input[17824]), .Z(n4838) );
  AND U7257 ( .A(p_input[7824]), .B(p_input[37824]), .Z(n4837) );
  AND U7258 ( .A(n4839), .B(n4840), .Z(o[7823]) );
  AND U7259 ( .A(p_input[27823]), .B(p_input[17823]), .Z(n4840) );
  AND U7260 ( .A(p_input[7823]), .B(p_input[37823]), .Z(n4839) );
  AND U7261 ( .A(n4841), .B(n4842), .Z(o[7822]) );
  AND U7262 ( .A(p_input[27822]), .B(p_input[17822]), .Z(n4842) );
  AND U7263 ( .A(p_input[7822]), .B(p_input[37822]), .Z(n4841) );
  AND U7264 ( .A(n4843), .B(n4844), .Z(o[7821]) );
  AND U7265 ( .A(p_input[27821]), .B(p_input[17821]), .Z(n4844) );
  AND U7266 ( .A(p_input[7821]), .B(p_input[37821]), .Z(n4843) );
  AND U7267 ( .A(n4845), .B(n4846), .Z(o[7820]) );
  AND U7268 ( .A(p_input[27820]), .B(p_input[17820]), .Z(n4846) );
  AND U7269 ( .A(p_input[7820]), .B(p_input[37820]), .Z(n4845) );
  AND U7270 ( .A(n4847), .B(n4848), .Z(o[781]) );
  AND U7271 ( .A(p_input[20781]), .B(p_input[10781]), .Z(n4848) );
  AND U7272 ( .A(p_input[781]), .B(p_input[30781]), .Z(n4847) );
  AND U7273 ( .A(n4849), .B(n4850), .Z(o[7819]) );
  AND U7274 ( .A(p_input[27819]), .B(p_input[17819]), .Z(n4850) );
  AND U7275 ( .A(p_input[7819]), .B(p_input[37819]), .Z(n4849) );
  AND U7276 ( .A(n4851), .B(n4852), .Z(o[7818]) );
  AND U7277 ( .A(p_input[27818]), .B(p_input[17818]), .Z(n4852) );
  AND U7278 ( .A(p_input[7818]), .B(p_input[37818]), .Z(n4851) );
  AND U7279 ( .A(n4853), .B(n4854), .Z(o[7817]) );
  AND U7280 ( .A(p_input[27817]), .B(p_input[17817]), .Z(n4854) );
  AND U7281 ( .A(p_input[7817]), .B(p_input[37817]), .Z(n4853) );
  AND U7282 ( .A(n4855), .B(n4856), .Z(o[7816]) );
  AND U7283 ( .A(p_input[27816]), .B(p_input[17816]), .Z(n4856) );
  AND U7284 ( .A(p_input[7816]), .B(p_input[37816]), .Z(n4855) );
  AND U7285 ( .A(n4857), .B(n4858), .Z(o[7815]) );
  AND U7286 ( .A(p_input[27815]), .B(p_input[17815]), .Z(n4858) );
  AND U7287 ( .A(p_input[7815]), .B(p_input[37815]), .Z(n4857) );
  AND U7288 ( .A(n4859), .B(n4860), .Z(o[7814]) );
  AND U7289 ( .A(p_input[27814]), .B(p_input[17814]), .Z(n4860) );
  AND U7290 ( .A(p_input[7814]), .B(p_input[37814]), .Z(n4859) );
  AND U7291 ( .A(n4861), .B(n4862), .Z(o[7813]) );
  AND U7292 ( .A(p_input[27813]), .B(p_input[17813]), .Z(n4862) );
  AND U7293 ( .A(p_input[7813]), .B(p_input[37813]), .Z(n4861) );
  AND U7294 ( .A(n4863), .B(n4864), .Z(o[7812]) );
  AND U7295 ( .A(p_input[27812]), .B(p_input[17812]), .Z(n4864) );
  AND U7296 ( .A(p_input[7812]), .B(p_input[37812]), .Z(n4863) );
  AND U7297 ( .A(n4865), .B(n4866), .Z(o[7811]) );
  AND U7298 ( .A(p_input[27811]), .B(p_input[17811]), .Z(n4866) );
  AND U7299 ( .A(p_input[7811]), .B(p_input[37811]), .Z(n4865) );
  AND U7300 ( .A(n4867), .B(n4868), .Z(o[7810]) );
  AND U7301 ( .A(p_input[27810]), .B(p_input[17810]), .Z(n4868) );
  AND U7302 ( .A(p_input[7810]), .B(p_input[37810]), .Z(n4867) );
  AND U7303 ( .A(n4869), .B(n4870), .Z(o[780]) );
  AND U7304 ( .A(p_input[20780]), .B(p_input[10780]), .Z(n4870) );
  AND U7305 ( .A(p_input[780]), .B(p_input[30780]), .Z(n4869) );
  AND U7306 ( .A(n4871), .B(n4872), .Z(o[7809]) );
  AND U7307 ( .A(p_input[27809]), .B(p_input[17809]), .Z(n4872) );
  AND U7308 ( .A(p_input[7809]), .B(p_input[37809]), .Z(n4871) );
  AND U7309 ( .A(n4873), .B(n4874), .Z(o[7808]) );
  AND U7310 ( .A(p_input[27808]), .B(p_input[17808]), .Z(n4874) );
  AND U7311 ( .A(p_input[7808]), .B(p_input[37808]), .Z(n4873) );
  AND U7312 ( .A(n4875), .B(n4876), .Z(o[7807]) );
  AND U7313 ( .A(p_input[27807]), .B(p_input[17807]), .Z(n4876) );
  AND U7314 ( .A(p_input[7807]), .B(p_input[37807]), .Z(n4875) );
  AND U7315 ( .A(n4877), .B(n4878), .Z(o[7806]) );
  AND U7316 ( .A(p_input[27806]), .B(p_input[17806]), .Z(n4878) );
  AND U7317 ( .A(p_input[7806]), .B(p_input[37806]), .Z(n4877) );
  AND U7318 ( .A(n4879), .B(n4880), .Z(o[7805]) );
  AND U7319 ( .A(p_input[27805]), .B(p_input[17805]), .Z(n4880) );
  AND U7320 ( .A(p_input[7805]), .B(p_input[37805]), .Z(n4879) );
  AND U7321 ( .A(n4881), .B(n4882), .Z(o[7804]) );
  AND U7322 ( .A(p_input[27804]), .B(p_input[17804]), .Z(n4882) );
  AND U7323 ( .A(p_input[7804]), .B(p_input[37804]), .Z(n4881) );
  AND U7324 ( .A(n4883), .B(n4884), .Z(o[7803]) );
  AND U7325 ( .A(p_input[27803]), .B(p_input[17803]), .Z(n4884) );
  AND U7326 ( .A(p_input[7803]), .B(p_input[37803]), .Z(n4883) );
  AND U7327 ( .A(n4885), .B(n4886), .Z(o[7802]) );
  AND U7328 ( .A(p_input[27802]), .B(p_input[17802]), .Z(n4886) );
  AND U7329 ( .A(p_input[7802]), .B(p_input[37802]), .Z(n4885) );
  AND U7330 ( .A(n4887), .B(n4888), .Z(o[7801]) );
  AND U7331 ( .A(p_input[27801]), .B(p_input[17801]), .Z(n4888) );
  AND U7332 ( .A(p_input[7801]), .B(p_input[37801]), .Z(n4887) );
  AND U7333 ( .A(n4889), .B(n4890), .Z(o[7800]) );
  AND U7334 ( .A(p_input[27800]), .B(p_input[17800]), .Z(n4890) );
  AND U7335 ( .A(p_input[7800]), .B(p_input[37800]), .Z(n4889) );
  AND U7336 ( .A(n4891), .B(n4892), .Z(o[77]) );
  AND U7337 ( .A(p_input[20077]), .B(p_input[10077]), .Z(n4892) );
  AND U7338 ( .A(p_input[77]), .B(p_input[30077]), .Z(n4891) );
  AND U7339 ( .A(n4893), .B(n4894), .Z(o[779]) );
  AND U7340 ( .A(p_input[20779]), .B(p_input[10779]), .Z(n4894) );
  AND U7341 ( .A(p_input[779]), .B(p_input[30779]), .Z(n4893) );
  AND U7342 ( .A(n4895), .B(n4896), .Z(o[7799]) );
  AND U7343 ( .A(p_input[27799]), .B(p_input[17799]), .Z(n4896) );
  AND U7344 ( .A(p_input[7799]), .B(p_input[37799]), .Z(n4895) );
  AND U7345 ( .A(n4897), .B(n4898), .Z(o[7798]) );
  AND U7346 ( .A(p_input[27798]), .B(p_input[17798]), .Z(n4898) );
  AND U7347 ( .A(p_input[7798]), .B(p_input[37798]), .Z(n4897) );
  AND U7348 ( .A(n4899), .B(n4900), .Z(o[7797]) );
  AND U7349 ( .A(p_input[27797]), .B(p_input[17797]), .Z(n4900) );
  AND U7350 ( .A(p_input[7797]), .B(p_input[37797]), .Z(n4899) );
  AND U7351 ( .A(n4901), .B(n4902), .Z(o[7796]) );
  AND U7352 ( .A(p_input[27796]), .B(p_input[17796]), .Z(n4902) );
  AND U7353 ( .A(p_input[7796]), .B(p_input[37796]), .Z(n4901) );
  AND U7354 ( .A(n4903), .B(n4904), .Z(o[7795]) );
  AND U7355 ( .A(p_input[27795]), .B(p_input[17795]), .Z(n4904) );
  AND U7356 ( .A(p_input[7795]), .B(p_input[37795]), .Z(n4903) );
  AND U7357 ( .A(n4905), .B(n4906), .Z(o[7794]) );
  AND U7358 ( .A(p_input[27794]), .B(p_input[17794]), .Z(n4906) );
  AND U7359 ( .A(p_input[7794]), .B(p_input[37794]), .Z(n4905) );
  AND U7360 ( .A(n4907), .B(n4908), .Z(o[7793]) );
  AND U7361 ( .A(p_input[27793]), .B(p_input[17793]), .Z(n4908) );
  AND U7362 ( .A(p_input[7793]), .B(p_input[37793]), .Z(n4907) );
  AND U7363 ( .A(n4909), .B(n4910), .Z(o[7792]) );
  AND U7364 ( .A(p_input[27792]), .B(p_input[17792]), .Z(n4910) );
  AND U7365 ( .A(p_input[7792]), .B(p_input[37792]), .Z(n4909) );
  AND U7366 ( .A(n4911), .B(n4912), .Z(o[7791]) );
  AND U7367 ( .A(p_input[27791]), .B(p_input[17791]), .Z(n4912) );
  AND U7368 ( .A(p_input[7791]), .B(p_input[37791]), .Z(n4911) );
  AND U7369 ( .A(n4913), .B(n4914), .Z(o[7790]) );
  AND U7370 ( .A(p_input[27790]), .B(p_input[17790]), .Z(n4914) );
  AND U7371 ( .A(p_input[7790]), .B(p_input[37790]), .Z(n4913) );
  AND U7372 ( .A(n4915), .B(n4916), .Z(o[778]) );
  AND U7373 ( .A(p_input[20778]), .B(p_input[10778]), .Z(n4916) );
  AND U7374 ( .A(p_input[778]), .B(p_input[30778]), .Z(n4915) );
  AND U7375 ( .A(n4917), .B(n4918), .Z(o[7789]) );
  AND U7376 ( .A(p_input[27789]), .B(p_input[17789]), .Z(n4918) );
  AND U7377 ( .A(p_input[7789]), .B(p_input[37789]), .Z(n4917) );
  AND U7378 ( .A(n4919), .B(n4920), .Z(o[7788]) );
  AND U7379 ( .A(p_input[27788]), .B(p_input[17788]), .Z(n4920) );
  AND U7380 ( .A(p_input[7788]), .B(p_input[37788]), .Z(n4919) );
  AND U7381 ( .A(n4921), .B(n4922), .Z(o[7787]) );
  AND U7382 ( .A(p_input[27787]), .B(p_input[17787]), .Z(n4922) );
  AND U7383 ( .A(p_input[7787]), .B(p_input[37787]), .Z(n4921) );
  AND U7384 ( .A(n4923), .B(n4924), .Z(o[7786]) );
  AND U7385 ( .A(p_input[27786]), .B(p_input[17786]), .Z(n4924) );
  AND U7386 ( .A(p_input[7786]), .B(p_input[37786]), .Z(n4923) );
  AND U7387 ( .A(n4925), .B(n4926), .Z(o[7785]) );
  AND U7388 ( .A(p_input[27785]), .B(p_input[17785]), .Z(n4926) );
  AND U7389 ( .A(p_input[7785]), .B(p_input[37785]), .Z(n4925) );
  AND U7390 ( .A(n4927), .B(n4928), .Z(o[7784]) );
  AND U7391 ( .A(p_input[27784]), .B(p_input[17784]), .Z(n4928) );
  AND U7392 ( .A(p_input[7784]), .B(p_input[37784]), .Z(n4927) );
  AND U7393 ( .A(n4929), .B(n4930), .Z(o[7783]) );
  AND U7394 ( .A(p_input[27783]), .B(p_input[17783]), .Z(n4930) );
  AND U7395 ( .A(p_input[7783]), .B(p_input[37783]), .Z(n4929) );
  AND U7396 ( .A(n4931), .B(n4932), .Z(o[7782]) );
  AND U7397 ( .A(p_input[27782]), .B(p_input[17782]), .Z(n4932) );
  AND U7398 ( .A(p_input[7782]), .B(p_input[37782]), .Z(n4931) );
  AND U7399 ( .A(n4933), .B(n4934), .Z(o[7781]) );
  AND U7400 ( .A(p_input[27781]), .B(p_input[17781]), .Z(n4934) );
  AND U7401 ( .A(p_input[7781]), .B(p_input[37781]), .Z(n4933) );
  AND U7402 ( .A(n4935), .B(n4936), .Z(o[7780]) );
  AND U7403 ( .A(p_input[27780]), .B(p_input[17780]), .Z(n4936) );
  AND U7404 ( .A(p_input[7780]), .B(p_input[37780]), .Z(n4935) );
  AND U7405 ( .A(n4937), .B(n4938), .Z(o[777]) );
  AND U7406 ( .A(p_input[20777]), .B(p_input[10777]), .Z(n4938) );
  AND U7407 ( .A(p_input[777]), .B(p_input[30777]), .Z(n4937) );
  AND U7408 ( .A(n4939), .B(n4940), .Z(o[7779]) );
  AND U7409 ( .A(p_input[27779]), .B(p_input[17779]), .Z(n4940) );
  AND U7410 ( .A(p_input[7779]), .B(p_input[37779]), .Z(n4939) );
  AND U7411 ( .A(n4941), .B(n4942), .Z(o[7778]) );
  AND U7412 ( .A(p_input[27778]), .B(p_input[17778]), .Z(n4942) );
  AND U7413 ( .A(p_input[7778]), .B(p_input[37778]), .Z(n4941) );
  AND U7414 ( .A(n4943), .B(n4944), .Z(o[7777]) );
  AND U7415 ( .A(p_input[27777]), .B(p_input[17777]), .Z(n4944) );
  AND U7416 ( .A(p_input[7777]), .B(p_input[37777]), .Z(n4943) );
  AND U7417 ( .A(n4945), .B(n4946), .Z(o[7776]) );
  AND U7418 ( .A(p_input[27776]), .B(p_input[17776]), .Z(n4946) );
  AND U7419 ( .A(p_input[7776]), .B(p_input[37776]), .Z(n4945) );
  AND U7420 ( .A(n4947), .B(n4948), .Z(o[7775]) );
  AND U7421 ( .A(p_input[27775]), .B(p_input[17775]), .Z(n4948) );
  AND U7422 ( .A(p_input[7775]), .B(p_input[37775]), .Z(n4947) );
  AND U7423 ( .A(n4949), .B(n4950), .Z(o[7774]) );
  AND U7424 ( .A(p_input[27774]), .B(p_input[17774]), .Z(n4950) );
  AND U7425 ( .A(p_input[7774]), .B(p_input[37774]), .Z(n4949) );
  AND U7426 ( .A(n4951), .B(n4952), .Z(o[7773]) );
  AND U7427 ( .A(p_input[27773]), .B(p_input[17773]), .Z(n4952) );
  AND U7428 ( .A(p_input[7773]), .B(p_input[37773]), .Z(n4951) );
  AND U7429 ( .A(n4953), .B(n4954), .Z(o[7772]) );
  AND U7430 ( .A(p_input[27772]), .B(p_input[17772]), .Z(n4954) );
  AND U7431 ( .A(p_input[7772]), .B(p_input[37772]), .Z(n4953) );
  AND U7432 ( .A(n4955), .B(n4956), .Z(o[7771]) );
  AND U7433 ( .A(p_input[27771]), .B(p_input[17771]), .Z(n4956) );
  AND U7434 ( .A(p_input[7771]), .B(p_input[37771]), .Z(n4955) );
  AND U7435 ( .A(n4957), .B(n4958), .Z(o[7770]) );
  AND U7436 ( .A(p_input[27770]), .B(p_input[17770]), .Z(n4958) );
  AND U7437 ( .A(p_input[7770]), .B(p_input[37770]), .Z(n4957) );
  AND U7438 ( .A(n4959), .B(n4960), .Z(o[776]) );
  AND U7439 ( .A(p_input[20776]), .B(p_input[10776]), .Z(n4960) );
  AND U7440 ( .A(p_input[776]), .B(p_input[30776]), .Z(n4959) );
  AND U7441 ( .A(n4961), .B(n4962), .Z(o[7769]) );
  AND U7442 ( .A(p_input[27769]), .B(p_input[17769]), .Z(n4962) );
  AND U7443 ( .A(p_input[7769]), .B(p_input[37769]), .Z(n4961) );
  AND U7444 ( .A(n4963), .B(n4964), .Z(o[7768]) );
  AND U7445 ( .A(p_input[27768]), .B(p_input[17768]), .Z(n4964) );
  AND U7446 ( .A(p_input[7768]), .B(p_input[37768]), .Z(n4963) );
  AND U7447 ( .A(n4965), .B(n4966), .Z(o[7767]) );
  AND U7448 ( .A(p_input[27767]), .B(p_input[17767]), .Z(n4966) );
  AND U7449 ( .A(p_input[7767]), .B(p_input[37767]), .Z(n4965) );
  AND U7450 ( .A(n4967), .B(n4968), .Z(o[7766]) );
  AND U7451 ( .A(p_input[27766]), .B(p_input[17766]), .Z(n4968) );
  AND U7452 ( .A(p_input[7766]), .B(p_input[37766]), .Z(n4967) );
  AND U7453 ( .A(n4969), .B(n4970), .Z(o[7765]) );
  AND U7454 ( .A(p_input[27765]), .B(p_input[17765]), .Z(n4970) );
  AND U7455 ( .A(p_input[7765]), .B(p_input[37765]), .Z(n4969) );
  AND U7456 ( .A(n4971), .B(n4972), .Z(o[7764]) );
  AND U7457 ( .A(p_input[27764]), .B(p_input[17764]), .Z(n4972) );
  AND U7458 ( .A(p_input[7764]), .B(p_input[37764]), .Z(n4971) );
  AND U7459 ( .A(n4973), .B(n4974), .Z(o[7763]) );
  AND U7460 ( .A(p_input[27763]), .B(p_input[17763]), .Z(n4974) );
  AND U7461 ( .A(p_input[7763]), .B(p_input[37763]), .Z(n4973) );
  AND U7462 ( .A(n4975), .B(n4976), .Z(o[7762]) );
  AND U7463 ( .A(p_input[27762]), .B(p_input[17762]), .Z(n4976) );
  AND U7464 ( .A(p_input[7762]), .B(p_input[37762]), .Z(n4975) );
  AND U7465 ( .A(n4977), .B(n4978), .Z(o[7761]) );
  AND U7466 ( .A(p_input[27761]), .B(p_input[17761]), .Z(n4978) );
  AND U7467 ( .A(p_input[7761]), .B(p_input[37761]), .Z(n4977) );
  AND U7468 ( .A(n4979), .B(n4980), .Z(o[7760]) );
  AND U7469 ( .A(p_input[27760]), .B(p_input[17760]), .Z(n4980) );
  AND U7470 ( .A(p_input[7760]), .B(p_input[37760]), .Z(n4979) );
  AND U7471 ( .A(n4981), .B(n4982), .Z(o[775]) );
  AND U7472 ( .A(p_input[20775]), .B(p_input[10775]), .Z(n4982) );
  AND U7473 ( .A(p_input[775]), .B(p_input[30775]), .Z(n4981) );
  AND U7474 ( .A(n4983), .B(n4984), .Z(o[7759]) );
  AND U7475 ( .A(p_input[27759]), .B(p_input[17759]), .Z(n4984) );
  AND U7476 ( .A(p_input[7759]), .B(p_input[37759]), .Z(n4983) );
  AND U7477 ( .A(n4985), .B(n4986), .Z(o[7758]) );
  AND U7478 ( .A(p_input[27758]), .B(p_input[17758]), .Z(n4986) );
  AND U7479 ( .A(p_input[7758]), .B(p_input[37758]), .Z(n4985) );
  AND U7480 ( .A(n4987), .B(n4988), .Z(o[7757]) );
  AND U7481 ( .A(p_input[27757]), .B(p_input[17757]), .Z(n4988) );
  AND U7482 ( .A(p_input[7757]), .B(p_input[37757]), .Z(n4987) );
  AND U7483 ( .A(n4989), .B(n4990), .Z(o[7756]) );
  AND U7484 ( .A(p_input[27756]), .B(p_input[17756]), .Z(n4990) );
  AND U7485 ( .A(p_input[7756]), .B(p_input[37756]), .Z(n4989) );
  AND U7486 ( .A(n4991), .B(n4992), .Z(o[7755]) );
  AND U7487 ( .A(p_input[27755]), .B(p_input[17755]), .Z(n4992) );
  AND U7488 ( .A(p_input[7755]), .B(p_input[37755]), .Z(n4991) );
  AND U7489 ( .A(n4993), .B(n4994), .Z(o[7754]) );
  AND U7490 ( .A(p_input[27754]), .B(p_input[17754]), .Z(n4994) );
  AND U7491 ( .A(p_input[7754]), .B(p_input[37754]), .Z(n4993) );
  AND U7492 ( .A(n4995), .B(n4996), .Z(o[7753]) );
  AND U7493 ( .A(p_input[27753]), .B(p_input[17753]), .Z(n4996) );
  AND U7494 ( .A(p_input[7753]), .B(p_input[37753]), .Z(n4995) );
  AND U7495 ( .A(n4997), .B(n4998), .Z(o[7752]) );
  AND U7496 ( .A(p_input[27752]), .B(p_input[17752]), .Z(n4998) );
  AND U7497 ( .A(p_input[7752]), .B(p_input[37752]), .Z(n4997) );
  AND U7498 ( .A(n4999), .B(n5000), .Z(o[7751]) );
  AND U7499 ( .A(p_input[27751]), .B(p_input[17751]), .Z(n5000) );
  AND U7500 ( .A(p_input[7751]), .B(p_input[37751]), .Z(n4999) );
  AND U7501 ( .A(n5001), .B(n5002), .Z(o[7750]) );
  AND U7502 ( .A(p_input[27750]), .B(p_input[17750]), .Z(n5002) );
  AND U7503 ( .A(p_input[7750]), .B(p_input[37750]), .Z(n5001) );
  AND U7504 ( .A(n5003), .B(n5004), .Z(o[774]) );
  AND U7505 ( .A(p_input[20774]), .B(p_input[10774]), .Z(n5004) );
  AND U7506 ( .A(p_input[774]), .B(p_input[30774]), .Z(n5003) );
  AND U7507 ( .A(n5005), .B(n5006), .Z(o[7749]) );
  AND U7508 ( .A(p_input[27749]), .B(p_input[17749]), .Z(n5006) );
  AND U7509 ( .A(p_input[7749]), .B(p_input[37749]), .Z(n5005) );
  AND U7510 ( .A(n5007), .B(n5008), .Z(o[7748]) );
  AND U7511 ( .A(p_input[27748]), .B(p_input[17748]), .Z(n5008) );
  AND U7512 ( .A(p_input[7748]), .B(p_input[37748]), .Z(n5007) );
  AND U7513 ( .A(n5009), .B(n5010), .Z(o[7747]) );
  AND U7514 ( .A(p_input[27747]), .B(p_input[17747]), .Z(n5010) );
  AND U7515 ( .A(p_input[7747]), .B(p_input[37747]), .Z(n5009) );
  AND U7516 ( .A(n5011), .B(n5012), .Z(o[7746]) );
  AND U7517 ( .A(p_input[27746]), .B(p_input[17746]), .Z(n5012) );
  AND U7518 ( .A(p_input[7746]), .B(p_input[37746]), .Z(n5011) );
  AND U7519 ( .A(n5013), .B(n5014), .Z(o[7745]) );
  AND U7520 ( .A(p_input[27745]), .B(p_input[17745]), .Z(n5014) );
  AND U7521 ( .A(p_input[7745]), .B(p_input[37745]), .Z(n5013) );
  AND U7522 ( .A(n5015), .B(n5016), .Z(o[7744]) );
  AND U7523 ( .A(p_input[27744]), .B(p_input[17744]), .Z(n5016) );
  AND U7524 ( .A(p_input[7744]), .B(p_input[37744]), .Z(n5015) );
  AND U7525 ( .A(n5017), .B(n5018), .Z(o[7743]) );
  AND U7526 ( .A(p_input[27743]), .B(p_input[17743]), .Z(n5018) );
  AND U7527 ( .A(p_input[7743]), .B(p_input[37743]), .Z(n5017) );
  AND U7528 ( .A(n5019), .B(n5020), .Z(o[7742]) );
  AND U7529 ( .A(p_input[27742]), .B(p_input[17742]), .Z(n5020) );
  AND U7530 ( .A(p_input[7742]), .B(p_input[37742]), .Z(n5019) );
  AND U7531 ( .A(n5021), .B(n5022), .Z(o[7741]) );
  AND U7532 ( .A(p_input[27741]), .B(p_input[17741]), .Z(n5022) );
  AND U7533 ( .A(p_input[7741]), .B(p_input[37741]), .Z(n5021) );
  AND U7534 ( .A(n5023), .B(n5024), .Z(o[7740]) );
  AND U7535 ( .A(p_input[27740]), .B(p_input[17740]), .Z(n5024) );
  AND U7536 ( .A(p_input[7740]), .B(p_input[37740]), .Z(n5023) );
  AND U7537 ( .A(n5025), .B(n5026), .Z(o[773]) );
  AND U7538 ( .A(p_input[20773]), .B(p_input[10773]), .Z(n5026) );
  AND U7539 ( .A(p_input[773]), .B(p_input[30773]), .Z(n5025) );
  AND U7540 ( .A(n5027), .B(n5028), .Z(o[7739]) );
  AND U7541 ( .A(p_input[27739]), .B(p_input[17739]), .Z(n5028) );
  AND U7542 ( .A(p_input[7739]), .B(p_input[37739]), .Z(n5027) );
  AND U7543 ( .A(n5029), .B(n5030), .Z(o[7738]) );
  AND U7544 ( .A(p_input[27738]), .B(p_input[17738]), .Z(n5030) );
  AND U7545 ( .A(p_input[7738]), .B(p_input[37738]), .Z(n5029) );
  AND U7546 ( .A(n5031), .B(n5032), .Z(o[7737]) );
  AND U7547 ( .A(p_input[27737]), .B(p_input[17737]), .Z(n5032) );
  AND U7548 ( .A(p_input[7737]), .B(p_input[37737]), .Z(n5031) );
  AND U7549 ( .A(n5033), .B(n5034), .Z(o[7736]) );
  AND U7550 ( .A(p_input[27736]), .B(p_input[17736]), .Z(n5034) );
  AND U7551 ( .A(p_input[7736]), .B(p_input[37736]), .Z(n5033) );
  AND U7552 ( .A(n5035), .B(n5036), .Z(o[7735]) );
  AND U7553 ( .A(p_input[27735]), .B(p_input[17735]), .Z(n5036) );
  AND U7554 ( .A(p_input[7735]), .B(p_input[37735]), .Z(n5035) );
  AND U7555 ( .A(n5037), .B(n5038), .Z(o[7734]) );
  AND U7556 ( .A(p_input[27734]), .B(p_input[17734]), .Z(n5038) );
  AND U7557 ( .A(p_input[7734]), .B(p_input[37734]), .Z(n5037) );
  AND U7558 ( .A(n5039), .B(n5040), .Z(o[7733]) );
  AND U7559 ( .A(p_input[27733]), .B(p_input[17733]), .Z(n5040) );
  AND U7560 ( .A(p_input[7733]), .B(p_input[37733]), .Z(n5039) );
  AND U7561 ( .A(n5041), .B(n5042), .Z(o[7732]) );
  AND U7562 ( .A(p_input[27732]), .B(p_input[17732]), .Z(n5042) );
  AND U7563 ( .A(p_input[7732]), .B(p_input[37732]), .Z(n5041) );
  AND U7564 ( .A(n5043), .B(n5044), .Z(o[7731]) );
  AND U7565 ( .A(p_input[27731]), .B(p_input[17731]), .Z(n5044) );
  AND U7566 ( .A(p_input[7731]), .B(p_input[37731]), .Z(n5043) );
  AND U7567 ( .A(n5045), .B(n5046), .Z(o[7730]) );
  AND U7568 ( .A(p_input[27730]), .B(p_input[17730]), .Z(n5046) );
  AND U7569 ( .A(p_input[7730]), .B(p_input[37730]), .Z(n5045) );
  AND U7570 ( .A(n5047), .B(n5048), .Z(o[772]) );
  AND U7571 ( .A(p_input[20772]), .B(p_input[10772]), .Z(n5048) );
  AND U7572 ( .A(p_input[772]), .B(p_input[30772]), .Z(n5047) );
  AND U7573 ( .A(n5049), .B(n5050), .Z(o[7729]) );
  AND U7574 ( .A(p_input[27729]), .B(p_input[17729]), .Z(n5050) );
  AND U7575 ( .A(p_input[7729]), .B(p_input[37729]), .Z(n5049) );
  AND U7576 ( .A(n5051), .B(n5052), .Z(o[7728]) );
  AND U7577 ( .A(p_input[27728]), .B(p_input[17728]), .Z(n5052) );
  AND U7578 ( .A(p_input[7728]), .B(p_input[37728]), .Z(n5051) );
  AND U7579 ( .A(n5053), .B(n5054), .Z(o[7727]) );
  AND U7580 ( .A(p_input[27727]), .B(p_input[17727]), .Z(n5054) );
  AND U7581 ( .A(p_input[7727]), .B(p_input[37727]), .Z(n5053) );
  AND U7582 ( .A(n5055), .B(n5056), .Z(o[7726]) );
  AND U7583 ( .A(p_input[27726]), .B(p_input[17726]), .Z(n5056) );
  AND U7584 ( .A(p_input[7726]), .B(p_input[37726]), .Z(n5055) );
  AND U7585 ( .A(n5057), .B(n5058), .Z(o[7725]) );
  AND U7586 ( .A(p_input[27725]), .B(p_input[17725]), .Z(n5058) );
  AND U7587 ( .A(p_input[7725]), .B(p_input[37725]), .Z(n5057) );
  AND U7588 ( .A(n5059), .B(n5060), .Z(o[7724]) );
  AND U7589 ( .A(p_input[27724]), .B(p_input[17724]), .Z(n5060) );
  AND U7590 ( .A(p_input[7724]), .B(p_input[37724]), .Z(n5059) );
  AND U7591 ( .A(n5061), .B(n5062), .Z(o[7723]) );
  AND U7592 ( .A(p_input[27723]), .B(p_input[17723]), .Z(n5062) );
  AND U7593 ( .A(p_input[7723]), .B(p_input[37723]), .Z(n5061) );
  AND U7594 ( .A(n5063), .B(n5064), .Z(o[7722]) );
  AND U7595 ( .A(p_input[27722]), .B(p_input[17722]), .Z(n5064) );
  AND U7596 ( .A(p_input[7722]), .B(p_input[37722]), .Z(n5063) );
  AND U7597 ( .A(n5065), .B(n5066), .Z(o[7721]) );
  AND U7598 ( .A(p_input[27721]), .B(p_input[17721]), .Z(n5066) );
  AND U7599 ( .A(p_input[7721]), .B(p_input[37721]), .Z(n5065) );
  AND U7600 ( .A(n5067), .B(n5068), .Z(o[7720]) );
  AND U7601 ( .A(p_input[27720]), .B(p_input[17720]), .Z(n5068) );
  AND U7602 ( .A(p_input[7720]), .B(p_input[37720]), .Z(n5067) );
  AND U7603 ( .A(n5069), .B(n5070), .Z(o[771]) );
  AND U7604 ( .A(p_input[20771]), .B(p_input[10771]), .Z(n5070) );
  AND U7605 ( .A(p_input[771]), .B(p_input[30771]), .Z(n5069) );
  AND U7606 ( .A(n5071), .B(n5072), .Z(o[7719]) );
  AND U7607 ( .A(p_input[27719]), .B(p_input[17719]), .Z(n5072) );
  AND U7608 ( .A(p_input[7719]), .B(p_input[37719]), .Z(n5071) );
  AND U7609 ( .A(n5073), .B(n5074), .Z(o[7718]) );
  AND U7610 ( .A(p_input[27718]), .B(p_input[17718]), .Z(n5074) );
  AND U7611 ( .A(p_input[7718]), .B(p_input[37718]), .Z(n5073) );
  AND U7612 ( .A(n5075), .B(n5076), .Z(o[7717]) );
  AND U7613 ( .A(p_input[27717]), .B(p_input[17717]), .Z(n5076) );
  AND U7614 ( .A(p_input[7717]), .B(p_input[37717]), .Z(n5075) );
  AND U7615 ( .A(n5077), .B(n5078), .Z(o[7716]) );
  AND U7616 ( .A(p_input[27716]), .B(p_input[17716]), .Z(n5078) );
  AND U7617 ( .A(p_input[7716]), .B(p_input[37716]), .Z(n5077) );
  AND U7618 ( .A(n5079), .B(n5080), .Z(o[7715]) );
  AND U7619 ( .A(p_input[27715]), .B(p_input[17715]), .Z(n5080) );
  AND U7620 ( .A(p_input[7715]), .B(p_input[37715]), .Z(n5079) );
  AND U7621 ( .A(n5081), .B(n5082), .Z(o[7714]) );
  AND U7622 ( .A(p_input[27714]), .B(p_input[17714]), .Z(n5082) );
  AND U7623 ( .A(p_input[7714]), .B(p_input[37714]), .Z(n5081) );
  AND U7624 ( .A(n5083), .B(n5084), .Z(o[7713]) );
  AND U7625 ( .A(p_input[27713]), .B(p_input[17713]), .Z(n5084) );
  AND U7626 ( .A(p_input[7713]), .B(p_input[37713]), .Z(n5083) );
  AND U7627 ( .A(n5085), .B(n5086), .Z(o[7712]) );
  AND U7628 ( .A(p_input[27712]), .B(p_input[17712]), .Z(n5086) );
  AND U7629 ( .A(p_input[7712]), .B(p_input[37712]), .Z(n5085) );
  AND U7630 ( .A(n5087), .B(n5088), .Z(o[7711]) );
  AND U7631 ( .A(p_input[27711]), .B(p_input[17711]), .Z(n5088) );
  AND U7632 ( .A(p_input[7711]), .B(p_input[37711]), .Z(n5087) );
  AND U7633 ( .A(n5089), .B(n5090), .Z(o[7710]) );
  AND U7634 ( .A(p_input[27710]), .B(p_input[17710]), .Z(n5090) );
  AND U7635 ( .A(p_input[7710]), .B(p_input[37710]), .Z(n5089) );
  AND U7636 ( .A(n5091), .B(n5092), .Z(o[770]) );
  AND U7637 ( .A(p_input[20770]), .B(p_input[10770]), .Z(n5092) );
  AND U7638 ( .A(p_input[770]), .B(p_input[30770]), .Z(n5091) );
  AND U7639 ( .A(n5093), .B(n5094), .Z(o[7709]) );
  AND U7640 ( .A(p_input[27709]), .B(p_input[17709]), .Z(n5094) );
  AND U7641 ( .A(p_input[7709]), .B(p_input[37709]), .Z(n5093) );
  AND U7642 ( .A(n5095), .B(n5096), .Z(o[7708]) );
  AND U7643 ( .A(p_input[27708]), .B(p_input[17708]), .Z(n5096) );
  AND U7644 ( .A(p_input[7708]), .B(p_input[37708]), .Z(n5095) );
  AND U7645 ( .A(n5097), .B(n5098), .Z(o[7707]) );
  AND U7646 ( .A(p_input[27707]), .B(p_input[17707]), .Z(n5098) );
  AND U7647 ( .A(p_input[7707]), .B(p_input[37707]), .Z(n5097) );
  AND U7648 ( .A(n5099), .B(n5100), .Z(o[7706]) );
  AND U7649 ( .A(p_input[27706]), .B(p_input[17706]), .Z(n5100) );
  AND U7650 ( .A(p_input[7706]), .B(p_input[37706]), .Z(n5099) );
  AND U7651 ( .A(n5101), .B(n5102), .Z(o[7705]) );
  AND U7652 ( .A(p_input[27705]), .B(p_input[17705]), .Z(n5102) );
  AND U7653 ( .A(p_input[7705]), .B(p_input[37705]), .Z(n5101) );
  AND U7654 ( .A(n5103), .B(n5104), .Z(o[7704]) );
  AND U7655 ( .A(p_input[27704]), .B(p_input[17704]), .Z(n5104) );
  AND U7656 ( .A(p_input[7704]), .B(p_input[37704]), .Z(n5103) );
  AND U7657 ( .A(n5105), .B(n5106), .Z(o[7703]) );
  AND U7658 ( .A(p_input[27703]), .B(p_input[17703]), .Z(n5106) );
  AND U7659 ( .A(p_input[7703]), .B(p_input[37703]), .Z(n5105) );
  AND U7660 ( .A(n5107), .B(n5108), .Z(o[7702]) );
  AND U7661 ( .A(p_input[27702]), .B(p_input[17702]), .Z(n5108) );
  AND U7662 ( .A(p_input[7702]), .B(p_input[37702]), .Z(n5107) );
  AND U7663 ( .A(n5109), .B(n5110), .Z(o[7701]) );
  AND U7664 ( .A(p_input[27701]), .B(p_input[17701]), .Z(n5110) );
  AND U7665 ( .A(p_input[7701]), .B(p_input[37701]), .Z(n5109) );
  AND U7666 ( .A(n5111), .B(n5112), .Z(o[7700]) );
  AND U7667 ( .A(p_input[27700]), .B(p_input[17700]), .Z(n5112) );
  AND U7668 ( .A(p_input[7700]), .B(p_input[37700]), .Z(n5111) );
  AND U7669 ( .A(n5113), .B(n5114), .Z(o[76]) );
  AND U7670 ( .A(p_input[20076]), .B(p_input[10076]), .Z(n5114) );
  AND U7671 ( .A(p_input[76]), .B(p_input[30076]), .Z(n5113) );
  AND U7672 ( .A(n5115), .B(n5116), .Z(o[769]) );
  AND U7673 ( .A(p_input[20769]), .B(p_input[10769]), .Z(n5116) );
  AND U7674 ( .A(p_input[769]), .B(p_input[30769]), .Z(n5115) );
  AND U7675 ( .A(n5117), .B(n5118), .Z(o[7699]) );
  AND U7676 ( .A(p_input[27699]), .B(p_input[17699]), .Z(n5118) );
  AND U7677 ( .A(p_input[7699]), .B(p_input[37699]), .Z(n5117) );
  AND U7678 ( .A(n5119), .B(n5120), .Z(o[7698]) );
  AND U7679 ( .A(p_input[27698]), .B(p_input[17698]), .Z(n5120) );
  AND U7680 ( .A(p_input[7698]), .B(p_input[37698]), .Z(n5119) );
  AND U7681 ( .A(n5121), .B(n5122), .Z(o[7697]) );
  AND U7682 ( .A(p_input[27697]), .B(p_input[17697]), .Z(n5122) );
  AND U7683 ( .A(p_input[7697]), .B(p_input[37697]), .Z(n5121) );
  AND U7684 ( .A(n5123), .B(n5124), .Z(o[7696]) );
  AND U7685 ( .A(p_input[27696]), .B(p_input[17696]), .Z(n5124) );
  AND U7686 ( .A(p_input[7696]), .B(p_input[37696]), .Z(n5123) );
  AND U7687 ( .A(n5125), .B(n5126), .Z(o[7695]) );
  AND U7688 ( .A(p_input[27695]), .B(p_input[17695]), .Z(n5126) );
  AND U7689 ( .A(p_input[7695]), .B(p_input[37695]), .Z(n5125) );
  AND U7690 ( .A(n5127), .B(n5128), .Z(o[7694]) );
  AND U7691 ( .A(p_input[27694]), .B(p_input[17694]), .Z(n5128) );
  AND U7692 ( .A(p_input[7694]), .B(p_input[37694]), .Z(n5127) );
  AND U7693 ( .A(n5129), .B(n5130), .Z(o[7693]) );
  AND U7694 ( .A(p_input[27693]), .B(p_input[17693]), .Z(n5130) );
  AND U7695 ( .A(p_input[7693]), .B(p_input[37693]), .Z(n5129) );
  AND U7696 ( .A(n5131), .B(n5132), .Z(o[7692]) );
  AND U7697 ( .A(p_input[27692]), .B(p_input[17692]), .Z(n5132) );
  AND U7698 ( .A(p_input[7692]), .B(p_input[37692]), .Z(n5131) );
  AND U7699 ( .A(n5133), .B(n5134), .Z(o[7691]) );
  AND U7700 ( .A(p_input[27691]), .B(p_input[17691]), .Z(n5134) );
  AND U7701 ( .A(p_input[7691]), .B(p_input[37691]), .Z(n5133) );
  AND U7702 ( .A(n5135), .B(n5136), .Z(o[7690]) );
  AND U7703 ( .A(p_input[27690]), .B(p_input[17690]), .Z(n5136) );
  AND U7704 ( .A(p_input[7690]), .B(p_input[37690]), .Z(n5135) );
  AND U7705 ( .A(n5137), .B(n5138), .Z(o[768]) );
  AND U7706 ( .A(p_input[20768]), .B(p_input[10768]), .Z(n5138) );
  AND U7707 ( .A(p_input[768]), .B(p_input[30768]), .Z(n5137) );
  AND U7708 ( .A(n5139), .B(n5140), .Z(o[7689]) );
  AND U7709 ( .A(p_input[27689]), .B(p_input[17689]), .Z(n5140) );
  AND U7710 ( .A(p_input[7689]), .B(p_input[37689]), .Z(n5139) );
  AND U7711 ( .A(n5141), .B(n5142), .Z(o[7688]) );
  AND U7712 ( .A(p_input[27688]), .B(p_input[17688]), .Z(n5142) );
  AND U7713 ( .A(p_input[7688]), .B(p_input[37688]), .Z(n5141) );
  AND U7714 ( .A(n5143), .B(n5144), .Z(o[7687]) );
  AND U7715 ( .A(p_input[27687]), .B(p_input[17687]), .Z(n5144) );
  AND U7716 ( .A(p_input[7687]), .B(p_input[37687]), .Z(n5143) );
  AND U7717 ( .A(n5145), .B(n5146), .Z(o[7686]) );
  AND U7718 ( .A(p_input[27686]), .B(p_input[17686]), .Z(n5146) );
  AND U7719 ( .A(p_input[7686]), .B(p_input[37686]), .Z(n5145) );
  AND U7720 ( .A(n5147), .B(n5148), .Z(o[7685]) );
  AND U7721 ( .A(p_input[27685]), .B(p_input[17685]), .Z(n5148) );
  AND U7722 ( .A(p_input[7685]), .B(p_input[37685]), .Z(n5147) );
  AND U7723 ( .A(n5149), .B(n5150), .Z(o[7684]) );
  AND U7724 ( .A(p_input[27684]), .B(p_input[17684]), .Z(n5150) );
  AND U7725 ( .A(p_input[7684]), .B(p_input[37684]), .Z(n5149) );
  AND U7726 ( .A(n5151), .B(n5152), .Z(o[7683]) );
  AND U7727 ( .A(p_input[27683]), .B(p_input[17683]), .Z(n5152) );
  AND U7728 ( .A(p_input[7683]), .B(p_input[37683]), .Z(n5151) );
  AND U7729 ( .A(n5153), .B(n5154), .Z(o[7682]) );
  AND U7730 ( .A(p_input[27682]), .B(p_input[17682]), .Z(n5154) );
  AND U7731 ( .A(p_input[7682]), .B(p_input[37682]), .Z(n5153) );
  AND U7732 ( .A(n5155), .B(n5156), .Z(o[7681]) );
  AND U7733 ( .A(p_input[27681]), .B(p_input[17681]), .Z(n5156) );
  AND U7734 ( .A(p_input[7681]), .B(p_input[37681]), .Z(n5155) );
  AND U7735 ( .A(n5157), .B(n5158), .Z(o[7680]) );
  AND U7736 ( .A(p_input[27680]), .B(p_input[17680]), .Z(n5158) );
  AND U7737 ( .A(p_input[7680]), .B(p_input[37680]), .Z(n5157) );
  AND U7738 ( .A(n5159), .B(n5160), .Z(o[767]) );
  AND U7739 ( .A(p_input[20767]), .B(p_input[10767]), .Z(n5160) );
  AND U7740 ( .A(p_input[767]), .B(p_input[30767]), .Z(n5159) );
  AND U7741 ( .A(n5161), .B(n5162), .Z(o[7679]) );
  AND U7742 ( .A(p_input[27679]), .B(p_input[17679]), .Z(n5162) );
  AND U7743 ( .A(p_input[7679]), .B(p_input[37679]), .Z(n5161) );
  AND U7744 ( .A(n5163), .B(n5164), .Z(o[7678]) );
  AND U7745 ( .A(p_input[27678]), .B(p_input[17678]), .Z(n5164) );
  AND U7746 ( .A(p_input[7678]), .B(p_input[37678]), .Z(n5163) );
  AND U7747 ( .A(n5165), .B(n5166), .Z(o[7677]) );
  AND U7748 ( .A(p_input[27677]), .B(p_input[17677]), .Z(n5166) );
  AND U7749 ( .A(p_input[7677]), .B(p_input[37677]), .Z(n5165) );
  AND U7750 ( .A(n5167), .B(n5168), .Z(o[7676]) );
  AND U7751 ( .A(p_input[27676]), .B(p_input[17676]), .Z(n5168) );
  AND U7752 ( .A(p_input[7676]), .B(p_input[37676]), .Z(n5167) );
  AND U7753 ( .A(n5169), .B(n5170), .Z(o[7675]) );
  AND U7754 ( .A(p_input[27675]), .B(p_input[17675]), .Z(n5170) );
  AND U7755 ( .A(p_input[7675]), .B(p_input[37675]), .Z(n5169) );
  AND U7756 ( .A(n5171), .B(n5172), .Z(o[7674]) );
  AND U7757 ( .A(p_input[27674]), .B(p_input[17674]), .Z(n5172) );
  AND U7758 ( .A(p_input[7674]), .B(p_input[37674]), .Z(n5171) );
  AND U7759 ( .A(n5173), .B(n5174), .Z(o[7673]) );
  AND U7760 ( .A(p_input[27673]), .B(p_input[17673]), .Z(n5174) );
  AND U7761 ( .A(p_input[7673]), .B(p_input[37673]), .Z(n5173) );
  AND U7762 ( .A(n5175), .B(n5176), .Z(o[7672]) );
  AND U7763 ( .A(p_input[27672]), .B(p_input[17672]), .Z(n5176) );
  AND U7764 ( .A(p_input[7672]), .B(p_input[37672]), .Z(n5175) );
  AND U7765 ( .A(n5177), .B(n5178), .Z(o[7671]) );
  AND U7766 ( .A(p_input[27671]), .B(p_input[17671]), .Z(n5178) );
  AND U7767 ( .A(p_input[7671]), .B(p_input[37671]), .Z(n5177) );
  AND U7768 ( .A(n5179), .B(n5180), .Z(o[7670]) );
  AND U7769 ( .A(p_input[27670]), .B(p_input[17670]), .Z(n5180) );
  AND U7770 ( .A(p_input[7670]), .B(p_input[37670]), .Z(n5179) );
  AND U7771 ( .A(n5181), .B(n5182), .Z(o[766]) );
  AND U7772 ( .A(p_input[20766]), .B(p_input[10766]), .Z(n5182) );
  AND U7773 ( .A(p_input[766]), .B(p_input[30766]), .Z(n5181) );
  AND U7774 ( .A(n5183), .B(n5184), .Z(o[7669]) );
  AND U7775 ( .A(p_input[27669]), .B(p_input[17669]), .Z(n5184) );
  AND U7776 ( .A(p_input[7669]), .B(p_input[37669]), .Z(n5183) );
  AND U7777 ( .A(n5185), .B(n5186), .Z(o[7668]) );
  AND U7778 ( .A(p_input[27668]), .B(p_input[17668]), .Z(n5186) );
  AND U7779 ( .A(p_input[7668]), .B(p_input[37668]), .Z(n5185) );
  AND U7780 ( .A(n5187), .B(n5188), .Z(o[7667]) );
  AND U7781 ( .A(p_input[27667]), .B(p_input[17667]), .Z(n5188) );
  AND U7782 ( .A(p_input[7667]), .B(p_input[37667]), .Z(n5187) );
  AND U7783 ( .A(n5189), .B(n5190), .Z(o[7666]) );
  AND U7784 ( .A(p_input[27666]), .B(p_input[17666]), .Z(n5190) );
  AND U7785 ( .A(p_input[7666]), .B(p_input[37666]), .Z(n5189) );
  AND U7786 ( .A(n5191), .B(n5192), .Z(o[7665]) );
  AND U7787 ( .A(p_input[27665]), .B(p_input[17665]), .Z(n5192) );
  AND U7788 ( .A(p_input[7665]), .B(p_input[37665]), .Z(n5191) );
  AND U7789 ( .A(n5193), .B(n5194), .Z(o[7664]) );
  AND U7790 ( .A(p_input[27664]), .B(p_input[17664]), .Z(n5194) );
  AND U7791 ( .A(p_input[7664]), .B(p_input[37664]), .Z(n5193) );
  AND U7792 ( .A(n5195), .B(n5196), .Z(o[7663]) );
  AND U7793 ( .A(p_input[27663]), .B(p_input[17663]), .Z(n5196) );
  AND U7794 ( .A(p_input[7663]), .B(p_input[37663]), .Z(n5195) );
  AND U7795 ( .A(n5197), .B(n5198), .Z(o[7662]) );
  AND U7796 ( .A(p_input[27662]), .B(p_input[17662]), .Z(n5198) );
  AND U7797 ( .A(p_input[7662]), .B(p_input[37662]), .Z(n5197) );
  AND U7798 ( .A(n5199), .B(n5200), .Z(o[7661]) );
  AND U7799 ( .A(p_input[27661]), .B(p_input[17661]), .Z(n5200) );
  AND U7800 ( .A(p_input[7661]), .B(p_input[37661]), .Z(n5199) );
  AND U7801 ( .A(n5201), .B(n5202), .Z(o[7660]) );
  AND U7802 ( .A(p_input[27660]), .B(p_input[17660]), .Z(n5202) );
  AND U7803 ( .A(p_input[7660]), .B(p_input[37660]), .Z(n5201) );
  AND U7804 ( .A(n5203), .B(n5204), .Z(o[765]) );
  AND U7805 ( .A(p_input[20765]), .B(p_input[10765]), .Z(n5204) );
  AND U7806 ( .A(p_input[765]), .B(p_input[30765]), .Z(n5203) );
  AND U7807 ( .A(n5205), .B(n5206), .Z(o[7659]) );
  AND U7808 ( .A(p_input[27659]), .B(p_input[17659]), .Z(n5206) );
  AND U7809 ( .A(p_input[7659]), .B(p_input[37659]), .Z(n5205) );
  AND U7810 ( .A(n5207), .B(n5208), .Z(o[7658]) );
  AND U7811 ( .A(p_input[27658]), .B(p_input[17658]), .Z(n5208) );
  AND U7812 ( .A(p_input[7658]), .B(p_input[37658]), .Z(n5207) );
  AND U7813 ( .A(n5209), .B(n5210), .Z(o[7657]) );
  AND U7814 ( .A(p_input[27657]), .B(p_input[17657]), .Z(n5210) );
  AND U7815 ( .A(p_input[7657]), .B(p_input[37657]), .Z(n5209) );
  AND U7816 ( .A(n5211), .B(n5212), .Z(o[7656]) );
  AND U7817 ( .A(p_input[27656]), .B(p_input[17656]), .Z(n5212) );
  AND U7818 ( .A(p_input[7656]), .B(p_input[37656]), .Z(n5211) );
  AND U7819 ( .A(n5213), .B(n5214), .Z(o[7655]) );
  AND U7820 ( .A(p_input[27655]), .B(p_input[17655]), .Z(n5214) );
  AND U7821 ( .A(p_input[7655]), .B(p_input[37655]), .Z(n5213) );
  AND U7822 ( .A(n5215), .B(n5216), .Z(o[7654]) );
  AND U7823 ( .A(p_input[27654]), .B(p_input[17654]), .Z(n5216) );
  AND U7824 ( .A(p_input[7654]), .B(p_input[37654]), .Z(n5215) );
  AND U7825 ( .A(n5217), .B(n5218), .Z(o[7653]) );
  AND U7826 ( .A(p_input[27653]), .B(p_input[17653]), .Z(n5218) );
  AND U7827 ( .A(p_input[7653]), .B(p_input[37653]), .Z(n5217) );
  AND U7828 ( .A(n5219), .B(n5220), .Z(o[7652]) );
  AND U7829 ( .A(p_input[27652]), .B(p_input[17652]), .Z(n5220) );
  AND U7830 ( .A(p_input[7652]), .B(p_input[37652]), .Z(n5219) );
  AND U7831 ( .A(n5221), .B(n5222), .Z(o[7651]) );
  AND U7832 ( .A(p_input[27651]), .B(p_input[17651]), .Z(n5222) );
  AND U7833 ( .A(p_input[7651]), .B(p_input[37651]), .Z(n5221) );
  AND U7834 ( .A(n5223), .B(n5224), .Z(o[7650]) );
  AND U7835 ( .A(p_input[27650]), .B(p_input[17650]), .Z(n5224) );
  AND U7836 ( .A(p_input[7650]), .B(p_input[37650]), .Z(n5223) );
  AND U7837 ( .A(n5225), .B(n5226), .Z(o[764]) );
  AND U7838 ( .A(p_input[20764]), .B(p_input[10764]), .Z(n5226) );
  AND U7839 ( .A(p_input[764]), .B(p_input[30764]), .Z(n5225) );
  AND U7840 ( .A(n5227), .B(n5228), .Z(o[7649]) );
  AND U7841 ( .A(p_input[27649]), .B(p_input[17649]), .Z(n5228) );
  AND U7842 ( .A(p_input[7649]), .B(p_input[37649]), .Z(n5227) );
  AND U7843 ( .A(n5229), .B(n5230), .Z(o[7648]) );
  AND U7844 ( .A(p_input[27648]), .B(p_input[17648]), .Z(n5230) );
  AND U7845 ( .A(p_input[7648]), .B(p_input[37648]), .Z(n5229) );
  AND U7846 ( .A(n5231), .B(n5232), .Z(o[7647]) );
  AND U7847 ( .A(p_input[27647]), .B(p_input[17647]), .Z(n5232) );
  AND U7848 ( .A(p_input[7647]), .B(p_input[37647]), .Z(n5231) );
  AND U7849 ( .A(n5233), .B(n5234), .Z(o[7646]) );
  AND U7850 ( .A(p_input[27646]), .B(p_input[17646]), .Z(n5234) );
  AND U7851 ( .A(p_input[7646]), .B(p_input[37646]), .Z(n5233) );
  AND U7852 ( .A(n5235), .B(n5236), .Z(o[7645]) );
  AND U7853 ( .A(p_input[27645]), .B(p_input[17645]), .Z(n5236) );
  AND U7854 ( .A(p_input[7645]), .B(p_input[37645]), .Z(n5235) );
  AND U7855 ( .A(n5237), .B(n5238), .Z(o[7644]) );
  AND U7856 ( .A(p_input[27644]), .B(p_input[17644]), .Z(n5238) );
  AND U7857 ( .A(p_input[7644]), .B(p_input[37644]), .Z(n5237) );
  AND U7858 ( .A(n5239), .B(n5240), .Z(o[7643]) );
  AND U7859 ( .A(p_input[27643]), .B(p_input[17643]), .Z(n5240) );
  AND U7860 ( .A(p_input[7643]), .B(p_input[37643]), .Z(n5239) );
  AND U7861 ( .A(n5241), .B(n5242), .Z(o[7642]) );
  AND U7862 ( .A(p_input[27642]), .B(p_input[17642]), .Z(n5242) );
  AND U7863 ( .A(p_input[7642]), .B(p_input[37642]), .Z(n5241) );
  AND U7864 ( .A(n5243), .B(n5244), .Z(o[7641]) );
  AND U7865 ( .A(p_input[27641]), .B(p_input[17641]), .Z(n5244) );
  AND U7866 ( .A(p_input[7641]), .B(p_input[37641]), .Z(n5243) );
  AND U7867 ( .A(n5245), .B(n5246), .Z(o[7640]) );
  AND U7868 ( .A(p_input[27640]), .B(p_input[17640]), .Z(n5246) );
  AND U7869 ( .A(p_input[7640]), .B(p_input[37640]), .Z(n5245) );
  AND U7870 ( .A(n5247), .B(n5248), .Z(o[763]) );
  AND U7871 ( .A(p_input[20763]), .B(p_input[10763]), .Z(n5248) );
  AND U7872 ( .A(p_input[763]), .B(p_input[30763]), .Z(n5247) );
  AND U7873 ( .A(n5249), .B(n5250), .Z(o[7639]) );
  AND U7874 ( .A(p_input[27639]), .B(p_input[17639]), .Z(n5250) );
  AND U7875 ( .A(p_input[7639]), .B(p_input[37639]), .Z(n5249) );
  AND U7876 ( .A(n5251), .B(n5252), .Z(o[7638]) );
  AND U7877 ( .A(p_input[27638]), .B(p_input[17638]), .Z(n5252) );
  AND U7878 ( .A(p_input[7638]), .B(p_input[37638]), .Z(n5251) );
  AND U7879 ( .A(n5253), .B(n5254), .Z(o[7637]) );
  AND U7880 ( .A(p_input[27637]), .B(p_input[17637]), .Z(n5254) );
  AND U7881 ( .A(p_input[7637]), .B(p_input[37637]), .Z(n5253) );
  AND U7882 ( .A(n5255), .B(n5256), .Z(o[7636]) );
  AND U7883 ( .A(p_input[27636]), .B(p_input[17636]), .Z(n5256) );
  AND U7884 ( .A(p_input[7636]), .B(p_input[37636]), .Z(n5255) );
  AND U7885 ( .A(n5257), .B(n5258), .Z(o[7635]) );
  AND U7886 ( .A(p_input[27635]), .B(p_input[17635]), .Z(n5258) );
  AND U7887 ( .A(p_input[7635]), .B(p_input[37635]), .Z(n5257) );
  AND U7888 ( .A(n5259), .B(n5260), .Z(o[7634]) );
  AND U7889 ( .A(p_input[27634]), .B(p_input[17634]), .Z(n5260) );
  AND U7890 ( .A(p_input[7634]), .B(p_input[37634]), .Z(n5259) );
  AND U7891 ( .A(n5261), .B(n5262), .Z(o[7633]) );
  AND U7892 ( .A(p_input[27633]), .B(p_input[17633]), .Z(n5262) );
  AND U7893 ( .A(p_input[7633]), .B(p_input[37633]), .Z(n5261) );
  AND U7894 ( .A(n5263), .B(n5264), .Z(o[7632]) );
  AND U7895 ( .A(p_input[27632]), .B(p_input[17632]), .Z(n5264) );
  AND U7896 ( .A(p_input[7632]), .B(p_input[37632]), .Z(n5263) );
  AND U7897 ( .A(n5265), .B(n5266), .Z(o[7631]) );
  AND U7898 ( .A(p_input[27631]), .B(p_input[17631]), .Z(n5266) );
  AND U7899 ( .A(p_input[7631]), .B(p_input[37631]), .Z(n5265) );
  AND U7900 ( .A(n5267), .B(n5268), .Z(o[7630]) );
  AND U7901 ( .A(p_input[27630]), .B(p_input[17630]), .Z(n5268) );
  AND U7902 ( .A(p_input[7630]), .B(p_input[37630]), .Z(n5267) );
  AND U7903 ( .A(n5269), .B(n5270), .Z(o[762]) );
  AND U7904 ( .A(p_input[20762]), .B(p_input[10762]), .Z(n5270) );
  AND U7905 ( .A(p_input[762]), .B(p_input[30762]), .Z(n5269) );
  AND U7906 ( .A(n5271), .B(n5272), .Z(o[7629]) );
  AND U7907 ( .A(p_input[27629]), .B(p_input[17629]), .Z(n5272) );
  AND U7908 ( .A(p_input[7629]), .B(p_input[37629]), .Z(n5271) );
  AND U7909 ( .A(n5273), .B(n5274), .Z(o[7628]) );
  AND U7910 ( .A(p_input[27628]), .B(p_input[17628]), .Z(n5274) );
  AND U7911 ( .A(p_input[7628]), .B(p_input[37628]), .Z(n5273) );
  AND U7912 ( .A(n5275), .B(n5276), .Z(o[7627]) );
  AND U7913 ( .A(p_input[27627]), .B(p_input[17627]), .Z(n5276) );
  AND U7914 ( .A(p_input[7627]), .B(p_input[37627]), .Z(n5275) );
  AND U7915 ( .A(n5277), .B(n5278), .Z(o[7626]) );
  AND U7916 ( .A(p_input[27626]), .B(p_input[17626]), .Z(n5278) );
  AND U7917 ( .A(p_input[7626]), .B(p_input[37626]), .Z(n5277) );
  AND U7918 ( .A(n5279), .B(n5280), .Z(o[7625]) );
  AND U7919 ( .A(p_input[27625]), .B(p_input[17625]), .Z(n5280) );
  AND U7920 ( .A(p_input[7625]), .B(p_input[37625]), .Z(n5279) );
  AND U7921 ( .A(n5281), .B(n5282), .Z(o[7624]) );
  AND U7922 ( .A(p_input[27624]), .B(p_input[17624]), .Z(n5282) );
  AND U7923 ( .A(p_input[7624]), .B(p_input[37624]), .Z(n5281) );
  AND U7924 ( .A(n5283), .B(n5284), .Z(o[7623]) );
  AND U7925 ( .A(p_input[27623]), .B(p_input[17623]), .Z(n5284) );
  AND U7926 ( .A(p_input[7623]), .B(p_input[37623]), .Z(n5283) );
  AND U7927 ( .A(n5285), .B(n5286), .Z(o[7622]) );
  AND U7928 ( .A(p_input[27622]), .B(p_input[17622]), .Z(n5286) );
  AND U7929 ( .A(p_input[7622]), .B(p_input[37622]), .Z(n5285) );
  AND U7930 ( .A(n5287), .B(n5288), .Z(o[7621]) );
  AND U7931 ( .A(p_input[27621]), .B(p_input[17621]), .Z(n5288) );
  AND U7932 ( .A(p_input[7621]), .B(p_input[37621]), .Z(n5287) );
  AND U7933 ( .A(n5289), .B(n5290), .Z(o[7620]) );
  AND U7934 ( .A(p_input[27620]), .B(p_input[17620]), .Z(n5290) );
  AND U7935 ( .A(p_input[7620]), .B(p_input[37620]), .Z(n5289) );
  AND U7936 ( .A(n5291), .B(n5292), .Z(o[761]) );
  AND U7937 ( .A(p_input[20761]), .B(p_input[10761]), .Z(n5292) );
  AND U7938 ( .A(p_input[761]), .B(p_input[30761]), .Z(n5291) );
  AND U7939 ( .A(n5293), .B(n5294), .Z(o[7619]) );
  AND U7940 ( .A(p_input[27619]), .B(p_input[17619]), .Z(n5294) );
  AND U7941 ( .A(p_input[7619]), .B(p_input[37619]), .Z(n5293) );
  AND U7942 ( .A(n5295), .B(n5296), .Z(o[7618]) );
  AND U7943 ( .A(p_input[27618]), .B(p_input[17618]), .Z(n5296) );
  AND U7944 ( .A(p_input[7618]), .B(p_input[37618]), .Z(n5295) );
  AND U7945 ( .A(n5297), .B(n5298), .Z(o[7617]) );
  AND U7946 ( .A(p_input[27617]), .B(p_input[17617]), .Z(n5298) );
  AND U7947 ( .A(p_input[7617]), .B(p_input[37617]), .Z(n5297) );
  AND U7948 ( .A(n5299), .B(n5300), .Z(o[7616]) );
  AND U7949 ( .A(p_input[27616]), .B(p_input[17616]), .Z(n5300) );
  AND U7950 ( .A(p_input[7616]), .B(p_input[37616]), .Z(n5299) );
  AND U7951 ( .A(n5301), .B(n5302), .Z(o[7615]) );
  AND U7952 ( .A(p_input[27615]), .B(p_input[17615]), .Z(n5302) );
  AND U7953 ( .A(p_input[7615]), .B(p_input[37615]), .Z(n5301) );
  AND U7954 ( .A(n5303), .B(n5304), .Z(o[7614]) );
  AND U7955 ( .A(p_input[27614]), .B(p_input[17614]), .Z(n5304) );
  AND U7956 ( .A(p_input[7614]), .B(p_input[37614]), .Z(n5303) );
  AND U7957 ( .A(n5305), .B(n5306), .Z(o[7613]) );
  AND U7958 ( .A(p_input[27613]), .B(p_input[17613]), .Z(n5306) );
  AND U7959 ( .A(p_input[7613]), .B(p_input[37613]), .Z(n5305) );
  AND U7960 ( .A(n5307), .B(n5308), .Z(o[7612]) );
  AND U7961 ( .A(p_input[27612]), .B(p_input[17612]), .Z(n5308) );
  AND U7962 ( .A(p_input[7612]), .B(p_input[37612]), .Z(n5307) );
  AND U7963 ( .A(n5309), .B(n5310), .Z(o[7611]) );
  AND U7964 ( .A(p_input[27611]), .B(p_input[17611]), .Z(n5310) );
  AND U7965 ( .A(p_input[7611]), .B(p_input[37611]), .Z(n5309) );
  AND U7966 ( .A(n5311), .B(n5312), .Z(o[7610]) );
  AND U7967 ( .A(p_input[27610]), .B(p_input[17610]), .Z(n5312) );
  AND U7968 ( .A(p_input[7610]), .B(p_input[37610]), .Z(n5311) );
  AND U7969 ( .A(n5313), .B(n5314), .Z(o[760]) );
  AND U7970 ( .A(p_input[20760]), .B(p_input[10760]), .Z(n5314) );
  AND U7971 ( .A(p_input[760]), .B(p_input[30760]), .Z(n5313) );
  AND U7972 ( .A(n5315), .B(n5316), .Z(o[7609]) );
  AND U7973 ( .A(p_input[27609]), .B(p_input[17609]), .Z(n5316) );
  AND U7974 ( .A(p_input[7609]), .B(p_input[37609]), .Z(n5315) );
  AND U7975 ( .A(n5317), .B(n5318), .Z(o[7608]) );
  AND U7976 ( .A(p_input[27608]), .B(p_input[17608]), .Z(n5318) );
  AND U7977 ( .A(p_input[7608]), .B(p_input[37608]), .Z(n5317) );
  AND U7978 ( .A(n5319), .B(n5320), .Z(o[7607]) );
  AND U7979 ( .A(p_input[27607]), .B(p_input[17607]), .Z(n5320) );
  AND U7980 ( .A(p_input[7607]), .B(p_input[37607]), .Z(n5319) );
  AND U7981 ( .A(n5321), .B(n5322), .Z(o[7606]) );
  AND U7982 ( .A(p_input[27606]), .B(p_input[17606]), .Z(n5322) );
  AND U7983 ( .A(p_input[7606]), .B(p_input[37606]), .Z(n5321) );
  AND U7984 ( .A(n5323), .B(n5324), .Z(o[7605]) );
  AND U7985 ( .A(p_input[27605]), .B(p_input[17605]), .Z(n5324) );
  AND U7986 ( .A(p_input[7605]), .B(p_input[37605]), .Z(n5323) );
  AND U7987 ( .A(n5325), .B(n5326), .Z(o[7604]) );
  AND U7988 ( .A(p_input[27604]), .B(p_input[17604]), .Z(n5326) );
  AND U7989 ( .A(p_input[7604]), .B(p_input[37604]), .Z(n5325) );
  AND U7990 ( .A(n5327), .B(n5328), .Z(o[7603]) );
  AND U7991 ( .A(p_input[27603]), .B(p_input[17603]), .Z(n5328) );
  AND U7992 ( .A(p_input[7603]), .B(p_input[37603]), .Z(n5327) );
  AND U7993 ( .A(n5329), .B(n5330), .Z(o[7602]) );
  AND U7994 ( .A(p_input[27602]), .B(p_input[17602]), .Z(n5330) );
  AND U7995 ( .A(p_input[7602]), .B(p_input[37602]), .Z(n5329) );
  AND U7996 ( .A(n5331), .B(n5332), .Z(o[7601]) );
  AND U7997 ( .A(p_input[27601]), .B(p_input[17601]), .Z(n5332) );
  AND U7998 ( .A(p_input[7601]), .B(p_input[37601]), .Z(n5331) );
  AND U7999 ( .A(n5333), .B(n5334), .Z(o[7600]) );
  AND U8000 ( .A(p_input[27600]), .B(p_input[17600]), .Z(n5334) );
  AND U8001 ( .A(p_input[7600]), .B(p_input[37600]), .Z(n5333) );
  AND U8002 ( .A(n5335), .B(n5336), .Z(o[75]) );
  AND U8003 ( .A(p_input[20075]), .B(p_input[10075]), .Z(n5336) );
  AND U8004 ( .A(p_input[75]), .B(p_input[30075]), .Z(n5335) );
  AND U8005 ( .A(n5337), .B(n5338), .Z(o[759]) );
  AND U8006 ( .A(p_input[20759]), .B(p_input[10759]), .Z(n5338) );
  AND U8007 ( .A(p_input[759]), .B(p_input[30759]), .Z(n5337) );
  AND U8008 ( .A(n5339), .B(n5340), .Z(o[7599]) );
  AND U8009 ( .A(p_input[27599]), .B(p_input[17599]), .Z(n5340) );
  AND U8010 ( .A(p_input[7599]), .B(p_input[37599]), .Z(n5339) );
  AND U8011 ( .A(n5341), .B(n5342), .Z(o[7598]) );
  AND U8012 ( .A(p_input[27598]), .B(p_input[17598]), .Z(n5342) );
  AND U8013 ( .A(p_input[7598]), .B(p_input[37598]), .Z(n5341) );
  AND U8014 ( .A(n5343), .B(n5344), .Z(o[7597]) );
  AND U8015 ( .A(p_input[27597]), .B(p_input[17597]), .Z(n5344) );
  AND U8016 ( .A(p_input[7597]), .B(p_input[37597]), .Z(n5343) );
  AND U8017 ( .A(n5345), .B(n5346), .Z(o[7596]) );
  AND U8018 ( .A(p_input[27596]), .B(p_input[17596]), .Z(n5346) );
  AND U8019 ( .A(p_input[7596]), .B(p_input[37596]), .Z(n5345) );
  AND U8020 ( .A(n5347), .B(n5348), .Z(o[7595]) );
  AND U8021 ( .A(p_input[27595]), .B(p_input[17595]), .Z(n5348) );
  AND U8022 ( .A(p_input[7595]), .B(p_input[37595]), .Z(n5347) );
  AND U8023 ( .A(n5349), .B(n5350), .Z(o[7594]) );
  AND U8024 ( .A(p_input[27594]), .B(p_input[17594]), .Z(n5350) );
  AND U8025 ( .A(p_input[7594]), .B(p_input[37594]), .Z(n5349) );
  AND U8026 ( .A(n5351), .B(n5352), .Z(o[7593]) );
  AND U8027 ( .A(p_input[27593]), .B(p_input[17593]), .Z(n5352) );
  AND U8028 ( .A(p_input[7593]), .B(p_input[37593]), .Z(n5351) );
  AND U8029 ( .A(n5353), .B(n5354), .Z(o[7592]) );
  AND U8030 ( .A(p_input[27592]), .B(p_input[17592]), .Z(n5354) );
  AND U8031 ( .A(p_input[7592]), .B(p_input[37592]), .Z(n5353) );
  AND U8032 ( .A(n5355), .B(n5356), .Z(o[7591]) );
  AND U8033 ( .A(p_input[27591]), .B(p_input[17591]), .Z(n5356) );
  AND U8034 ( .A(p_input[7591]), .B(p_input[37591]), .Z(n5355) );
  AND U8035 ( .A(n5357), .B(n5358), .Z(o[7590]) );
  AND U8036 ( .A(p_input[27590]), .B(p_input[17590]), .Z(n5358) );
  AND U8037 ( .A(p_input[7590]), .B(p_input[37590]), .Z(n5357) );
  AND U8038 ( .A(n5359), .B(n5360), .Z(o[758]) );
  AND U8039 ( .A(p_input[20758]), .B(p_input[10758]), .Z(n5360) );
  AND U8040 ( .A(p_input[758]), .B(p_input[30758]), .Z(n5359) );
  AND U8041 ( .A(n5361), .B(n5362), .Z(o[7589]) );
  AND U8042 ( .A(p_input[27589]), .B(p_input[17589]), .Z(n5362) );
  AND U8043 ( .A(p_input[7589]), .B(p_input[37589]), .Z(n5361) );
  AND U8044 ( .A(n5363), .B(n5364), .Z(o[7588]) );
  AND U8045 ( .A(p_input[27588]), .B(p_input[17588]), .Z(n5364) );
  AND U8046 ( .A(p_input[7588]), .B(p_input[37588]), .Z(n5363) );
  AND U8047 ( .A(n5365), .B(n5366), .Z(o[7587]) );
  AND U8048 ( .A(p_input[27587]), .B(p_input[17587]), .Z(n5366) );
  AND U8049 ( .A(p_input[7587]), .B(p_input[37587]), .Z(n5365) );
  AND U8050 ( .A(n5367), .B(n5368), .Z(o[7586]) );
  AND U8051 ( .A(p_input[27586]), .B(p_input[17586]), .Z(n5368) );
  AND U8052 ( .A(p_input[7586]), .B(p_input[37586]), .Z(n5367) );
  AND U8053 ( .A(n5369), .B(n5370), .Z(o[7585]) );
  AND U8054 ( .A(p_input[27585]), .B(p_input[17585]), .Z(n5370) );
  AND U8055 ( .A(p_input[7585]), .B(p_input[37585]), .Z(n5369) );
  AND U8056 ( .A(n5371), .B(n5372), .Z(o[7584]) );
  AND U8057 ( .A(p_input[27584]), .B(p_input[17584]), .Z(n5372) );
  AND U8058 ( .A(p_input[7584]), .B(p_input[37584]), .Z(n5371) );
  AND U8059 ( .A(n5373), .B(n5374), .Z(o[7583]) );
  AND U8060 ( .A(p_input[27583]), .B(p_input[17583]), .Z(n5374) );
  AND U8061 ( .A(p_input[7583]), .B(p_input[37583]), .Z(n5373) );
  AND U8062 ( .A(n5375), .B(n5376), .Z(o[7582]) );
  AND U8063 ( .A(p_input[27582]), .B(p_input[17582]), .Z(n5376) );
  AND U8064 ( .A(p_input[7582]), .B(p_input[37582]), .Z(n5375) );
  AND U8065 ( .A(n5377), .B(n5378), .Z(o[7581]) );
  AND U8066 ( .A(p_input[27581]), .B(p_input[17581]), .Z(n5378) );
  AND U8067 ( .A(p_input[7581]), .B(p_input[37581]), .Z(n5377) );
  AND U8068 ( .A(n5379), .B(n5380), .Z(o[7580]) );
  AND U8069 ( .A(p_input[27580]), .B(p_input[17580]), .Z(n5380) );
  AND U8070 ( .A(p_input[7580]), .B(p_input[37580]), .Z(n5379) );
  AND U8071 ( .A(n5381), .B(n5382), .Z(o[757]) );
  AND U8072 ( .A(p_input[20757]), .B(p_input[10757]), .Z(n5382) );
  AND U8073 ( .A(p_input[757]), .B(p_input[30757]), .Z(n5381) );
  AND U8074 ( .A(n5383), .B(n5384), .Z(o[7579]) );
  AND U8075 ( .A(p_input[27579]), .B(p_input[17579]), .Z(n5384) );
  AND U8076 ( .A(p_input[7579]), .B(p_input[37579]), .Z(n5383) );
  AND U8077 ( .A(n5385), .B(n5386), .Z(o[7578]) );
  AND U8078 ( .A(p_input[27578]), .B(p_input[17578]), .Z(n5386) );
  AND U8079 ( .A(p_input[7578]), .B(p_input[37578]), .Z(n5385) );
  AND U8080 ( .A(n5387), .B(n5388), .Z(o[7577]) );
  AND U8081 ( .A(p_input[27577]), .B(p_input[17577]), .Z(n5388) );
  AND U8082 ( .A(p_input[7577]), .B(p_input[37577]), .Z(n5387) );
  AND U8083 ( .A(n5389), .B(n5390), .Z(o[7576]) );
  AND U8084 ( .A(p_input[27576]), .B(p_input[17576]), .Z(n5390) );
  AND U8085 ( .A(p_input[7576]), .B(p_input[37576]), .Z(n5389) );
  AND U8086 ( .A(n5391), .B(n5392), .Z(o[7575]) );
  AND U8087 ( .A(p_input[27575]), .B(p_input[17575]), .Z(n5392) );
  AND U8088 ( .A(p_input[7575]), .B(p_input[37575]), .Z(n5391) );
  AND U8089 ( .A(n5393), .B(n5394), .Z(o[7574]) );
  AND U8090 ( .A(p_input[27574]), .B(p_input[17574]), .Z(n5394) );
  AND U8091 ( .A(p_input[7574]), .B(p_input[37574]), .Z(n5393) );
  AND U8092 ( .A(n5395), .B(n5396), .Z(o[7573]) );
  AND U8093 ( .A(p_input[27573]), .B(p_input[17573]), .Z(n5396) );
  AND U8094 ( .A(p_input[7573]), .B(p_input[37573]), .Z(n5395) );
  AND U8095 ( .A(n5397), .B(n5398), .Z(o[7572]) );
  AND U8096 ( .A(p_input[27572]), .B(p_input[17572]), .Z(n5398) );
  AND U8097 ( .A(p_input[7572]), .B(p_input[37572]), .Z(n5397) );
  AND U8098 ( .A(n5399), .B(n5400), .Z(o[7571]) );
  AND U8099 ( .A(p_input[27571]), .B(p_input[17571]), .Z(n5400) );
  AND U8100 ( .A(p_input[7571]), .B(p_input[37571]), .Z(n5399) );
  AND U8101 ( .A(n5401), .B(n5402), .Z(o[7570]) );
  AND U8102 ( .A(p_input[27570]), .B(p_input[17570]), .Z(n5402) );
  AND U8103 ( .A(p_input[7570]), .B(p_input[37570]), .Z(n5401) );
  AND U8104 ( .A(n5403), .B(n5404), .Z(o[756]) );
  AND U8105 ( .A(p_input[20756]), .B(p_input[10756]), .Z(n5404) );
  AND U8106 ( .A(p_input[756]), .B(p_input[30756]), .Z(n5403) );
  AND U8107 ( .A(n5405), .B(n5406), .Z(o[7569]) );
  AND U8108 ( .A(p_input[27569]), .B(p_input[17569]), .Z(n5406) );
  AND U8109 ( .A(p_input[7569]), .B(p_input[37569]), .Z(n5405) );
  AND U8110 ( .A(n5407), .B(n5408), .Z(o[7568]) );
  AND U8111 ( .A(p_input[27568]), .B(p_input[17568]), .Z(n5408) );
  AND U8112 ( .A(p_input[7568]), .B(p_input[37568]), .Z(n5407) );
  AND U8113 ( .A(n5409), .B(n5410), .Z(o[7567]) );
  AND U8114 ( .A(p_input[27567]), .B(p_input[17567]), .Z(n5410) );
  AND U8115 ( .A(p_input[7567]), .B(p_input[37567]), .Z(n5409) );
  AND U8116 ( .A(n5411), .B(n5412), .Z(o[7566]) );
  AND U8117 ( .A(p_input[27566]), .B(p_input[17566]), .Z(n5412) );
  AND U8118 ( .A(p_input[7566]), .B(p_input[37566]), .Z(n5411) );
  AND U8119 ( .A(n5413), .B(n5414), .Z(o[7565]) );
  AND U8120 ( .A(p_input[27565]), .B(p_input[17565]), .Z(n5414) );
  AND U8121 ( .A(p_input[7565]), .B(p_input[37565]), .Z(n5413) );
  AND U8122 ( .A(n5415), .B(n5416), .Z(o[7564]) );
  AND U8123 ( .A(p_input[27564]), .B(p_input[17564]), .Z(n5416) );
  AND U8124 ( .A(p_input[7564]), .B(p_input[37564]), .Z(n5415) );
  AND U8125 ( .A(n5417), .B(n5418), .Z(o[7563]) );
  AND U8126 ( .A(p_input[27563]), .B(p_input[17563]), .Z(n5418) );
  AND U8127 ( .A(p_input[7563]), .B(p_input[37563]), .Z(n5417) );
  AND U8128 ( .A(n5419), .B(n5420), .Z(o[7562]) );
  AND U8129 ( .A(p_input[27562]), .B(p_input[17562]), .Z(n5420) );
  AND U8130 ( .A(p_input[7562]), .B(p_input[37562]), .Z(n5419) );
  AND U8131 ( .A(n5421), .B(n5422), .Z(o[7561]) );
  AND U8132 ( .A(p_input[27561]), .B(p_input[17561]), .Z(n5422) );
  AND U8133 ( .A(p_input[7561]), .B(p_input[37561]), .Z(n5421) );
  AND U8134 ( .A(n5423), .B(n5424), .Z(o[7560]) );
  AND U8135 ( .A(p_input[27560]), .B(p_input[17560]), .Z(n5424) );
  AND U8136 ( .A(p_input[7560]), .B(p_input[37560]), .Z(n5423) );
  AND U8137 ( .A(n5425), .B(n5426), .Z(o[755]) );
  AND U8138 ( .A(p_input[20755]), .B(p_input[10755]), .Z(n5426) );
  AND U8139 ( .A(p_input[755]), .B(p_input[30755]), .Z(n5425) );
  AND U8140 ( .A(n5427), .B(n5428), .Z(o[7559]) );
  AND U8141 ( .A(p_input[27559]), .B(p_input[17559]), .Z(n5428) );
  AND U8142 ( .A(p_input[7559]), .B(p_input[37559]), .Z(n5427) );
  AND U8143 ( .A(n5429), .B(n5430), .Z(o[7558]) );
  AND U8144 ( .A(p_input[27558]), .B(p_input[17558]), .Z(n5430) );
  AND U8145 ( .A(p_input[7558]), .B(p_input[37558]), .Z(n5429) );
  AND U8146 ( .A(n5431), .B(n5432), .Z(o[7557]) );
  AND U8147 ( .A(p_input[27557]), .B(p_input[17557]), .Z(n5432) );
  AND U8148 ( .A(p_input[7557]), .B(p_input[37557]), .Z(n5431) );
  AND U8149 ( .A(n5433), .B(n5434), .Z(o[7556]) );
  AND U8150 ( .A(p_input[27556]), .B(p_input[17556]), .Z(n5434) );
  AND U8151 ( .A(p_input[7556]), .B(p_input[37556]), .Z(n5433) );
  AND U8152 ( .A(n5435), .B(n5436), .Z(o[7555]) );
  AND U8153 ( .A(p_input[27555]), .B(p_input[17555]), .Z(n5436) );
  AND U8154 ( .A(p_input[7555]), .B(p_input[37555]), .Z(n5435) );
  AND U8155 ( .A(n5437), .B(n5438), .Z(o[7554]) );
  AND U8156 ( .A(p_input[27554]), .B(p_input[17554]), .Z(n5438) );
  AND U8157 ( .A(p_input[7554]), .B(p_input[37554]), .Z(n5437) );
  AND U8158 ( .A(n5439), .B(n5440), .Z(o[7553]) );
  AND U8159 ( .A(p_input[27553]), .B(p_input[17553]), .Z(n5440) );
  AND U8160 ( .A(p_input[7553]), .B(p_input[37553]), .Z(n5439) );
  AND U8161 ( .A(n5441), .B(n5442), .Z(o[7552]) );
  AND U8162 ( .A(p_input[27552]), .B(p_input[17552]), .Z(n5442) );
  AND U8163 ( .A(p_input[7552]), .B(p_input[37552]), .Z(n5441) );
  AND U8164 ( .A(n5443), .B(n5444), .Z(o[7551]) );
  AND U8165 ( .A(p_input[27551]), .B(p_input[17551]), .Z(n5444) );
  AND U8166 ( .A(p_input[7551]), .B(p_input[37551]), .Z(n5443) );
  AND U8167 ( .A(n5445), .B(n5446), .Z(o[7550]) );
  AND U8168 ( .A(p_input[27550]), .B(p_input[17550]), .Z(n5446) );
  AND U8169 ( .A(p_input[7550]), .B(p_input[37550]), .Z(n5445) );
  AND U8170 ( .A(n5447), .B(n5448), .Z(o[754]) );
  AND U8171 ( .A(p_input[20754]), .B(p_input[10754]), .Z(n5448) );
  AND U8172 ( .A(p_input[754]), .B(p_input[30754]), .Z(n5447) );
  AND U8173 ( .A(n5449), .B(n5450), .Z(o[7549]) );
  AND U8174 ( .A(p_input[27549]), .B(p_input[17549]), .Z(n5450) );
  AND U8175 ( .A(p_input[7549]), .B(p_input[37549]), .Z(n5449) );
  AND U8176 ( .A(n5451), .B(n5452), .Z(o[7548]) );
  AND U8177 ( .A(p_input[27548]), .B(p_input[17548]), .Z(n5452) );
  AND U8178 ( .A(p_input[7548]), .B(p_input[37548]), .Z(n5451) );
  AND U8179 ( .A(n5453), .B(n5454), .Z(o[7547]) );
  AND U8180 ( .A(p_input[27547]), .B(p_input[17547]), .Z(n5454) );
  AND U8181 ( .A(p_input[7547]), .B(p_input[37547]), .Z(n5453) );
  AND U8182 ( .A(n5455), .B(n5456), .Z(o[7546]) );
  AND U8183 ( .A(p_input[27546]), .B(p_input[17546]), .Z(n5456) );
  AND U8184 ( .A(p_input[7546]), .B(p_input[37546]), .Z(n5455) );
  AND U8185 ( .A(n5457), .B(n5458), .Z(o[7545]) );
  AND U8186 ( .A(p_input[27545]), .B(p_input[17545]), .Z(n5458) );
  AND U8187 ( .A(p_input[7545]), .B(p_input[37545]), .Z(n5457) );
  AND U8188 ( .A(n5459), .B(n5460), .Z(o[7544]) );
  AND U8189 ( .A(p_input[27544]), .B(p_input[17544]), .Z(n5460) );
  AND U8190 ( .A(p_input[7544]), .B(p_input[37544]), .Z(n5459) );
  AND U8191 ( .A(n5461), .B(n5462), .Z(o[7543]) );
  AND U8192 ( .A(p_input[27543]), .B(p_input[17543]), .Z(n5462) );
  AND U8193 ( .A(p_input[7543]), .B(p_input[37543]), .Z(n5461) );
  AND U8194 ( .A(n5463), .B(n5464), .Z(o[7542]) );
  AND U8195 ( .A(p_input[27542]), .B(p_input[17542]), .Z(n5464) );
  AND U8196 ( .A(p_input[7542]), .B(p_input[37542]), .Z(n5463) );
  AND U8197 ( .A(n5465), .B(n5466), .Z(o[7541]) );
  AND U8198 ( .A(p_input[27541]), .B(p_input[17541]), .Z(n5466) );
  AND U8199 ( .A(p_input[7541]), .B(p_input[37541]), .Z(n5465) );
  AND U8200 ( .A(n5467), .B(n5468), .Z(o[7540]) );
  AND U8201 ( .A(p_input[27540]), .B(p_input[17540]), .Z(n5468) );
  AND U8202 ( .A(p_input[7540]), .B(p_input[37540]), .Z(n5467) );
  AND U8203 ( .A(n5469), .B(n5470), .Z(o[753]) );
  AND U8204 ( .A(p_input[20753]), .B(p_input[10753]), .Z(n5470) );
  AND U8205 ( .A(p_input[753]), .B(p_input[30753]), .Z(n5469) );
  AND U8206 ( .A(n5471), .B(n5472), .Z(o[7539]) );
  AND U8207 ( .A(p_input[27539]), .B(p_input[17539]), .Z(n5472) );
  AND U8208 ( .A(p_input[7539]), .B(p_input[37539]), .Z(n5471) );
  AND U8209 ( .A(n5473), .B(n5474), .Z(o[7538]) );
  AND U8210 ( .A(p_input[27538]), .B(p_input[17538]), .Z(n5474) );
  AND U8211 ( .A(p_input[7538]), .B(p_input[37538]), .Z(n5473) );
  AND U8212 ( .A(n5475), .B(n5476), .Z(o[7537]) );
  AND U8213 ( .A(p_input[27537]), .B(p_input[17537]), .Z(n5476) );
  AND U8214 ( .A(p_input[7537]), .B(p_input[37537]), .Z(n5475) );
  AND U8215 ( .A(n5477), .B(n5478), .Z(o[7536]) );
  AND U8216 ( .A(p_input[27536]), .B(p_input[17536]), .Z(n5478) );
  AND U8217 ( .A(p_input[7536]), .B(p_input[37536]), .Z(n5477) );
  AND U8218 ( .A(n5479), .B(n5480), .Z(o[7535]) );
  AND U8219 ( .A(p_input[27535]), .B(p_input[17535]), .Z(n5480) );
  AND U8220 ( .A(p_input[7535]), .B(p_input[37535]), .Z(n5479) );
  AND U8221 ( .A(n5481), .B(n5482), .Z(o[7534]) );
  AND U8222 ( .A(p_input[27534]), .B(p_input[17534]), .Z(n5482) );
  AND U8223 ( .A(p_input[7534]), .B(p_input[37534]), .Z(n5481) );
  AND U8224 ( .A(n5483), .B(n5484), .Z(o[7533]) );
  AND U8225 ( .A(p_input[27533]), .B(p_input[17533]), .Z(n5484) );
  AND U8226 ( .A(p_input[7533]), .B(p_input[37533]), .Z(n5483) );
  AND U8227 ( .A(n5485), .B(n5486), .Z(o[7532]) );
  AND U8228 ( .A(p_input[27532]), .B(p_input[17532]), .Z(n5486) );
  AND U8229 ( .A(p_input[7532]), .B(p_input[37532]), .Z(n5485) );
  AND U8230 ( .A(n5487), .B(n5488), .Z(o[7531]) );
  AND U8231 ( .A(p_input[27531]), .B(p_input[17531]), .Z(n5488) );
  AND U8232 ( .A(p_input[7531]), .B(p_input[37531]), .Z(n5487) );
  AND U8233 ( .A(n5489), .B(n5490), .Z(o[7530]) );
  AND U8234 ( .A(p_input[27530]), .B(p_input[17530]), .Z(n5490) );
  AND U8235 ( .A(p_input[7530]), .B(p_input[37530]), .Z(n5489) );
  AND U8236 ( .A(n5491), .B(n5492), .Z(o[752]) );
  AND U8237 ( .A(p_input[20752]), .B(p_input[10752]), .Z(n5492) );
  AND U8238 ( .A(p_input[752]), .B(p_input[30752]), .Z(n5491) );
  AND U8239 ( .A(n5493), .B(n5494), .Z(o[7529]) );
  AND U8240 ( .A(p_input[27529]), .B(p_input[17529]), .Z(n5494) );
  AND U8241 ( .A(p_input[7529]), .B(p_input[37529]), .Z(n5493) );
  AND U8242 ( .A(n5495), .B(n5496), .Z(o[7528]) );
  AND U8243 ( .A(p_input[27528]), .B(p_input[17528]), .Z(n5496) );
  AND U8244 ( .A(p_input[7528]), .B(p_input[37528]), .Z(n5495) );
  AND U8245 ( .A(n5497), .B(n5498), .Z(o[7527]) );
  AND U8246 ( .A(p_input[27527]), .B(p_input[17527]), .Z(n5498) );
  AND U8247 ( .A(p_input[7527]), .B(p_input[37527]), .Z(n5497) );
  AND U8248 ( .A(n5499), .B(n5500), .Z(o[7526]) );
  AND U8249 ( .A(p_input[27526]), .B(p_input[17526]), .Z(n5500) );
  AND U8250 ( .A(p_input[7526]), .B(p_input[37526]), .Z(n5499) );
  AND U8251 ( .A(n5501), .B(n5502), .Z(o[7525]) );
  AND U8252 ( .A(p_input[27525]), .B(p_input[17525]), .Z(n5502) );
  AND U8253 ( .A(p_input[7525]), .B(p_input[37525]), .Z(n5501) );
  AND U8254 ( .A(n5503), .B(n5504), .Z(o[7524]) );
  AND U8255 ( .A(p_input[27524]), .B(p_input[17524]), .Z(n5504) );
  AND U8256 ( .A(p_input[7524]), .B(p_input[37524]), .Z(n5503) );
  AND U8257 ( .A(n5505), .B(n5506), .Z(o[7523]) );
  AND U8258 ( .A(p_input[27523]), .B(p_input[17523]), .Z(n5506) );
  AND U8259 ( .A(p_input[7523]), .B(p_input[37523]), .Z(n5505) );
  AND U8260 ( .A(n5507), .B(n5508), .Z(o[7522]) );
  AND U8261 ( .A(p_input[27522]), .B(p_input[17522]), .Z(n5508) );
  AND U8262 ( .A(p_input[7522]), .B(p_input[37522]), .Z(n5507) );
  AND U8263 ( .A(n5509), .B(n5510), .Z(o[7521]) );
  AND U8264 ( .A(p_input[27521]), .B(p_input[17521]), .Z(n5510) );
  AND U8265 ( .A(p_input[7521]), .B(p_input[37521]), .Z(n5509) );
  AND U8266 ( .A(n5511), .B(n5512), .Z(o[7520]) );
  AND U8267 ( .A(p_input[27520]), .B(p_input[17520]), .Z(n5512) );
  AND U8268 ( .A(p_input[7520]), .B(p_input[37520]), .Z(n5511) );
  AND U8269 ( .A(n5513), .B(n5514), .Z(o[751]) );
  AND U8270 ( .A(p_input[20751]), .B(p_input[10751]), .Z(n5514) );
  AND U8271 ( .A(p_input[751]), .B(p_input[30751]), .Z(n5513) );
  AND U8272 ( .A(n5515), .B(n5516), .Z(o[7519]) );
  AND U8273 ( .A(p_input[27519]), .B(p_input[17519]), .Z(n5516) );
  AND U8274 ( .A(p_input[7519]), .B(p_input[37519]), .Z(n5515) );
  AND U8275 ( .A(n5517), .B(n5518), .Z(o[7518]) );
  AND U8276 ( .A(p_input[27518]), .B(p_input[17518]), .Z(n5518) );
  AND U8277 ( .A(p_input[7518]), .B(p_input[37518]), .Z(n5517) );
  AND U8278 ( .A(n5519), .B(n5520), .Z(o[7517]) );
  AND U8279 ( .A(p_input[27517]), .B(p_input[17517]), .Z(n5520) );
  AND U8280 ( .A(p_input[7517]), .B(p_input[37517]), .Z(n5519) );
  AND U8281 ( .A(n5521), .B(n5522), .Z(o[7516]) );
  AND U8282 ( .A(p_input[27516]), .B(p_input[17516]), .Z(n5522) );
  AND U8283 ( .A(p_input[7516]), .B(p_input[37516]), .Z(n5521) );
  AND U8284 ( .A(n5523), .B(n5524), .Z(o[7515]) );
  AND U8285 ( .A(p_input[27515]), .B(p_input[17515]), .Z(n5524) );
  AND U8286 ( .A(p_input[7515]), .B(p_input[37515]), .Z(n5523) );
  AND U8287 ( .A(n5525), .B(n5526), .Z(o[7514]) );
  AND U8288 ( .A(p_input[27514]), .B(p_input[17514]), .Z(n5526) );
  AND U8289 ( .A(p_input[7514]), .B(p_input[37514]), .Z(n5525) );
  AND U8290 ( .A(n5527), .B(n5528), .Z(o[7513]) );
  AND U8291 ( .A(p_input[27513]), .B(p_input[17513]), .Z(n5528) );
  AND U8292 ( .A(p_input[7513]), .B(p_input[37513]), .Z(n5527) );
  AND U8293 ( .A(n5529), .B(n5530), .Z(o[7512]) );
  AND U8294 ( .A(p_input[27512]), .B(p_input[17512]), .Z(n5530) );
  AND U8295 ( .A(p_input[7512]), .B(p_input[37512]), .Z(n5529) );
  AND U8296 ( .A(n5531), .B(n5532), .Z(o[7511]) );
  AND U8297 ( .A(p_input[27511]), .B(p_input[17511]), .Z(n5532) );
  AND U8298 ( .A(p_input[7511]), .B(p_input[37511]), .Z(n5531) );
  AND U8299 ( .A(n5533), .B(n5534), .Z(o[7510]) );
  AND U8300 ( .A(p_input[27510]), .B(p_input[17510]), .Z(n5534) );
  AND U8301 ( .A(p_input[7510]), .B(p_input[37510]), .Z(n5533) );
  AND U8302 ( .A(n5535), .B(n5536), .Z(o[750]) );
  AND U8303 ( .A(p_input[20750]), .B(p_input[10750]), .Z(n5536) );
  AND U8304 ( .A(p_input[750]), .B(p_input[30750]), .Z(n5535) );
  AND U8305 ( .A(n5537), .B(n5538), .Z(o[7509]) );
  AND U8306 ( .A(p_input[27509]), .B(p_input[17509]), .Z(n5538) );
  AND U8307 ( .A(p_input[7509]), .B(p_input[37509]), .Z(n5537) );
  AND U8308 ( .A(n5539), .B(n5540), .Z(o[7508]) );
  AND U8309 ( .A(p_input[27508]), .B(p_input[17508]), .Z(n5540) );
  AND U8310 ( .A(p_input[7508]), .B(p_input[37508]), .Z(n5539) );
  AND U8311 ( .A(n5541), .B(n5542), .Z(o[7507]) );
  AND U8312 ( .A(p_input[27507]), .B(p_input[17507]), .Z(n5542) );
  AND U8313 ( .A(p_input[7507]), .B(p_input[37507]), .Z(n5541) );
  AND U8314 ( .A(n5543), .B(n5544), .Z(o[7506]) );
  AND U8315 ( .A(p_input[27506]), .B(p_input[17506]), .Z(n5544) );
  AND U8316 ( .A(p_input[7506]), .B(p_input[37506]), .Z(n5543) );
  AND U8317 ( .A(n5545), .B(n5546), .Z(o[7505]) );
  AND U8318 ( .A(p_input[27505]), .B(p_input[17505]), .Z(n5546) );
  AND U8319 ( .A(p_input[7505]), .B(p_input[37505]), .Z(n5545) );
  AND U8320 ( .A(n5547), .B(n5548), .Z(o[7504]) );
  AND U8321 ( .A(p_input[27504]), .B(p_input[17504]), .Z(n5548) );
  AND U8322 ( .A(p_input[7504]), .B(p_input[37504]), .Z(n5547) );
  AND U8323 ( .A(n5549), .B(n5550), .Z(o[7503]) );
  AND U8324 ( .A(p_input[27503]), .B(p_input[17503]), .Z(n5550) );
  AND U8325 ( .A(p_input[7503]), .B(p_input[37503]), .Z(n5549) );
  AND U8326 ( .A(n5551), .B(n5552), .Z(o[7502]) );
  AND U8327 ( .A(p_input[27502]), .B(p_input[17502]), .Z(n5552) );
  AND U8328 ( .A(p_input[7502]), .B(p_input[37502]), .Z(n5551) );
  AND U8329 ( .A(n5553), .B(n5554), .Z(o[7501]) );
  AND U8330 ( .A(p_input[27501]), .B(p_input[17501]), .Z(n5554) );
  AND U8331 ( .A(p_input[7501]), .B(p_input[37501]), .Z(n5553) );
  AND U8332 ( .A(n5555), .B(n5556), .Z(o[7500]) );
  AND U8333 ( .A(p_input[27500]), .B(p_input[17500]), .Z(n5556) );
  AND U8334 ( .A(p_input[7500]), .B(p_input[37500]), .Z(n5555) );
  AND U8335 ( .A(n5557), .B(n5558), .Z(o[74]) );
  AND U8336 ( .A(p_input[20074]), .B(p_input[10074]), .Z(n5558) );
  AND U8337 ( .A(p_input[74]), .B(p_input[30074]), .Z(n5557) );
  AND U8338 ( .A(n5559), .B(n5560), .Z(o[749]) );
  AND U8339 ( .A(p_input[20749]), .B(p_input[10749]), .Z(n5560) );
  AND U8340 ( .A(p_input[749]), .B(p_input[30749]), .Z(n5559) );
  AND U8341 ( .A(n5561), .B(n5562), .Z(o[7499]) );
  AND U8342 ( .A(p_input[27499]), .B(p_input[17499]), .Z(n5562) );
  AND U8343 ( .A(p_input[7499]), .B(p_input[37499]), .Z(n5561) );
  AND U8344 ( .A(n5563), .B(n5564), .Z(o[7498]) );
  AND U8345 ( .A(p_input[27498]), .B(p_input[17498]), .Z(n5564) );
  AND U8346 ( .A(p_input[7498]), .B(p_input[37498]), .Z(n5563) );
  AND U8347 ( .A(n5565), .B(n5566), .Z(o[7497]) );
  AND U8348 ( .A(p_input[27497]), .B(p_input[17497]), .Z(n5566) );
  AND U8349 ( .A(p_input[7497]), .B(p_input[37497]), .Z(n5565) );
  AND U8350 ( .A(n5567), .B(n5568), .Z(o[7496]) );
  AND U8351 ( .A(p_input[27496]), .B(p_input[17496]), .Z(n5568) );
  AND U8352 ( .A(p_input[7496]), .B(p_input[37496]), .Z(n5567) );
  AND U8353 ( .A(n5569), .B(n5570), .Z(o[7495]) );
  AND U8354 ( .A(p_input[27495]), .B(p_input[17495]), .Z(n5570) );
  AND U8355 ( .A(p_input[7495]), .B(p_input[37495]), .Z(n5569) );
  AND U8356 ( .A(n5571), .B(n5572), .Z(o[7494]) );
  AND U8357 ( .A(p_input[27494]), .B(p_input[17494]), .Z(n5572) );
  AND U8358 ( .A(p_input[7494]), .B(p_input[37494]), .Z(n5571) );
  AND U8359 ( .A(n5573), .B(n5574), .Z(o[7493]) );
  AND U8360 ( .A(p_input[27493]), .B(p_input[17493]), .Z(n5574) );
  AND U8361 ( .A(p_input[7493]), .B(p_input[37493]), .Z(n5573) );
  AND U8362 ( .A(n5575), .B(n5576), .Z(o[7492]) );
  AND U8363 ( .A(p_input[27492]), .B(p_input[17492]), .Z(n5576) );
  AND U8364 ( .A(p_input[7492]), .B(p_input[37492]), .Z(n5575) );
  AND U8365 ( .A(n5577), .B(n5578), .Z(o[7491]) );
  AND U8366 ( .A(p_input[27491]), .B(p_input[17491]), .Z(n5578) );
  AND U8367 ( .A(p_input[7491]), .B(p_input[37491]), .Z(n5577) );
  AND U8368 ( .A(n5579), .B(n5580), .Z(o[7490]) );
  AND U8369 ( .A(p_input[27490]), .B(p_input[17490]), .Z(n5580) );
  AND U8370 ( .A(p_input[7490]), .B(p_input[37490]), .Z(n5579) );
  AND U8371 ( .A(n5581), .B(n5582), .Z(o[748]) );
  AND U8372 ( .A(p_input[20748]), .B(p_input[10748]), .Z(n5582) );
  AND U8373 ( .A(p_input[748]), .B(p_input[30748]), .Z(n5581) );
  AND U8374 ( .A(n5583), .B(n5584), .Z(o[7489]) );
  AND U8375 ( .A(p_input[27489]), .B(p_input[17489]), .Z(n5584) );
  AND U8376 ( .A(p_input[7489]), .B(p_input[37489]), .Z(n5583) );
  AND U8377 ( .A(n5585), .B(n5586), .Z(o[7488]) );
  AND U8378 ( .A(p_input[27488]), .B(p_input[17488]), .Z(n5586) );
  AND U8379 ( .A(p_input[7488]), .B(p_input[37488]), .Z(n5585) );
  AND U8380 ( .A(n5587), .B(n5588), .Z(o[7487]) );
  AND U8381 ( .A(p_input[27487]), .B(p_input[17487]), .Z(n5588) );
  AND U8382 ( .A(p_input[7487]), .B(p_input[37487]), .Z(n5587) );
  AND U8383 ( .A(n5589), .B(n5590), .Z(o[7486]) );
  AND U8384 ( .A(p_input[27486]), .B(p_input[17486]), .Z(n5590) );
  AND U8385 ( .A(p_input[7486]), .B(p_input[37486]), .Z(n5589) );
  AND U8386 ( .A(n5591), .B(n5592), .Z(o[7485]) );
  AND U8387 ( .A(p_input[27485]), .B(p_input[17485]), .Z(n5592) );
  AND U8388 ( .A(p_input[7485]), .B(p_input[37485]), .Z(n5591) );
  AND U8389 ( .A(n5593), .B(n5594), .Z(o[7484]) );
  AND U8390 ( .A(p_input[27484]), .B(p_input[17484]), .Z(n5594) );
  AND U8391 ( .A(p_input[7484]), .B(p_input[37484]), .Z(n5593) );
  AND U8392 ( .A(n5595), .B(n5596), .Z(o[7483]) );
  AND U8393 ( .A(p_input[27483]), .B(p_input[17483]), .Z(n5596) );
  AND U8394 ( .A(p_input[7483]), .B(p_input[37483]), .Z(n5595) );
  AND U8395 ( .A(n5597), .B(n5598), .Z(o[7482]) );
  AND U8396 ( .A(p_input[27482]), .B(p_input[17482]), .Z(n5598) );
  AND U8397 ( .A(p_input[7482]), .B(p_input[37482]), .Z(n5597) );
  AND U8398 ( .A(n5599), .B(n5600), .Z(o[7481]) );
  AND U8399 ( .A(p_input[27481]), .B(p_input[17481]), .Z(n5600) );
  AND U8400 ( .A(p_input[7481]), .B(p_input[37481]), .Z(n5599) );
  AND U8401 ( .A(n5601), .B(n5602), .Z(o[7480]) );
  AND U8402 ( .A(p_input[27480]), .B(p_input[17480]), .Z(n5602) );
  AND U8403 ( .A(p_input[7480]), .B(p_input[37480]), .Z(n5601) );
  AND U8404 ( .A(n5603), .B(n5604), .Z(o[747]) );
  AND U8405 ( .A(p_input[20747]), .B(p_input[10747]), .Z(n5604) );
  AND U8406 ( .A(p_input[747]), .B(p_input[30747]), .Z(n5603) );
  AND U8407 ( .A(n5605), .B(n5606), .Z(o[7479]) );
  AND U8408 ( .A(p_input[27479]), .B(p_input[17479]), .Z(n5606) );
  AND U8409 ( .A(p_input[7479]), .B(p_input[37479]), .Z(n5605) );
  AND U8410 ( .A(n5607), .B(n5608), .Z(o[7478]) );
  AND U8411 ( .A(p_input[27478]), .B(p_input[17478]), .Z(n5608) );
  AND U8412 ( .A(p_input[7478]), .B(p_input[37478]), .Z(n5607) );
  AND U8413 ( .A(n5609), .B(n5610), .Z(o[7477]) );
  AND U8414 ( .A(p_input[27477]), .B(p_input[17477]), .Z(n5610) );
  AND U8415 ( .A(p_input[7477]), .B(p_input[37477]), .Z(n5609) );
  AND U8416 ( .A(n5611), .B(n5612), .Z(o[7476]) );
  AND U8417 ( .A(p_input[27476]), .B(p_input[17476]), .Z(n5612) );
  AND U8418 ( .A(p_input[7476]), .B(p_input[37476]), .Z(n5611) );
  AND U8419 ( .A(n5613), .B(n5614), .Z(o[7475]) );
  AND U8420 ( .A(p_input[27475]), .B(p_input[17475]), .Z(n5614) );
  AND U8421 ( .A(p_input[7475]), .B(p_input[37475]), .Z(n5613) );
  AND U8422 ( .A(n5615), .B(n5616), .Z(o[7474]) );
  AND U8423 ( .A(p_input[27474]), .B(p_input[17474]), .Z(n5616) );
  AND U8424 ( .A(p_input[7474]), .B(p_input[37474]), .Z(n5615) );
  AND U8425 ( .A(n5617), .B(n5618), .Z(o[7473]) );
  AND U8426 ( .A(p_input[27473]), .B(p_input[17473]), .Z(n5618) );
  AND U8427 ( .A(p_input[7473]), .B(p_input[37473]), .Z(n5617) );
  AND U8428 ( .A(n5619), .B(n5620), .Z(o[7472]) );
  AND U8429 ( .A(p_input[27472]), .B(p_input[17472]), .Z(n5620) );
  AND U8430 ( .A(p_input[7472]), .B(p_input[37472]), .Z(n5619) );
  AND U8431 ( .A(n5621), .B(n5622), .Z(o[7471]) );
  AND U8432 ( .A(p_input[27471]), .B(p_input[17471]), .Z(n5622) );
  AND U8433 ( .A(p_input[7471]), .B(p_input[37471]), .Z(n5621) );
  AND U8434 ( .A(n5623), .B(n5624), .Z(o[7470]) );
  AND U8435 ( .A(p_input[27470]), .B(p_input[17470]), .Z(n5624) );
  AND U8436 ( .A(p_input[7470]), .B(p_input[37470]), .Z(n5623) );
  AND U8437 ( .A(n5625), .B(n5626), .Z(o[746]) );
  AND U8438 ( .A(p_input[20746]), .B(p_input[10746]), .Z(n5626) );
  AND U8439 ( .A(p_input[746]), .B(p_input[30746]), .Z(n5625) );
  AND U8440 ( .A(n5627), .B(n5628), .Z(o[7469]) );
  AND U8441 ( .A(p_input[27469]), .B(p_input[17469]), .Z(n5628) );
  AND U8442 ( .A(p_input[7469]), .B(p_input[37469]), .Z(n5627) );
  AND U8443 ( .A(n5629), .B(n5630), .Z(o[7468]) );
  AND U8444 ( .A(p_input[27468]), .B(p_input[17468]), .Z(n5630) );
  AND U8445 ( .A(p_input[7468]), .B(p_input[37468]), .Z(n5629) );
  AND U8446 ( .A(n5631), .B(n5632), .Z(o[7467]) );
  AND U8447 ( .A(p_input[27467]), .B(p_input[17467]), .Z(n5632) );
  AND U8448 ( .A(p_input[7467]), .B(p_input[37467]), .Z(n5631) );
  AND U8449 ( .A(n5633), .B(n5634), .Z(o[7466]) );
  AND U8450 ( .A(p_input[27466]), .B(p_input[17466]), .Z(n5634) );
  AND U8451 ( .A(p_input[7466]), .B(p_input[37466]), .Z(n5633) );
  AND U8452 ( .A(n5635), .B(n5636), .Z(o[7465]) );
  AND U8453 ( .A(p_input[27465]), .B(p_input[17465]), .Z(n5636) );
  AND U8454 ( .A(p_input[7465]), .B(p_input[37465]), .Z(n5635) );
  AND U8455 ( .A(n5637), .B(n5638), .Z(o[7464]) );
  AND U8456 ( .A(p_input[27464]), .B(p_input[17464]), .Z(n5638) );
  AND U8457 ( .A(p_input[7464]), .B(p_input[37464]), .Z(n5637) );
  AND U8458 ( .A(n5639), .B(n5640), .Z(o[7463]) );
  AND U8459 ( .A(p_input[27463]), .B(p_input[17463]), .Z(n5640) );
  AND U8460 ( .A(p_input[7463]), .B(p_input[37463]), .Z(n5639) );
  AND U8461 ( .A(n5641), .B(n5642), .Z(o[7462]) );
  AND U8462 ( .A(p_input[27462]), .B(p_input[17462]), .Z(n5642) );
  AND U8463 ( .A(p_input[7462]), .B(p_input[37462]), .Z(n5641) );
  AND U8464 ( .A(n5643), .B(n5644), .Z(o[7461]) );
  AND U8465 ( .A(p_input[27461]), .B(p_input[17461]), .Z(n5644) );
  AND U8466 ( .A(p_input[7461]), .B(p_input[37461]), .Z(n5643) );
  AND U8467 ( .A(n5645), .B(n5646), .Z(o[7460]) );
  AND U8468 ( .A(p_input[27460]), .B(p_input[17460]), .Z(n5646) );
  AND U8469 ( .A(p_input[7460]), .B(p_input[37460]), .Z(n5645) );
  AND U8470 ( .A(n5647), .B(n5648), .Z(o[745]) );
  AND U8471 ( .A(p_input[20745]), .B(p_input[10745]), .Z(n5648) );
  AND U8472 ( .A(p_input[745]), .B(p_input[30745]), .Z(n5647) );
  AND U8473 ( .A(n5649), .B(n5650), .Z(o[7459]) );
  AND U8474 ( .A(p_input[27459]), .B(p_input[17459]), .Z(n5650) );
  AND U8475 ( .A(p_input[7459]), .B(p_input[37459]), .Z(n5649) );
  AND U8476 ( .A(n5651), .B(n5652), .Z(o[7458]) );
  AND U8477 ( .A(p_input[27458]), .B(p_input[17458]), .Z(n5652) );
  AND U8478 ( .A(p_input[7458]), .B(p_input[37458]), .Z(n5651) );
  AND U8479 ( .A(n5653), .B(n5654), .Z(o[7457]) );
  AND U8480 ( .A(p_input[27457]), .B(p_input[17457]), .Z(n5654) );
  AND U8481 ( .A(p_input[7457]), .B(p_input[37457]), .Z(n5653) );
  AND U8482 ( .A(n5655), .B(n5656), .Z(o[7456]) );
  AND U8483 ( .A(p_input[27456]), .B(p_input[17456]), .Z(n5656) );
  AND U8484 ( .A(p_input[7456]), .B(p_input[37456]), .Z(n5655) );
  AND U8485 ( .A(n5657), .B(n5658), .Z(o[7455]) );
  AND U8486 ( .A(p_input[27455]), .B(p_input[17455]), .Z(n5658) );
  AND U8487 ( .A(p_input[7455]), .B(p_input[37455]), .Z(n5657) );
  AND U8488 ( .A(n5659), .B(n5660), .Z(o[7454]) );
  AND U8489 ( .A(p_input[27454]), .B(p_input[17454]), .Z(n5660) );
  AND U8490 ( .A(p_input[7454]), .B(p_input[37454]), .Z(n5659) );
  AND U8491 ( .A(n5661), .B(n5662), .Z(o[7453]) );
  AND U8492 ( .A(p_input[27453]), .B(p_input[17453]), .Z(n5662) );
  AND U8493 ( .A(p_input[7453]), .B(p_input[37453]), .Z(n5661) );
  AND U8494 ( .A(n5663), .B(n5664), .Z(o[7452]) );
  AND U8495 ( .A(p_input[27452]), .B(p_input[17452]), .Z(n5664) );
  AND U8496 ( .A(p_input[7452]), .B(p_input[37452]), .Z(n5663) );
  AND U8497 ( .A(n5665), .B(n5666), .Z(o[7451]) );
  AND U8498 ( .A(p_input[27451]), .B(p_input[17451]), .Z(n5666) );
  AND U8499 ( .A(p_input[7451]), .B(p_input[37451]), .Z(n5665) );
  AND U8500 ( .A(n5667), .B(n5668), .Z(o[7450]) );
  AND U8501 ( .A(p_input[27450]), .B(p_input[17450]), .Z(n5668) );
  AND U8502 ( .A(p_input[7450]), .B(p_input[37450]), .Z(n5667) );
  AND U8503 ( .A(n5669), .B(n5670), .Z(o[744]) );
  AND U8504 ( .A(p_input[20744]), .B(p_input[10744]), .Z(n5670) );
  AND U8505 ( .A(p_input[744]), .B(p_input[30744]), .Z(n5669) );
  AND U8506 ( .A(n5671), .B(n5672), .Z(o[7449]) );
  AND U8507 ( .A(p_input[27449]), .B(p_input[17449]), .Z(n5672) );
  AND U8508 ( .A(p_input[7449]), .B(p_input[37449]), .Z(n5671) );
  AND U8509 ( .A(n5673), .B(n5674), .Z(o[7448]) );
  AND U8510 ( .A(p_input[27448]), .B(p_input[17448]), .Z(n5674) );
  AND U8511 ( .A(p_input[7448]), .B(p_input[37448]), .Z(n5673) );
  AND U8512 ( .A(n5675), .B(n5676), .Z(o[7447]) );
  AND U8513 ( .A(p_input[27447]), .B(p_input[17447]), .Z(n5676) );
  AND U8514 ( .A(p_input[7447]), .B(p_input[37447]), .Z(n5675) );
  AND U8515 ( .A(n5677), .B(n5678), .Z(o[7446]) );
  AND U8516 ( .A(p_input[27446]), .B(p_input[17446]), .Z(n5678) );
  AND U8517 ( .A(p_input[7446]), .B(p_input[37446]), .Z(n5677) );
  AND U8518 ( .A(n5679), .B(n5680), .Z(o[7445]) );
  AND U8519 ( .A(p_input[27445]), .B(p_input[17445]), .Z(n5680) );
  AND U8520 ( .A(p_input[7445]), .B(p_input[37445]), .Z(n5679) );
  AND U8521 ( .A(n5681), .B(n5682), .Z(o[7444]) );
  AND U8522 ( .A(p_input[27444]), .B(p_input[17444]), .Z(n5682) );
  AND U8523 ( .A(p_input[7444]), .B(p_input[37444]), .Z(n5681) );
  AND U8524 ( .A(n5683), .B(n5684), .Z(o[7443]) );
  AND U8525 ( .A(p_input[27443]), .B(p_input[17443]), .Z(n5684) );
  AND U8526 ( .A(p_input[7443]), .B(p_input[37443]), .Z(n5683) );
  AND U8527 ( .A(n5685), .B(n5686), .Z(o[7442]) );
  AND U8528 ( .A(p_input[27442]), .B(p_input[17442]), .Z(n5686) );
  AND U8529 ( .A(p_input[7442]), .B(p_input[37442]), .Z(n5685) );
  AND U8530 ( .A(n5687), .B(n5688), .Z(o[7441]) );
  AND U8531 ( .A(p_input[27441]), .B(p_input[17441]), .Z(n5688) );
  AND U8532 ( .A(p_input[7441]), .B(p_input[37441]), .Z(n5687) );
  AND U8533 ( .A(n5689), .B(n5690), .Z(o[7440]) );
  AND U8534 ( .A(p_input[27440]), .B(p_input[17440]), .Z(n5690) );
  AND U8535 ( .A(p_input[7440]), .B(p_input[37440]), .Z(n5689) );
  AND U8536 ( .A(n5691), .B(n5692), .Z(o[743]) );
  AND U8537 ( .A(p_input[20743]), .B(p_input[10743]), .Z(n5692) );
  AND U8538 ( .A(p_input[743]), .B(p_input[30743]), .Z(n5691) );
  AND U8539 ( .A(n5693), .B(n5694), .Z(o[7439]) );
  AND U8540 ( .A(p_input[27439]), .B(p_input[17439]), .Z(n5694) );
  AND U8541 ( .A(p_input[7439]), .B(p_input[37439]), .Z(n5693) );
  AND U8542 ( .A(n5695), .B(n5696), .Z(o[7438]) );
  AND U8543 ( .A(p_input[27438]), .B(p_input[17438]), .Z(n5696) );
  AND U8544 ( .A(p_input[7438]), .B(p_input[37438]), .Z(n5695) );
  AND U8545 ( .A(n5697), .B(n5698), .Z(o[7437]) );
  AND U8546 ( .A(p_input[27437]), .B(p_input[17437]), .Z(n5698) );
  AND U8547 ( .A(p_input[7437]), .B(p_input[37437]), .Z(n5697) );
  AND U8548 ( .A(n5699), .B(n5700), .Z(o[7436]) );
  AND U8549 ( .A(p_input[27436]), .B(p_input[17436]), .Z(n5700) );
  AND U8550 ( .A(p_input[7436]), .B(p_input[37436]), .Z(n5699) );
  AND U8551 ( .A(n5701), .B(n5702), .Z(o[7435]) );
  AND U8552 ( .A(p_input[27435]), .B(p_input[17435]), .Z(n5702) );
  AND U8553 ( .A(p_input[7435]), .B(p_input[37435]), .Z(n5701) );
  AND U8554 ( .A(n5703), .B(n5704), .Z(o[7434]) );
  AND U8555 ( .A(p_input[27434]), .B(p_input[17434]), .Z(n5704) );
  AND U8556 ( .A(p_input[7434]), .B(p_input[37434]), .Z(n5703) );
  AND U8557 ( .A(n5705), .B(n5706), .Z(o[7433]) );
  AND U8558 ( .A(p_input[27433]), .B(p_input[17433]), .Z(n5706) );
  AND U8559 ( .A(p_input[7433]), .B(p_input[37433]), .Z(n5705) );
  AND U8560 ( .A(n5707), .B(n5708), .Z(o[7432]) );
  AND U8561 ( .A(p_input[27432]), .B(p_input[17432]), .Z(n5708) );
  AND U8562 ( .A(p_input[7432]), .B(p_input[37432]), .Z(n5707) );
  AND U8563 ( .A(n5709), .B(n5710), .Z(o[7431]) );
  AND U8564 ( .A(p_input[27431]), .B(p_input[17431]), .Z(n5710) );
  AND U8565 ( .A(p_input[7431]), .B(p_input[37431]), .Z(n5709) );
  AND U8566 ( .A(n5711), .B(n5712), .Z(o[7430]) );
  AND U8567 ( .A(p_input[27430]), .B(p_input[17430]), .Z(n5712) );
  AND U8568 ( .A(p_input[7430]), .B(p_input[37430]), .Z(n5711) );
  AND U8569 ( .A(n5713), .B(n5714), .Z(o[742]) );
  AND U8570 ( .A(p_input[20742]), .B(p_input[10742]), .Z(n5714) );
  AND U8571 ( .A(p_input[742]), .B(p_input[30742]), .Z(n5713) );
  AND U8572 ( .A(n5715), .B(n5716), .Z(o[7429]) );
  AND U8573 ( .A(p_input[27429]), .B(p_input[17429]), .Z(n5716) );
  AND U8574 ( .A(p_input[7429]), .B(p_input[37429]), .Z(n5715) );
  AND U8575 ( .A(n5717), .B(n5718), .Z(o[7428]) );
  AND U8576 ( .A(p_input[27428]), .B(p_input[17428]), .Z(n5718) );
  AND U8577 ( .A(p_input[7428]), .B(p_input[37428]), .Z(n5717) );
  AND U8578 ( .A(n5719), .B(n5720), .Z(o[7427]) );
  AND U8579 ( .A(p_input[27427]), .B(p_input[17427]), .Z(n5720) );
  AND U8580 ( .A(p_input[7427]), .B(p_input[37427]), .Z(n5719) );
  AND U8581 ( .A(n5721), .B(n5722), .Z(o[7426]) );
  AND U8582 ( .A(p_input[27426]), .B(p_input[17426]), .Z(n5722) );
  AND U8583 ( .A(p_input[7426]), .B(p_input[37426]), .Z(n5721) );
  AND U8584 ( .A(n5723), .B(n5724), .Z(o[7425]) );
  AND U8585 ( .A(p_input[27425]), .B(p_input[17425]), .Z(n5724) );
  AND U8586 ( .A(p_input[7425]), .B(p_input[37425]), .Z(n5723) );
  AND U8587 ( .A(n5725), .B(n5726), .Z(o[7424]) );
  AND U8588 ( .A(p_input[27424]), .B(p_input[17424]), .Z(n5726) );
  AND U8589 ( .A(p_input[7424]), .B(p_input[37424]), .Z(n5725) );
  AND U8590 ( .A(n5727), .B(n5728), .Z(o[7423]) );
  AND U8591 ( .A(p_input[27423]), .B(p_input[17423]), .Z(n5728) );
  AND U8592 ( .A(p_input[7423]), .B(p_input[37423]), .Z(n5727) );
  AND U8593 ( .A(n5729), .B(n5730), .Z(o[7422]) );
  AND U8594 ( .A(p_input[27422]), .B(p_input[17422]), .Z(n5730) );
  AND U8595 ( .A(p_input[7422]), .B(p_input[37422]), .Z(n5729) );
  AND U8596 ( .A(n5731), .B(n5732), .Z(o[7421]) );
  AND U8597 ( .A(p_input[27421]), .B(p_input[17421]), .Z(n5732) );
  AND U8598 ( .A(p_input[7421]), .B(p_input[37421]), .Z(n5731) );
  AND U8599 ( .A(n5733), .B(n5734), .Z(o[7420]) );
  AND U8600 ( .A(p_input[27420]), .B(p_input[17420]), .Z(n5734) );
  AND U8601 ( .A(p_input[7420]), .B(p_input[37420]), .Z(n5733) );
  AND U8602 ( .A(n5735), .B(n5736), .Z(o[741]) );
  AND U8603 ( .A(p_input[20741]), .B(p_input[10741]), .Z(n5736) );
  AND U8604 ( .A(p_input[741]), .B(p_input[30741]), .Z(n5735) );
  AND U8605 ( .A(n5737), .B(n5738), .Z(o[7419]) );
  AND U8606 ( .A(p_input[27419]), .B(p_input[17419]), .Z(n5738) );
  AND U8607 ( .A(p_input[7419]), .B(p_input[37419]), .Z(n5737) );
  AND U8608 ( .A(n5739), .B(n5740), .Z(o[7418]) );
  AND U8609 ( .A(p_input[27418]), .B(p_input[17418]), .Z(n5740) );
  AND U8610 ( .A(p_input[7418]), .B(p_input[37418]), .Z(n5739) );
  AND U8611 ( .A(n5741), .B(n5742), .Z(o[7417]) );
  AND U8612 ( .A(p_input[27417]), .B(p_input[17417]), .Z(n5742) );
  AND U8613 ( .A(p_input[7417]), .B(p_input[37417]), .Z(n5741) );
  AND U8614 ( .A(n5743), .B(n5744), .Z(o[7416]) );
  AND U8615 ( .A(p_input[27416]), .B(p_input[17416]), .Z(n5744) );
  AND U8616 ( .A(p_input[7416]), .B(p_input[37416]), .Z(n5743) );
  AND U8617 ( .A(n5745), .B(n5746), .Z(o[7415]) );
  AND U8618 ( .A(p_input[27415]), .B(p_input[17415]), .Z(n5746) );
  AND U8619 ( .A(p_input[7415]), .B(p_input[37415]), .Z(n5745) );
  AND U8620 ( .A(n5747), .B(n5748), .Z(o[7414]) );
  AND U8621 ( .A(p_input[27414]), .B(p_input[17414]), .Z(n5748) );
  AND U8622 ( .A(p_input[7414]), .B(p_input[37414]), .Z(n5747) );
  AND U8623 ( .A(n5749), .B(n5750), .Z(o[7413]) );
  AND U8624 ( .A(p_input[27413]), .B(p_input[17413]), .Z(n5750) );
  AND U8625 ( .A(p_input[7413]), .B(p_input[37413]), .Z(n5749) );
  AND U8626 ( .A(n5751), .B(n5752), .Z(o[7412]) );
  AND U8627 ( .A(p_input[27412]), .B(p_input[17412]), .Z(n5752) );
  AND U8628 ( .A(p_input[7412]), .B(p_input[37412]), .Z(n5751) );
  AND U8629 ( .A(n5753), .B(n5754), .Z(o[7411]) );
  AND U8630 ( .A(p_input[27411]), .B(p_input[17411]), .Z(n5754) );
  AND U8631 ( .A(p_input[7411]), .B(p_input[37411]), .Z(n5753) );
  AND U8632 ( .A(n5755), .B(n5756), .Z(o[7410]) );
  AND U8633 ( .A(p_input[27410]), .B(p_input[17410]), .Z(n5756) );
  AND U8634 ( .A(p_input[7410]), .B(p_input[37410]), .Z(n5755) );
  AND U8635 ( .A(n5757), .B(n5758), .Z(o[740]) );
  AND U8636 ( .A(p_input[20740]), .B(p_input[10740]), .Z(n5758) );
  AND U8637 ( .A(p_input[740]), .B(p_input[30740]), .Z(n5757) );
  AND U8638 ( .A(n5759), .B(n5760), .Z(o[7409]) );
  AND U8639 ( .A(p_input[27409]), .B(p_input[17409]), .Z(n5760) );
  AND U8640 ( .A(p_input[7409]), .B(p_input[37409]), .Z(n5759) );
  AND U8641 ( .A(n5761), .B(n5762), .Z(o[7408]) );
  AND U8642 ( .A(p_input[27408]), .B(p_input[17408]), .Z(n5762) );
  AND U8643 ( .A(p_input[7408]), .B(p_input[37408]), .Z(n5761) );
  AND U8644 ( .A(n5763), .B(n5764), .Z(o[7407]) );
  AND U8645 ( .A(p_input[27407]), .B(p_input[17407]), .Z(n5764) );
  AND U8646 ( .A(p_input[7407]), .B(p_input[37407]), .Z(n5763) );
  AND U8647 ( .A(n5765), .B(n5766), .Z(o[7406]) );
  AND U8648 ( .A(p_input[27406]), .B(p_input[17406]), .Z(n5766) );
  AND U8649 ( .A(p_input[7406]), .B(p_input[37406]), .Z(n5765) );
  AND U8650 ( .A(n5767), .B(n5768), .Z(o[7405]) );
  AND U8651 ( .A(p_input[27405]), .B(p_input[17405]), .Z(n5768) );
  AND U8652 ( .A(p_input[7405]), .B(p_input[37405]), .Z(n5767) );
  AND U8653 ( .A(n5769), .B(n5770), .Z(o[7404]) );
  AND U8654 ( .A(p_input[27404]), .B(p_input[17404]), .Z(n5770) );
  AND U8655 ( .A(p_input[7404]), .B(p_input[37404]), .Z(n5769) );
  AND U8656 ( .A(n5771), .B(n5772), .Z(o[7403]) );
  AND U8657 ( .A(p_input[27403]), .B(p_input[17403]), .Z(n5772) );
  AND U8658 ( .A(p_input[7403]), .B(p_input[37403]), .Z(n5771) );
  AND U8659 ( .A(n5773), .B(n5774), .Z(o[7402]) );
  AND U8660 ( .A(p_input[27402]), .B(p_input[17402]), .Z(n5774) );
  AND U8661 ( .A(p_input[7402]), .B(p_input[37402]), .Z(n5773) );
  AND U8662 ( .A(n5775), .B(n5776), .Z(o[7401]) );
  AND U8663 ( .A(p_input[27401]), .B(p_input[17401]), .Z(n5776) );
  AND U8664 ( .A(p_input[7401]), .B(p_input[37401]), .Z(n5775) );
  AND U8665 ( .A(n5777), .B(n5778), .Z(o[7400]) );
  AND U8666 ( .A(p_input[27400]), .B(p_input[17400]), .Z(n5778) );
  AND U8667 ( .A(p_input[7400]), .B(p_input[37400]), .Z(n5777) );
  AND U8668 ( .A(n5779), .B(n5780), .Z(o[73]) );
  AND U8669 ( .A(p_input[20073]), .B(p_input[10073]), .Z(n5780) );
  AND U8670 ( .A(p_input[73]), .B(p_input[30073]), .Z(n5779) );
  AND U8671 ( .A(n5781), .B(n5782), .Z(o[739]) );
  AND U8672 ( .A(p_input[20739]), .B(p_input[10739]), .Z(n5782) );
  AND U8673 ( .A(p_input[739]), .B(p_input[30739]), .Z(n5781) );
  AND U8674 ( .A(n5783), .B(n5784), .Z(o[7399]) );
  AND U8675 ( .A(p_input[27399]), .B(p_input[17399]), .Z(n5784) );
  AND U8676 ( .A(p_input[7399]), .B(p_input[37399]), .Z(n5783) );
  AND U8677 ( .A(n5785), .B(n5786), .Z(o[7398]) );
  AND U8678 ( .A(p_input[27398]), .B(p_input[17398]), .Z(n5786) );
  AND U8679 ( .A(p_input[7398]), .B(p_input[37398]), .Z(n5785) );
  AND U8680 ( .A(n5787), .B(n5788), .Z(o[7397]) );
  AND U8681 ( .A(p_input[27397]), .B(p_input[17397]), .Z(n5788) );
  AND U8682 ( .A(p_input[7397]), .B(p_input[37397]), .Z(n5787) );
  AND U8683 ( .A(n5789), .B(n5790), .Z(o[7396]) );
  AND U8684 ( .A(p_input[27396]), .B(p_input[17396]), .Z(n5790) );
  AND U8685 ( .A(p_input[7396]), .B(p_input[37396]), .Z(n5789) );
  AND U8686 ( .A(n5791), .B(n5792), .Z(o[7395]) );
  AND U8687 ( .A(p_input[27395]), .B(p_input[17395]), .Z(n5792) );
  AND U8688 ( .A(p_input[7395]), .B(p_input[37395]), .Z(n5791) );
  AND U8689 ( .A(n5793), .B(n5794), .Z(o[7394]) );
  AND U8690 ( .A(p_input[27394]), .B(p_input[17394]), .Z(n5794) );
  AND U8691 ( .A(p_input[7394]), .B(p_input[37394]), .Z(n5793) );
  AND U8692 ( .A(n5795), .B(n5796), .Z(o[7393]) );
  AND U8693 ( .A(p_input[27393]), .B(p_input[17393]), .Z(n5796) );
  AND U8694 ( .A(p_input[7393]), .B(p_input[37393]), .Z(n5795) );
  AND U8695 ( .A(n5797), .B(n5798), .Z(o[7392]) );
  AND U8696 ( .A(p_input[27392]), .B(p_input[17392]), .Z(n5798) );
  AND U8697 ( .A(p_input[7392]), .B(p_input[37392]), .Z(n5797) );
  AND U8698 ( .A(n5799), .B(n5800), .Z(o[7391]) );
  AND U8699 ( .A(p_input[27391]), .B(p_input[17391]), .Z(n5800) );
  AND U8700 ( .A(p_input[7391]), .B(p_input[37391]), .Z(n5799) );
  AND U8701 ( .A(n5801), .B(n5802), .Z(o[7390]) );
  AND U8702 ( .A(p_input[27390]), .B(p_input[17390]), .Z(n5802) );
  AND U8703 ( .A(p_input[7390]), .B(p_input[37390]), .Z(n5801) );
  AND U8704 ( .A(n5803), .B(n5804), .Z(o[738]) );
  AND U8705 ( .A(p_input[20738]), .B(p_input[10738]), .Z(n5804) );
  AND U8706 ( .A(p_input[738]), .B(p_input[30738]), .Z(n5803) );
  AND U8707 ( .A(n5805), .B(n5806), .Z(o[7389]) );
  AND U8708 ( .A(p_input[27389]), .B(p_input[17389]), .Z(n5806) );
  AND U8709 ( .A(p_input[7389]), .B(p_input[37389]), .Z(n5805) );
  AND U8710 ( .A(n5807), .B(n5808), .Z(o[7388]) );
  AND U8711 ( .A(p_input[27388]), .B(p_input[17388]), .Z(n5808) );
  AND U8712 ( .A(p_input[7388]), .B(p_input[37388]), .Z(n5807) );
  AND U8713 ( .A(n5809), .B(n5810), .Z(o[7387]) );
  AND U8714 ( .A(p_input[27387]), .B(p_input[17387]), .Z(n5810) );
  AND U8715 ( .A(p_input[7387]), .B(p_input[37387]), .Z(n5809) );
  AND U8716 ( .A(n5811), .B(n5812), .Z(o[7386]) );
  AND U8717 ( .A(p_input[27386]), .B(p_input[17386]), .Z(n5812) );
  AND U8718 ( .A(p_input[7386]), .B(p_input[37386]), .Z(n5811) );
  AND U8719 ( .A(n5813), .B(n5814), .Z(o[7385]) );
  AND U8720 ( .A(p_input[27385]), .B(p_input[17385]), .Z(n5814) );
  AND U8721 ( .A(p_input[7385]), .B(p_input[37385]), .Z(n5813) );
  AND U8722 ( .A(n5815), .B(n5816), .Z(o[7384]) );
  AND U8723 ( .A(p_input[27384]), .B(p_input[17384]), .Z(n5816) );
  AND U8724 ( .A(p_input[7384]), .B(p_input[37384]), .Z(n5815) );
  AND U8725 ( .A(n5817), .B(n5818), .Z(o[7383]) );
  AND U8726 ( .A(p_input[27383]), .B(p_input[17383]), .Z(n5818) );
  AND U8727 ( .A(p_input[7383]), .B(p_input[37383]), .Z(n5817) );
  AND U8728 ( .A(n5819), .B(n5820), .Z(o[7382]) );
  AND U8729 ( .A(p_input[27382]), .B(p_input[17382]), .Z(n5820) );
  AND U8730 ( .A(p_input[7382]), .B(p_input[37382]), .Z(n5819) );
  AND U8731 ( .A(n5821), .B(n5822), .Z(o[7381]) );
  AND U8732 ( .A(p_input[27381]), .B(p_input[17381]), .Z(n5822) );
  AND U8733 ( .A(p_input[7381]), .B(p_input[37381]), .Z(n5821) );
  AND U8734 ( .A(n5823), .B(n5824), .Z(o[7380]) );
  AND U8735 ( .A(p_input[27380]), .B(p_input[17380]), .Z(n5824) );
  AND U8736 ( .A(p_input[7380]), .B(p_input[37380]), .Z(n5823) );
  AND U8737 ( .A(n5825), .B(n5826), .Z(o[737]) );
  AND U8738 ( .A(p_input[20737]), .B(p_input[10737]), .Z(n5826) );
  AND U8739 ( .A(p_input[737]), .B(p_input[30737]), .Z(n5825) );
  AND U8740 ( .A(n5827), .B(n5828), .Z(o[7379]) );
  AND U8741 ( .A(p_input[27379]), .B(p_input[17379]), .Z(n5828) );
  AND U8742 ( .A(p_input[7379]), .B(p_input[37379]), .Z(n5827) );
  AND U8743 ( .A(n5829), .B(n5830), .Z(o[7378]) );
  AND U8744 ( .A(p_input[27378]), .B(p_input[17378]), .Z(n5830) );
  AND U8745 ( .A(p_input[7378]), .B(p_input[37378]), .Z(n5829) );
  AND U8746 ( .A(n5831), .B(n5832), .Z(o[7377]) );
  AND U8747 ( .A(p_input[27377]), .B(p_input[17377]), .Z(n5832) );
  AND U8748 ( .A(p_input[7377]), .B(p_input[37377]), .Z(n5831) );
  AND U8749 ( .A(n5833), .B(n5834), .Z(o[7376]) );
  AND U8750 ( .A(p_input[27376]), .B(p_input[17376]), .Z(n5834) );
  AND U8751 ( .A(p_input[7376]), .B(p_input[37376]), .Z(n5833) );
  AND U8752 ( .A(n5835), .B(n5836), .Z(o[7375]) );
  AND U8753 ( .A(p_input[27375]), .B(p_input[17375]), .Z(n5836) );
  AND U8754 ( .A(p_input[7375]), .B(p_input[37375]), .Z(n5835) );
  AND U8755 ( .A(n5837), .B(n5838), .Z(o[7374]) );
  AND U8756 ( .A(p_input[27374]), .B(p_input[17374]), .Z(n5838) );
  AND U8757 ( .A(p_input[7374]), .B(p_input[37374]), .Z(n5837) );
  AND U8758 ( .A(n5839), .B(n5840), .Z(o[7373]) );
  AND U8759 ( .A(p_input[27373]), .B(p_input[17373]), .Z(n5840) );
  AND U8760 ( .A(p_input[7373]), .B(p_input[37373]), .Z(n5839) );
  AND U8761 ( .A(n5841), .B(n5842), .Z(o[7372]) );
  AND U8762 ( .A(p_input[27372]), .B(p_input[17372]), .Z(n5842) );
  AND U8763 ( .A(p_input[7372]), .B(p_input[37372]), .Z(n5841) );
  AND U8764 ( .A(n5843), .B(n5844), .Z(o[7371]) );
  AND U8765 ( .A(p_input[27371]), .B(p_input[17371]), .Z(n5844) );
  AND U8766 ( .A(p_input[7371]), .B(p_input[37371]), .Z(n5843) );
  AND U8767 ( .A(n5845), .B(n5846), .Z(o[7370]) );
  AND U8768 ( .A(p_input[27370]), .B(p_input[17370]), .Z(n5846) );
  AND U8769 ( .A(p_input[7370]), .B(p_input[37370]), .Z(n5845) );
  AND U8770 ( .A(n5847), .B(n5848), .Z(o[736]) );
  AND U8771 ( .A(p_input[20736]), .B(p_input[10736]), .Z(n5848) );
  AND U8772 ( .A(p_input[736]), .B(p_input[30736]), .Z(n5847) );
  AND U8773 ( .A(n5849), .B(n5850), .Z(o[7369]) );
  AND U8774 ( .A(p_input[27369]), .B(p_input[17369]), .Z(n5850) );
  AND U8775 ( .A(p_input[7369]), .B(p_input[37369]), .Z(n5849) );
  AND U8776 ( .A(n5851), .B(n5852), .Z(o[7368]) );
  AND U8777 ( .A(p_input[27368]), .B(p_input[17368]), .Z(n5852) );
  AND U8778 ( .A(p_input[7368]), .B(p_input[37368]), .Z(n5851) );
  AND U8779 ( .A(n5853), .B(n5854), .Z(o[7367]) );
  AND U8780 ( .A(p_input[27367]), .B(p_input[17367]), .Z(n5854) );
  AND U8781 ( .A(p_input[7367]), .B(p_input[37367]), .Z(n5853) );
  AND U8782 ( .A(n5855), .B(n5856), .Z(o[7366]) );
  AND U8783 ( .A(p_input[27366]), .B(p_input[17366]), .Z(n5856) );
  AND U8784 ( .A(p_input[7366]), .B(p_input[37366]), .Z(n5855) );
  AND U8785 ( .A(n5857), .B(n5858), .Z(o[7365]) );
  AND U8786 ( .A(p_input[27365]), .B(p_input[17365]), .Z(n5858) );
  AND U8787 ( .A(p_input[7365]), .B(p_input[37365]), .Z(n5857) );
  AND U8788 ( .A(n5859), .B(n5860), .Z(o[7364]) );
  AND U8789 ( .A(p_input[27364]), .B(p_input[17364]), .Z(n5860) );
  AND U8790 ( .A(p_input[7364]), .B(p_input[37364]), .Z(n5859) );
  AND U8791 ( .A(n5861), .B(n5862), .Z(o[7363]) );
  AND U8792 ( .A(p_input[27363]), .B(p_input[17363]), .Z(n5862) );
  AND U8793 ( .A(p_input[7363]), .B(p_input[37363]), .Z(n5861) );
  AND U8794 ( .A(n5863), .B(n5864), .Z(o[7362]) );
  AND U8795 ( .A(p_input[27362]), .B(p_input[17362]), .Z(n5864) );
  AND U8796 ( .A(p_input[7362]), .B(p_input[37362]), .Z(n5863) );
  AND U8797 ( .A(n5865), .B(n5866), .Z(o[7361]) );
  AND U8798 ( .A(p_input[27361]), .B(p_input[17361]), .Z(n5866) );
  AND U8799 ( .A(p_input[7361]), .B(p_input[37361]), .Z(n5865) );
  AND U8800 ( .A(n5867), .B(n5868), .Z(o[7360]) );
  AND U8801 ( .A(p_input[27360]), .B(p_input[17360]), .Z(n5868) );
  AND U8802 ( .A(p_input[7360]), .B(p_input[37360]), .Z(n5867) );
  AND U8803 ( .A(n5869), .B(n5870), .Z(o[735]) );
  AND U8804 ( .A(p_input[20735]), .B(p_input[10735]), .Z(n5870) );
  AND U8805 ( .A(p_input[735]), .B(p_input[30735]), .Z(n5869) );
  AND U8806 ( .A(n5871), .B(n5872), .Z(o[7359]) );
  AND U8807 ( .A(p_input[27359]), .B(p_input[17359]), .Z(n5872) );
  AND U8808 ( .A(p_input[7359]), .B(p_input[37359]), .Z(n5871) );
  AND U8809 ( .A(n5873), .B(n5874), .Z(o[7358]) );
  AND U8810 ( .A(p_input[27358]), .B(p_input[17358]), .Z(n5874) );
  AND U8811 ( .A(p_input[7358]), .B(p_input[37358]), .Z(n5873) );
  AND U8812 ( .A(n5875), .B(n5876), .Z(o[7357]) );
  AND U8813 ( .A(p_input[27357]), .B(p_input[17357]), .Z(n5876) );
  AND U8814 ( .A(p_input[7357]), .B(p_input[37357]), .Z(n5875) );
  AND U8815 ( .A(n5877), .B(n5878), .Z(o[7356]) );
  AND U8816 ( .A(p_input[27356]), .B(p_input[17356]), .Z(n5878) );
  AND U8817 ( .A(p_input[7356]), .B(p_input[37356]), .Z(n5877) );
  AND U8818 ( .A(n5879), .B(n5880), .Z(o[7355]) );
  AND U8819 ( .A(p_input[27355]), .B(p_input[17355]), .Z(n5880) );
  AND U8820 ( .A(p_input[7355]), .B(p_input[37355]), .Z(n5879) );
  AND U8821 ( .A(n5881), .B(n5882), .Z(o[7354]) );
  AND U8822 ( .A(p_input[27354]), .B(p_input[17354]), .Z(n5882) );
  AND U8823 ( .A(p_input[7354]), .B(p_input[37354]), .Z(n5881) );
  AND U8824 ( .A(n5883), .B(n5884), .Z(o[7353]) );
  AND U8825 ( .A(p_input[27353]), .B(p_input[17353]), .Z(n5884) );
  AND U8826 ( .A(p_input[7353]), .B(p_input[37353]), .Z(n5883) );
  AND U8827 ( .A(n5885), .B(n5886), .Z(o[7352]) );
  AND U8828 ( .A(p_input[27352]), .B(p_input[17352]), .Z(n5886) );
  AND U8829 ( .A(p_input[7352]), .B(p_input[37352]), .Z(n5885) );
  AND U8830 ( .A(n5887), .B(n5888), .Z(o[7351]) );
  AND U8831 ( .A(p_input[27351]), .B(p_input[17351]), .Z(n5888) );
  AND U8832 ( .A(p_input[7351]), .B(p_input[37351]), .Z(n5887) );
  AND U8833 ( .A(n5889), .B(n5890), .Z(o[7350]) );
  AND U8834 ( .A(p_input[27350]), .B(p_input[17350]), .Z(n5890) );
  AND U8835 ( .A(p_input[7350]), .B(p_input[37350]), .Z(n5889) );
  AND U8836 ( .A(n5891), .B(n5892), .Z(o[734]) );
  AND U8837 ( .A(p_input[20734]), .B(p_input[10734]), .Z(n5892) );
  AND U8838 ( .A(p_input[734]), .B(p_input[30734]), .Z(n5891) );
  AND U8839 ( .A(n5893), .B(n5894), .Z(o[7349]) );
  AND U8840 ( .A(p_input[27349]), .B(p_input[17349]), .Z(n5894) );
  AND U8841 ( .A(p_input[7349]), .B(p_input[37349]), .Z(n5893) );
  AND U8842 ( .A(n5895), .B(n5896), .Z(o[7348]) );
  AND U8843 ( .A(p_input[27348]), .B(p_input[17348]), .Z(n5896) );
  AND U8844 ( .A(p_input[7348]), .B(p_input[37348]), .Z(n5895) );
  AND U8845 ( .A(n5897), .B(n5898), .Z(o[7347]) );
  AND U8846 ( .A(p_input[27347]), .B(p_input[17347]), .Z(n5898) );
  AND U8847 ( .A(p_input[7347]), .B(p_input[37347]), .Z(n5897) );
  AND U8848 ( .A(n5899), .B(n5900), .Z(o[7346]) );
  AND U8849 ( .A(p_input[27346]), .B(p_input[17346]), .Z(n5900) );
  AND U8850 ( .A(p_input[7346]), .B(p_input[37346]), .Z(n5899) );
  AND U8851 ( .A(n5901), .B(n5902), .Z(o[7345]) );
  AND U8852 ( .A(p_input[27345]), .B(p_input[17345]), .Z(n5902) );
  AND U8853 ( .A(p_input[7345]), .B(p_input[37345]), .Z(n5901) );
  AND U8854 ( .A(n5903), .B(n5904), .Z(o[7344]) );
  AND U8855 ( .A(p_input[27344]), .B(p_input[17344]), .Z(n5904) );
  AND U8856 ( .A(p_input[7344]), .B(p_input[37344]), .Z(n5903) );
  AND U8857 ( .A(n5905), .B(n5906), .Z(o[7343]) );
  AND U8858 ( .A(p_input[27343]), .B(p_input[17343]), .Z(n5906) );
  AND U8859 ( .A(p_input[7343]), .B(p_input[37343]), .Z(n5905) );
  AND U8860 ( .A(n5907), .B(n5908), .Z(o[7342]) );
  AND U8861 ( .A(p_input[27342]), .B(p_input[17342]), .Z(n5908) );
  AND U8862 ( .A(p_input[7342]), .B(p_input[37342]), .Z(n5907) );
  AND U8863 ( .A(n5909), .B(n5910), .Z(o[7341]) );
  AND U8864 ( .A(p_input[27341]), .B(p_input[17341]), .Z(n5910) );
  AND U8865 ( .A(p_input[7341]), .B(p_input[37341]), .Z(n5909) );
  AND U8866 ( .A(n5911), .B(n5912), .Z(o[7340]) );
  AND U8867 ( .A(p_input[27340]), .B(p_input[17340]), .Z(n5912) );
  AND U8868 ( .A(p_input[7340]), .B(p_input[37340]), .Z(n5911) );
  AND U8869 ( .A(n5913), .B(n5914), .Z(o[733]) );
  AND U8870 ( .A(p_input[20733]), .B(p_input[10733]), .Z(n5914) );
  AND U8871 ( .A(p_input[733]), .B(p_input[30733]), .Z(n5913) );
  AND U8872 ( .A(n5915), .B(n5916), .Z(o[7339]) );
  AND U8873 ( .A(p_input[27339]), .B(p_input[17339]), .Z(n5916) );
  AND U8874 ( .A(p_input[7339]), .B(p_input[37339]), .Z(n5915) );
  AND U8875 ( .A(n5917), .B(n5918), .Z(o[7338]) );
  AND U8876 ( .A(p_input[27338]), .B(p_input[17338]), .Z(n5918) );
  AND U8877 ( .A(p_input[7338]), .B(p_input[37338]), .Z(n5917) );
  AND U8878 ( .A(n5919), .B(n5920), .Z(o[7337]) );
  AND U8879 ( .A(p_input[27337]), .B(p_input[17337]), .Z(n5920) );
  AND U8880 ( .A(p_input[7337]), .B(p_input[37337]), .Z(n5919) );
  AND U8881 ( .A(n5921), .B(n5922), .Z(o[7336]) );
  AND U8882 ( .A(p_input[27336]), .B(p_input[17336]), .Z(n5922) );
  AND U8883 ( .A(p_input[7336]), .B(p_input[37336]), .Z(n5921) );
  AND U8884 ( .A(n5923), .B(n5924), .Z(o[7335]) );
  AND U8885 ( .A(p_input[27335]), .B(p_input[17335]), .Z(n5924) );
  AND U8886 ( .A(p_input[7335]), .B(p_input[37335]), .Z(n5923) );
  AND U8887 ( .A(n5925), .B(n5926), .Z(o[7334]) );
  AND U8888 ( .A(p_input[27334]), .B(p_input[17334]), .Z(n5926) );
  AND U8889 ( .A(p_input[7334]), .B(p_input[37334]), .Z(n5925) );
  AND U8890 ( .A(n5927), .B(n5928), .Z(o[7333]) );
  AND U8891 ( .A(p_input[27333]), .B(p_input[17333]), .Z(n5928) );
  AND U8892 ( .A(p_input[7333]), .B(p_input[37333]), .Z(n5927) );
  AND U8893 ( .A(n5929), .B(n5930), .Z(o[7332]) );
  AND U8894 ( .A(p_input[27332]), .B(p_input[17332]), .Z(n5930) );
  AND U8895 ( .A(p_input[7332]), .B(p_input[37332]), .Z(n5929) );
  AND U8896 ( .A(n5931), .B(n5932), .Z(o[7331]) );
  AND U8897 ( .A(p_input[27331]), .B(p_input[17331]), .Z(n5932) );
  AND U8898 ( .A(p_input[7331]), .B(p_input[37331]), .Z(n5931) );
  AND U8899 ( .A(n5933), .B(n5934), .Z(o[7330]) );
  AND U8900 ( .A(p_input[27330]), .B(p_input[17330]), .Z(n5934) );
  AND U8901 ( .A(p_input[7330]), .B(p_input[37330]), .Z(n5933) );
  AND U8902 ( .A(n5935), .B(n5936), .Z(o[732]) );
  AND U8903 ( .A(p_input[20732]), .B(p_input[10732]), .Z(n5936) );
  AND U8904 ( .A(p_input[732]), .B(p_input[30732]), .Z(n5935) );
  AND U8905 ( .A(n5937), .B(n5938), .Z(o[7329]) );
  AND U8906 ( .A(p_input[27329]), .B(p_input[17329]), .Z(n5938) );
  AND U8907 ( .A(p_input[7329]), .B(p_input[37329]), .Z(n5937) );
  AND U8908 ( .A(n5939), .B(n5940), .Z(o[7328]) );
  AND U8909 ( .A(p_input[27328]), .B(p_input[17328]), .Z(n5940) );
  AND U8910 ( .A(p_input[7328]), .B(p_input[37328]), .Z(n5939) );
  AND U8911 ( .A(n5941), .B(n5942), .Z(o[7327]) );
  AND U8912 ( .A(p_input[27327]), .B(p_input[17327]), .Z(n5942) );
  AND U8913 ( .A(p_input[7327]), .B(p_input[37327]), .Z(n5941) );
  AND U8914 ( .A(n5943), .B(n5944), .Z(o[7326]) );
  AND U8915 ( .A(p_input[27326]), .B(p_input[17326]), .Z(n5944) );
  AND U8916 ( .A(p_input[7326]), .B(p_input[37326]), .Z(n5943) );
  AND U8917 ( .A(n5945), .B(n5946), .Z(o[7325]) );
  AND U8918 ( .A(p_input[27325]), .B(p_input[17325]), .Z(n5946) );
  AND U8919 ( .A(p_input[7325]), .B(p_input[37325]), .Z(n5945) );
  AND U8920 ( .A(n5947), .B(n5948), .Z(o[7324]) );
  AND U8921 ( .A(p_input[27324]), .B(p_input[17324]), .Z(n5948) );
  AND U8922 ( .A(p_input[7324]), .B(p_input[37324]), .Z(n5947) );
  AND U8923 ( .A(n5949), .B(n5950), .Z(o[7323]) );
  AND U8924 ( .A(p_input[27323]), .B(p_input[17323]), .Z(n5950) );
  AND U8925 ( .A(p_input[7323]), .B(p_input[37323]), .Z(n5949) );
  AND U8926 ( .A(n5951), .B(n5952), .Z(o[7322]) );
  AND U8927 ( .A(p_input[27322]), .B(p_input[17322]), .Z(n5952) );
  AND U8928 ( .A(p_input[7322]), .B(p_input[37322]), .Z(n5951) );
  AND U8929 ( .A(n5953), .B(n5954), .Z(o[7321]) );
  AND U8930 ( .A(p_input[27321]), .B(p_input[17321]), .Z(n5954) );
  AND U8931 ( .A(p_input[7321]), .B(p_input[37321]), .Z(n5953) );
  AND U8932 ( .A(n5955), .B(n5956), .Z(o[7320]) );
  AND U8933 ( .A(p_input[27320]), .B(p_input[17320]), .Z(n5956) );
  AND U8934 ( .A(p_input[7320]), .B(p_input[37320]), .Z(n5955) );
  AND U8935 ( .A(n5957), .B(n5958), .Z(o[731]) );
  AND U8936 ( .A(p_input[20731]), .B(p_input[10731]), .Z(n5958) );
  AND U8937 ( .A(p_input[731]), .B(p_input[30731]), .Z(n5957) );
  AND U8938 ( .A(n5959), .B(n5960), .Z(o[7319]) );
  AND U8939 ( .A(p_input[27319]), .B(p_input[17319]), .Z(n5960) );
  AND U8940 ( .A(p_input[7319]), .B(p_input[37319]), .Z(n5959) );
  AND U8941 ( .A(n5961), .B(n5962), .Z(o[7318]) );
  AND U8942 ( .A(p_input[27318]), .B(p_input[17318]), .Z(n5962) );
  AND U8943 ( .A(p_input[7318]), .B(p_input[37318]), .Z(n5961) );
  AND U8944 ( .A(n5963), .B(n5964), .Z(o[7317]) );
  AND U8945 ( .A(p_input[27317]), .B(p_input[17317]), .Z(n5964) );
  AND U8946 ( .A(p_input[7317]), .B(p_input[37317]), .Z(n5963) );
  AND U8947 ( .A(n5965), .B(n5966), .Z(o[7316]) );
  AND U8948 ( .A(p_input[27316]), .B(p_input[17316]), .Z(n5966) );
  AND U8949 ( .A(p_input[7316]), .B(p_input[37316]), .Z(n5965) );
  AND U8950 ( .A(n5967), .B(n5968), .Z(o[7315]) );
  AND U8951 ( .A(p_input[27315]), .B(p_input[17315]), .Z(n5968) );
  AND U8952 ( .A(p_input[7315]), .B(p_input[37315]), .Z(n5967) );
  AND U8953 ( .A(n5969), .B(n5970), .Z(o[7314]) );
  AND U8954 ( .A(p_input[27314]), .B(p_input[17314]), .Z(n5970) );
  AND U8955 ( .A(p_input[7314]), .B(p_input[37314]), .Z(n5969) );
  AND U8956 ( .A(n5971), .B(n5972), .Z(o[7313]) );
  AND U8957 ( .A(p_input[27313]), .B(p_input[17313]), .Z(n5972) );
  AND U8958 ( .A(p_input[7313]), .B(p_input[37313]), .Z(n5971) );
  AND U8959 ( .A(n5973), .B(n5974), .Z(o[7312]) );
  AND U8960 ( .A(p_input[27312]), .B(p_input[17312]), .Z(n5974) );
  AND U8961 ( .A(p_input[7312]), .B(p_input[37312]), .Z(n5973) );
  AND U8962 ( .A(n5975), .B(n5976), .Z(o[7311]) );
  AND U8963 ( .A(p_input[27311]), .B(p_input[17311]), .Z(n5976) );
  AND U8964 ( .A(p_input[7311]), .B(p_input[37311]), .Z(n5975) );
  AND U8965 ( .A(n5977), .B(n5978), .Z(o[7310]) );
  AND U8966 ( .A(p_input[27310]), .B(p_input[17310]), .Z(n5978) );
  AND U8967 ( .A(p_input[7310]), .B(p_input[37310]), .Z(n5977) );
  AND U8968 ( .A(n5979), .B(n5980), .Z(o[730]) );
  AND U8969 ( .A(p_input[20730]), .B(p_input[10730]), .Z(n5980) );
  AND U8970 ( .A(p_input[730]), .B(p_input[30730]), .Z(n5979) );
  AND U8971 ( .A(n5981), .B(n5982), .Z(o[7309]) );
  AND U8972 ( .A(p_input[27309]), .B(p_input[17309]), .Z(n5982) );
  AND U8973 ( .A(p_input[7309]), .B(p_input[37309]), .Z(n5981) );
  AND U8974 ( .A(n5983), .B(n5984), .Z(o[7308]) );
  AND U8975 ( .A(p_input[27308]), .B(p_input[17308]), .Z(n5984) );
  AND U8976 ( .A(p_input[7308]), .B(p_input[37308]), .Z(n5983) );
  AND U8977 ( .A(n5985), .B(n5986), .Z(o[7307]) );
  AND U8978 ( .A(p_input[27307]), .B(p_input[17307]), .Z(n5986) );
  AND U8979 ( .A(p_input[7307]), .B(p_input[37307]), .Z(n5985) );
  AND U8980 ( .A(n5987), .B(n5988), .Z(o[7306]) );
  AND U8981 ( .A(p_input[27306]), .B(p_input[17306]), .Z(n5988) );
  AND U8982 ( .A(p_input[7306]), .B(p_input[37306]), .Z(n5987) );
  AND U8983 ( .A(n5989), .B(n5990), .Z(o[7305]) );
  AND U8984 ( .A(p_input[27305]), .B(p_input[17305]), .Z(n5990) );
  AND U8985 ( .A(p_input[7305]), .B(p_input[37305]), .Z(n5989) );
  AND U8986 ( .A(n5991), .B(n5992), .Z(o[7304]) );
  AND U8987 ( .A(p_input[27304]), .B(p_input[17304]), .Z(n5992) );
  AND U8988 ( .A(p_input[7304]), .B(p_input[37304]), .Z(n5991) );
  AND U8989 ( .A(n5993), .B(n5994), .Z(o[7303]) );
  AND U8990 ( .A(p_input[27303]), .B(p_input[17303]), .Z(n5994) );
  AND U8991 ( .A(p_input[7303]), .B(p_input[37303]), .Z(n5993) );
  AND U8992 ( .A(n5995), .B(n5996), .Z(o[7302]) );
  AND U8993 ( .A(p_input[27302]), .B(p_input[17302]), .Z(n5996) );
  AND U8994 ( .A(p_input[7302]), .B(p_input[37302]), .Z(n5995) );
  AND U8995 ( .A(n5997), .B(n5998), .Z(o[7301]) );
  AND U8996 ( .A(p_input[27301]), .B(p_input[17301]), .Z(n5998) );
  AND U8997 ( .A(p_input[7301]), .B(p_input[37301]), .Z(n5997) );
  AND U8998 ( .A(n5999), .B(n6000), .Z(o[7300]) );
  AND U8999 ( .A(p_input[27300]), .B(p_input[17300]), .Z(n6000) );
  AND U9000 ( .A(p_input[7300]), .B(p_input[37300]), .Z(n5999) );
  AND U9001 ( .A(n6001), .B(n6002), .Z(o[72]) );
  AND U9002 ( .A(p_input[20072]), .B(p_input[10072]), .Z(n6002) );
  AND U9003 ( .A(p_input[72]), .B(p_input[30072]), .Z(n6001) );
  AND U9004 ( .A(n6003), .B(n6004), .Z(o[729]) );
  AND U9005 ( .A(p_input[20729]), .B(p_input[10729]), .Z(n6004) );
  AND U9006 ( .A(p_input[729]), .B(p_input[30729]), .Z(n6003) );
  AND U9007 ( .A(n6005), .B(n6006), .Z(o[7299]) );
  AND U9008 ( .A(p_input[27299]), .B(p_input[17299]), .Z(n6006) );
  AND U9009 ( .A(p_input[7299]), .B(p_input[37299]), .Z(n6005) );
  AND U9010 ( .A(n6007), .B(n6008), .Z(o[7298]) );
  AND U9011 ( .A(p_input[27298]), .B(p_input[17298]), .Z(n6008) );
  AND U9012 ( .A(p_input[7298]), .B(p_input[37298]), .Z(n6007) );
  AND U9013 ( .A(n6009), .B(n6010), .Z(o[7297]) );
  AND U9014 ( .A(p_input[27297]), .B(p_input[17297]), .Z(n6010) );
  AND U9015 ( .A(p_input[7297]), .B(p_input[37297]), .Z(n6009) );
  AND U9016 ( .A(n6011), .B(n6012), .Z(o[7296]) );
  AND U9017 ( .A(p_input[27296]), .B(p_input[17296]), .Z(n6012) );
  AND U9018 ( .A(p_input[7296]), .B(p_input[37296]), .Z(n6011) );
  AND U9019 ( .A(n6013), .B(n6014), .Z(o[7295]) );
  AND U9020 ( .A(p_input[27295]), .B(p_input[17295]), .Z(n6014) );
  AND U9021 ( .A(p_input[7295]), .B(p_input[37295]), .Z(n6013) );
  AND U9022 ( .A(n6015), .B(n6016), .Z(o[7294]) );
  AND U9023 ( .A(p_input[27294]), .B(p_input[17294]), .Z(n6016) );
  AND U9024 ( .A(p_input[7294]), .B(p_input[37294]), .Z(n6015) );
  AND U9025 ( .A(n6017), .B(n6018), .Z(o[7293]) );
  AND U9026 ( .A(p_input[27293]), .B(p_input[17293]), .Z(n6018) );
  AND U9027 ( .A(p_input[7293]), .B(p_input[37293]), .Z(n6017) );
  AND U9028 ( .A(n6019), .B(n6020), .Z(o[7292]) );
  AND U9029 ( .A(p_input[27292]), .B(p_input[17292]), .Z(n6020) );
  AND U9030 ( .A(p_input[7292]), .B(p_input[37292]), .Z(n6019) );
  AND U9031 ( .A(n6021), .B(n6022), .Z(o[7291]) );
  AND U9032 ( .A(p_input[27291]), .B(p_input[17291]), .Z(n6022) );
  AND U9033 ( .A(p_input[7291]), .B(p_input[37291]), .Z(n6021) );
  AND U9034 ( .A(n6023), .B(n6024), .Z(o[7290]) );
  AND U9035 ( .A(p_input[27290]), .B(p_input[17290]), .Z(n6024) );
  AND U9036 ( .A(p_input[7290]), .B(p_input[37290]), .Z(n6023) );
  AND U9037 ( .A(n6025), .B(n6026), .Z(o[728]) );
  AND U9038 ( .A(p_input[20728]), .B(p_input[10728]), .Z(n6026) );
  AND U9039 ( .A(p_input[728]), .B(p_input[30728]), .Z(n6025) );
  AND U9040 ( .A(n6027), .B(n6028), .Z(o[7289]) );
  AND U9041 ( .A(p_input[27289]), .B(p_input[17289]), .Z(n6028) );
  AND U9042 ( .A(p_input[7289]), .B(p_input[37289]), .Z(n6027) );
  AND U9043 ( .A(n6029), .B(n6030), .Z(o[7288]) );
  AND U9044 ( .A(p_input[27288]), .B(p_input[17288]), .Z(n6030) );
  AND U9045 ( .A(p_input[7288]), .B(p_input[37288]), .Z(n6029) );
  AND U9046 ( .A(n6031), .B(n6032), .Z(o[7287]) );
  AND U9047 ( .A(p_input[27287]), .B(p_input[17287]), .Z(n6032) );
  AND U9048 ( .A(p_input[7287]), .B(p_input[37287]), .Z(n6031) );
  AND U9049 ( .A(n6033), .B(n6034), .Z(o[7286]) );
  AND U9050 ( .A(p_input[27286]), .B(p_input[17286]), .Z(n6034) );
  AND U9051 ( .A(p_input[7286]), .B(p_input[37286]), .Z(n6033) );
  AND U9052 ( .A(n6035), .B(n6036), .Z(o[7285]) );
  AND U9053 ( .A(p_input[27285]), .B(p_input[17285]), .Z(n6036) );
  AND U9054 ( .A(p_input[7285]), .B(p_input[37285]), .Z(n6035) );
  AND U9055 ( .A(n6037), .B(n6038), .Z(o[7284]) );
  AND U9056 ( .A(p_input[27284]), .B(p_input[17284]), .Z(n6038) );
  AND U9057 ( .A(p_input[7284]), .B(p_input[37284]), .Z(n6037) );
  AND U9058 ( .A(n6039), .B(n6040), .Z(o[7283]) );
  AND U9059 ( .A(p_input[27283]), .B(p_input[17283]), .Z(n6040) );
  AND U9060 ( .A(p_input[7283]), .B(p_input[37283]), .Z(n6039) );
  AND U9061 ( .A(n6041), .B(n6042), .Z(o[7282]) );
  AND U9062 ( .A(p_input[27282]), .B(p_input[17282]), .Z(n6042) );
  AND U9063 ( .A(p_input[7282]), .B(p_input[37282]), .Z(n6041) );
  AND U9064 ( .A(n6043), .B(n6044), .Z(o[7281]) );
  AND U9065 ( .A(p_input[27281]), .B(p_input[17281]), .Z(n6044) );
  AND U9066 ( .A(p_input[7281]), .B(p_input[37281]), .Z(n6043) );
  AND U9067 ( .A(n6045), .B(n6046), .Z(o[7280]) );
  AND U9068 ( .A(p_input[27280]), .B(p_input[17280]), .Z(n6046) );
  AND U9069 ( .A(p_input[7280]), .B(p_input[37280]), .Z(n6045) );
  AND U9070 ( .A(n6047), .B(n6048), .Z(o[727]) );
  AND U9071 ( .A(p_input[20727]), .B(p_input[10727]), .Z(n6048) );
  AND U9072 ( .A(p_input[727]), .B(p_input[30727]), .Z(n6047) );
  AND U9073 ( .A(n6049), .B(n6050), .Z(o[7279]) );
  AND U9074 ( .A(p_input[27279]), .B(p_input[17279]), .Z(n6050) );
  AND U9075 ( .A(p_input[7279]), .B(p_input[37279]), .Z(n6049) );
  AND U9076 ( .A(n6051), .B(n6052), .Z(o[7278]) );
  AND U9077 ( .A(p_input[27278]), .B(p_input[17278]), .Z(n6052) );
  AND U9078 ( .A(p_input[7278]), .B(p_input[37278]), .Z(n6051) );
  AND U9079 ( .A(n6053), .B(n6054), .Z(o[7277]) );
  AND U9080 ( .A(p_input[27277]), .B(p_input[17277]), .Z(n6054) );
  AND U9081 ( .A(p_input[7277]), .B(p_input[37277]), .Z(n6053) );
  AND U9082 ( .A(n6055), .B(n6056), .Z(o[7276]) );
  AND U9083 ( .A(p_input[27276]), .B(p_input[17276]), .Z(n6056) );
  AND U9084 ( .A(p_input[7276]), .B(p_input[37276]), .Z(n6055) );
  AND U9085 ( .A(n6057), .B(n6058), .Z(o[7275]) );
  AND U9086 ( .A(p_input[27275]), .B(p_input[17275]), .Z(n6058) );
  AND U9087 ( .A(p_input[7275]), .B(p_input[37275]), .Z(n6057) );
  AND U9088 ( .A(n6059), .B(n6060), .Z(o[7274]) );
  AND U9089 ( .A(p_input[27274]), .B(p_input[17274]), .Z(n6060) );
  AND U9090 ( .A(p_input[7274]), .B(p_input[37274]), .Z(n6059) );
  AND U9091 ( .A(n6061), .B(n6062), .Z(o[7273]) );
  AND U9092 ( .A(p_input[27273]), .B(p_input[17273]), .Z(n6062) );
  AND U9093 ( .A(p_input[7273]), .B(p_input[37273]), .Z(n6061) );
  AND U9094 ( .A(n6063), .B(n6064), .Z(o[7272]) );
  AND U9095 ( .A(p_input[27272]), .B(p_input[17272]), .Z(n6064) );
  AND U9096 ( .A(p_input[7272]), .B(p_input[37272]), .Z(n6063) );
  AND U9097 ( .A(n6065), .B(n6066), .Z(o[7271]) );
  AND U9098 ( .A(p_input[27271]), .B(p_input[17271]), .Z(n6066) );
  AND U9099 ( .A(p_input[7271]), .B(p_input[37271]), .Z(n6065) );
  AND U9100 ( .A(n6067), .B(n6068), .Z(o[7270]) );
  AND U9101 ( .A(p_input[27270]), .B(p_input[17270]), .Z(n6068) );
  AND U9102 ( .A(p_input[7270]), .B(p_input[37270]), .Z(n6067) );
  AND U9103 ( .A(n6069), .B(n6070), .Z(o[726]) );
  AND U9104 ( .A(p_input[20726]), .B(p_input[10726]), .Z(n6070) );
  AND U9105 ( .A(p_input[726]), .B(p_input[30726]), .Z(n6069) );
  AND U9106 ( .A(n6071), .B(n6072), .Z(o[7269]) );
  AND U9107 ( .A(p_input[27269]), .B(p_input[17269]), .Z(n6072) );
  AND U9108 ( .A(p_input[7269]), .B(p_input[37269]), .Z(n6071) );
  AND U9109 ( .A(n6073), .B(n6074), .Z(o[7268]) );
  AND U9110 ( .A(p_input[27268]), .B(p_input[17268]), .Z(n6074) );
  AND U9111 ( .A(p_input[7268]), .B(p_input[37268]), .Z(n6073) );
  AND U9112 ( .A(n6075), .B(n6076), .Z(o[7267]) );
  AND U9113 ( .A(p_input[27267]), .B(p_input[17267]), .Z(n6076) );
  AND U9114 ( .A(p_input[7267]), .B(p_input[37267]), .Z(n6075) );
  AND U9115 ( .A(n6077), .B(n6078), .Z(o[7266]) );
  AND U9116 ( .A(p_input[27266]), .B(p_input[17266]), .Z(n6078) );
  AND U9117 ( .A(p_input[7266]), .B(p_input[37266]), .Z(n6077) );
  AND U9118 ( .A(n6079), .B(n6080), .Z(o[7265]) );
  AND U9119 ( .A(p_input[27265]), .B(p_input[17265]), .Z(n6080) );
  AND U9120 ( .A(p_input[7265]), .B(p_input[37265]), .Z(n6079) );
  AND U9121 ( .A(n6081), .B(n6082), .Z(o[7264]) );
  AND U9122 ( .A(p_input[27264]), .B(p_input[17264]), .Z(n6082) );
  AND U9123 ( .A(p_input[7264]), .B(p_input[37264]), .Z(n6081) );
  AND U9124 ( .A(n6083), .B(n6084), .Z(o[7263]) );
  AND U9125 ( .A(p_input[27263]), .B(p_input[17263]), .Z(n6084) );
  AND U9126 ( .A(p_input[7263]), .B(p_input[37263]), .Z(n6083) );
  AND U9127 ( .A(n6085), .B(n6086), .Z(o[7262]) );
  AND U9128 ( .A(p_input[27262]), .B(p_input[17262]), .Z(n6086) );
  AND U9129 ( .A(p_input[7262]), .B(p_input[37262]), .Z(n6085) );
  AND U9130 ( .A(n6087), .B(n6088), .Z(o[7261]) );
  AND U9131 ( .A(p_input[27261]), .B(p_input[17261]), .Z(n6088) );
  AND U9132 ( .A(p_input[7261]), .B(p_input[37261]), .Z(n6087) );
  AND U9133 ( .A(n6089), .B(n6090), .Z(o[7260]) );
  AND U9134 ( .A(p_input[27260]), .B(p_input[17260]), .Z(n6090) );
  AND U9135 ( .A(p_input[7260]), .B(p_input[37260]), .Z(n6089) );
  AND U9136 ( .A(n6091), .B(n6092), .Z(o[725]) );
  AND U9137 ( .A(p_input[20725]), .B(p_input[10725]), .Z(n6092) );
  AND U9138 ( .A(p_input[725]), .B(p_input[30725]), .Z(n6091) );
  AND U9139 ( .A(n6093), .B(n6094), .Z(o[7259]) );
  AND U9140 ( .A(p_input[27259]), .B(p_input[17259]), .Z(n6094) );
  AND U9141 ( .A(p_input[7259]), .B(p_input[37259]), .Z(n6093) );
  AND U9142 ( .A(n6095), .B(n6096), .Z(o[7258]) );
  AND U9143 ( .A(p_input[27258]), .B(p_input[17258]), .Z(n6096) );
  AND U9144 ( .A(p_input[7258]), .B(p_input[37258]), .Z(n6095) );
  AND U9145 ( .A(n6097), .B(n6098), .Z(o[7257]) );
  AND U9146 ( .A(p_input[27257]), .B(p_input[17257]), .Z(n6098) );
  AND U9147 ( .A(p_input[7257]), .B(p_input[37257]), .Z(n6097) );
  AND U9148 ( .A(n6099), .B(n6100), .Z(o[7256]) );
  AND U9149 ( .A(p_input[27256]), .B(p_input[17256]), .Z(n6100) );
  AND U9150 ( .A(p_input[7256]), .B(p_input[37256]), .Z(n6099) );
  AND U9151 ( .A(n6101), .B(n6102), .Z(o[7255]) );
  AND U9152 ( .A(p_input[27255]), .B(p_input[17255]), .Z(n6102) );
  AND U9153 ( .A(p_input[7255]), .B(p_input[37255]), .Z(n6101) );
  AND U9154 ( .A(n6103), .B(n6104), .Z(o[7254]) );
  AND U9155 ( .A(p_input[27254]), .B(p_input[17254]), .Z(n6104) );
  AND U9156 ( .A(p_input[7254]), .B(p_input[37254]), .Z(n6103) );
  AND U9157 ( .A(n6105), .B(n6106), .Z(o[7253]) );
  AND U9158 ( .A(p_input[27253]), .B(p_input[17253]), .Z(n6106) );
  AND U9159 ( .A(p_input[7253]), .B(p_input[37253]), .Z(n6105) );
  AND U9160 ( .A(n6107), .B(n6108), .Z(o[7252]) );
  AND U9161 ( .A(p_input[27252]), .B(p_input[17252]), .Z(n6108) );
  AND U9162 ( .A(p_input[7252]), .B(p_input[37252]), .Z(n6107) );
  AND U9163 ( .A(n6109), .B(n6110), .Z(o[7251]) );
  AND U9164 ( .A(p_input[27251]), .B(p_input[17251]), .Z(n6110) );
  AND U9165 ( .A(p_input[7251]), .B(p_input[37251]), .Z(n6109) );
  AND U9166 ( .A(n6111), .B(n6112), .Z(o[7250]) );
  AND U9167 ( .A(p_input[27250]), .B(p_input[17250]), .Z(n6112) );
  AND U9168 ( .A(p_input[7250]), .B(p_input[37250]), .Z(n6111) );
  AND U9169 ( .A(n6113), .B(n6114), .Z(o[724]) );
  AND U9170 ( .A(p_input[20724]), .B(p_input[10724]), .Z(n6114) );
  AND U9171 ( .A(p_input[724]), .B(p_input[30724]), .Z(n6113) );
  AND U9172 ( .A(n6115), .B(n6116), .Z(o[7249]) );
  AND U9173 ( .A(p_input[27249]), .B(p_input[17249]), .Z(n6116) );
  AND U9174 ( .A(p_input[7249]), .B(p_input[37249]), .Z(n6115) );
  AND U9175 ( .A(n6117), .B(n6118), .Z(o[7248]) );
  AND U9176 ( .A(p_input[27248]), .B(p_input[17248]), .Z(n6118) );
  AND U9177 ( .A(p_input[7248]), .B(p_input[37248]), .Z(n6117) );
  AND U9178 ( .A(n6119), .B(n6120), .Z(o[7247]) );
  AND U9179 ( .A(p_input[27247]), .B(p_input[17247]), .Z(n6120) );
  AND U9180 ( .A(p_input[7247]), .B(p_input[37247]), .Z(n6119) );
  AND U9181 ( .A(n6121), .B(n6122), .Z(o[7246]) );
  AND U9182 ( .A(p_input[27246]), .B(p_input[17246]), .Z(n6122) );
  AND U9183 ( .A(p_input[7246]), .B(p_input[37246]), .Z(n6121) );
  AND U9184 ( .A(n6123), .B(n6124), .Z(o[7245]) );
  AND U9185 ( .A(p_input[27245]), .B(p_input[17245]), .Z(n6124) );
  AND U9186 ( .A(p_input[7245]), .B(p_input[37245]), .Z(n6123) );
  AND U9187 ( .A(n6125), .B(n6126), .Z(o[7244]) );
  AND U9188 ( .A(p_input[27244]), .B(p_input[17244]), .Z(n6126) );
  AND U9189 ( .A(p_input[7244]), .B(p_input[37244]), .Z(n6125) );
  AND U9190 ( .A(n6127), .B(n6128), .Z(o[7243]) );
  AND U9191 ( .A(p_input[27243]), .B(p_input[17243]), .Z(n6128) );
  AND U9192 ( .A(p_input[7243]), .B(p_input[37243]), .Z(n6127) );
  AND U9193 ( .A(n6129), .B(n6130), .Z(o[7242]) );
  AND U9194 ( .A(p_input[27242]), .B(p_input[17242]), .Z(n6130) );
  AND U9195 ( .A(p_input[7242]), .B(p_input[37242]), .Z(n6129) );
  AND U9196 ( .A(n6131), .B(n6132), .Z(o[7241]) );
  AND U9197 ( .A(p_input[27241]), .B(p_input[17241]), .Z(n6132) );
  AND U9198 ( .A(p_input[7241]), .B(p_input[37241]), .Z(n6131) );
  AND U9199 ( .A(n6133), .B(n6134), .Z(o[7240]) );
  AND U9200 ( .A(p_input[27240]), .B(p_input[17240]), .Z(n6134) );
  AND U9201 ( .A(p_input[7240]), .B(p_input[37240]), .Z(n6133) );
  AND U9202 ( .A(n6135), .B(n6136), .Z(o[723]) );
  AND U9203 ( .A(p_input[20723]), .B(p_input[10723]), .Z(n6136) );
  AND U9204 ( .A(p_input[723]), .B(p_input[30723]), .Z(n6135) );
  AND U9205 ( .A(n6137), .B(n6138), .Z(o[7239]) );
  AND U9206 ( .A(p_input[27239]), .B(p_input[17239]), .Z(n6138) );
  AND U9207 ( .A(p_input[7239]), .B(p_input[37239]), .Z(n6137) );
  AND U9208 ( .A(n6139), .B(n6140), .Z(o[7238]) );
  AND U9209 ( .A(p_input[27238]), .B(p_input[17238]), .Z(n6140) );
  AND U9210 ( .A(p_input[7238]), .B(p_input[37238]), .Z(n6139) );
  AND U9211 ( .A(n6141), .B(n6142), .Z(o[7237]) );
  AND U9212 ( .A(p_input[27237]), .B(p_input[17237]), .Z(n6142) );
  AND U9213 ( .A(p_input[7237]), .B(p_input[37237]), .Z(n6141) );
  AND U9214 ( .A(n6143), .B(n6144), .Z(o[7236]) );
  AND U9215 ( .A(p_input[27236]), .B(p_input[17236]), .Z(n6144) );
  AND U9216 ( .A(p_input[7236]), .B(p_input[37236]), .Z(n6143) );
  AND U9217 ( .A(n6145), .B(n6146), .Z(o[7235]) );
  AND U9218 ( .A(p_input[27235]), .B(p_input[17235]), .Z(n6146) );
  AND U9219 ( .A(p_input[7235]), .B(p_input[37235]), .Z(n6145) );
  AND U9220 ( .A(n6147), .B(n6148), .Z(o[7234]) );
  AND U9221 ( .A(p_input[27234]), .B(p_input[17234]), .Z(n6148) );
  AND U9222 ( .A(p_input[7234]), .B(p_input[37234]), .Z(n6147) );
  AND U9223 ( .A(n6149), .B(n6150), .Z(o[7233]) );
  AND U9224 ( .A(p_input[27233]), .B(p_input[17233]), .Z(n6150) );
  AND U9225 ( .A(p_input[7233]), .B(p_input[37233]), .Z(n6149) );
  AND U9226 ( .A(n6151), .B(n6152), .Z(o[7232]) );
  AND U9227 ( .A(p_input[27232]), .B(p_input[17232]), .Z(n6152) );
  AND U9228 ( .A(p_input[7232]), .B(p_input[37232]), .Z(n6151) );
  AND U9229 ( .A(n6153), .B(n6154), .Z(o[7231]) );
  AND U9230 ( .A(p_input[27231]), .B(p_input[17231]), .Z(n6154) );
  AND U9231 ( .A(p_input[7231]), .B(p_input[37231]), .Z(n6153) );
  AND U9232 ( .A(n6155), .B(n6156), .Z(o[7230]) );
  AND U9233 ( .A(p_input[27230]), .B(p_input[17230]), .Z(n6156) );
  AND U9234 ( .A(p_input[7230]), .B(p_input[37230]), .Z(n6155) );
  AND U9235 ( .A(n6157), .B(n6158), .Z(o[722]) );
  AND U9236 ( .A(p_input[20722]), .B(p_input[10722]), .Z(n6158) );
  AND U9237 ( .A(p_input[722]), .B(p_input[30722]), .Z(n6157) );
  AND U9238 ( .A(n6159), .B(n6160), .Z(o[7229]) );
  AND U9239 ( .A(p_input[27229]), .B(p_input[17229]), .Z(n6160) );
  AND U9240 ( .A(p_input[7229]), .B(p_input[37229]), .Z(n6159) );
  AND U9241 ( .A(n6161), .B(n6162), .Z(o[7228]) );
  AND U9242 ( .A(p_input[27228]), .B(p_input[17228]), .Z(n6162) );
  AND U9243 ( .A(p_input[7228]), .B(p_input[37228]), .Z(n6161) );
  AND U9244 ( .A(n6163), .B(n6164), .Z(o[7227]) );
  AND U9245 ( .A(p_input[27227]), .B(p_input[17227]), .Z(n6164) );
  AND U9246 ( .A(p_input[7227]), .B(p_input[37227]), .Z(n6163) );
  AND U9247 ( .A(n6165), .B(n6166), .Z(o[7226]) );
  AND U9248 ( .A(p_input[27226]), .B(p_input[17226]), .Z(n6166) );
  AND U9249 ( .A(p_input[7226]), .B(p_input[37226]), .Z(n6165) );
  AND U9250 ( .A(n6167), .B(n6168), .Z(o[7225]) );
  AND U9251 ( .A(p_input[27225]), .B(p_input[17225]), .Z(n6168) );
  AND U9252 ( .A(p_input[7225]), .B(p_input[37225]), .Z(n6167) );
  AND U9253 ( .A(n6169), .B(n6170), .Z(o[7224]) );
  AND U9254 ( .A(p_input[27224]), .B(p_input[17224]), .Z(n6170) );
  AND U9255 ( .A(p_input[7224]), .B(p_input[37224]), .Z(n6169) );
  AND U9256 ( .A(n6171), .B(n6172), .Z(o[7223]) );
  AND U9257 ( .A(p_input[27223]), .B(p_input[17223]), .Z(n6172) );
  AND U9258 ( .A(p_input[7223]), .B(p_input[37223]), .Z(n6171) );
  AND U9259 ( .A(n6173), .B(n6174), .Z(o[7222]) );
  AND U9260 ( .A(p_input[27222]), .B(p_input[17222]), .Z(n6174) );
  AND U9261 ( .A(p_input[7222]), .B(p_input[37222]), .Z(n6173) );
  AND U9262 ( .A(n6175), .B(n6176), .Z(o[7221]) );
  AND U9263 ( .A(p_input[27221]), .B(p_input[17221]), .Z(n6176) );
  AND U9264 ( .A(p_input[7221]), .B(p_input[37221]), .Z(n6175) );
  AND U9265 ( .A(n6177), .B(n6178), .Z(o[7220]) );
  AND U9266 ( .A(p_input[27220]), .B(p_input[17220]), .Z(n6178) );
  AND U9267 ( .A(p_input[7220]), .B(p_input[37220]), .Z(n6177) );
  AND U9268 ( .A(n6179), .B(n6180), .Z(o[721]) );
  AND U9269 ( .A(p_input[20721]), .B(p_input[10721]), .Z(n6180) );
  AND U9270 ( .A(p_input[721]), .B(p_input[30721]), .Z(n6179) );
  AND U9271 ( .A(n6181), .B(n6182), .Z(o[7219]) );
  AND U9272 ( .A(p_input[27219]), .B(p_input[17219]), .Z(n6182) );
  AND U9273 ( .A(p_input[7219]), .B(p_input[37219]), .Z(n6181) );
  AND U9274 ( .A(n6183), .B(n6184), .Z(o[7218]) );
  AND U9275 ( .A(p_input[27218]), .B(p_input[17218]), .Z(n6184) );
  AND U9276 ( .A(p_input[7218]), .B(p_input[37218]), .Z(n6183) );
  AND U9277 ( .A(n6185), .B(n6186), .Z(o[7217]) );
  AND U9278 ( .A(p_input[27217]), .B(p_input[17217]), .Z(n6186) );
  AND U9279 ( .A(p_input[7217]), .B(p_input[37217]), .Z(n6185) );
  AND U9280 ( .A(n6187), .B(n6188), .Z(o[7216]) );
  AND U9281 ( .A(p_input[27216]), .B(p_input[17216]), .Z(n6188) );
  AND U9282 ( .A(p_input[7216]), .B(p_input[37216]), .Z(n6187) );
  AND U9283 ( .A(n6189), .B(n6190), .Z(o[7215]) );
  AND U9284 ( .A(p_input[27215]), .B(p_input[17215]), .Z(n6190) );
  AND U9285 ( .A(p_input[7215]), .B(p_input[37215]), .Z(n6189) );
  AND U9286 ( .A(n6191), .B(n6192), .Z(o[7214]) );
  AND U9287 ( .A(p_input[27214]), .B(p_input[17214]), .Z(n6192) );
  AND U9288 ( .A(p_input[7214]), .B(p_input[37214]), .Z(n6191) );
  AND U9289 ( .A(n6193), .B(n6194), .Z(o[7213]) );
  AND U9290 ( .A(p_input[27213]), .B(p_input[17213]), .Z(n6194) );
  AND U9291 ( .A(p_input[7213]), .B(p_input[37213]), .Z(n6193) );
  AND U9292 ( .A(n6195), .B(n6196), .Z(o[7212]) );
  AND U9293 ( .A(p_input[27212]), .B(p_input[17212]), .Z(n6196) );
  AND U9294 ( .A(p_input[7212]), .B(p_input[37212]), .Z(n6195) );
  AND U9295 ( .A(n6197), .B(n6198), .Z(o[7211]) );
  AND U9296 ( .A(p_input[27211]), .B(p_input[17211]), .Z(n6198) );
  AND U9297 ( .A(p_input[7211]), .B(p_input[37211]), .Z(n6197) );
  AND U9298 ( .A(n6199), .B(n6200), .Z(o[7210]) );
  AND U9299 ( .A(p_input[27210]), .B(p_input[17210]), .Z(n6200) );
  AND U9300 ( .A(p_input[7210]), .B(p_input[37210]), .Z(n6199) );
  AND U9301 ( .A(n6201), .B(n6202), .Z(o[720]) );
  AND U9302 ( .A(p_input[20720]), .B(p_input[10720]), .Z(n6202) );
  AND U9303 ( .A(p_input[720]), .B(p_input[30720]), .Z(n6201) );
  AND U9304 ( .A(n6203), .B(n6204), .Z(o[7209]) );
  AND U9305 ( .A(p_input[27209]), .B(p_input[17209]), .Z(n6204) );
  AND U9306 ( .A(p_input[7209]), .B(p_input[37209]), .Z(n6203) );
  AND U9307 ( .A(n6205), .B(n6206), .Z(o[7208]) );
  AND U9308 ( .A(p_input[27208]), .B(p_input[17208]), .Z(n6206) );
  AND U9309 ( .A(p_input[7208]), .B(p_input[37208]), .Z(n6205) );
  AND U9310 ( .A(n6207), .B(n6208), .Z(o[7207]) );
  AND U9311 ( .A(p_input[27207]), .B(p_input[17207]), .Z(n6208) );
  AND U9312 ( .A(p_input[7207]), .B(p_input[37207]), .Z(n6207) );
  AND U9313 ( .A(n6209), .B(n6210), .Z(o[7206]) );
  AND U9314 ( .A(p_input[27206]), .B(p_input[17206]), .Z(n6210) );
  AND U9315 ( .A(p_input[7206]), .B(p_input[37206]), .Z(n6209) );
  AND U9316 ( .A(n6211), .B(n6212), .Z(o[7205]) );
  AND U9317 ( .A(p_input[27205]), .B(p_input[17205]), .Z(n6212) );
  AND U9318 ( .A(p_input[7205]), .B(p_input[37205]), .Z(n6211) );
  AND U9319 ( .A(n6213), .B(n6214), .Z(o[7204]) );
  AND U9320 ( .A(p_input[27204]), .B(p_input[17204]), .Z(n6214) );
  AND U9321 ( .A(p_input[7204]), .B(p_input[37204]), .Z(n6213) );
  AND U9322 ( .A(n6215), .B(n6216), .Z(o[7203]) );
  AND U9323 ( .A(p_input[27203]), .B(p_input[17203]), .Z(n6216) );
  AND U9324 ( .A(p_input[7203]), .B(p_input[37203]), .Z(n6215) );
  AND U9325 ( .A(n6217), .B(n6218), .Z(o[7202]) );
  AND U9326 ( .A(p_input[27202]), .B(p_input[17202]), .Z(n6218) );
  AND U9327 ( .A(p_input[7202]), .B(p_input[37202]), .Z(n6217) );
  AND U9328 ( .A(n6219), .B(n6220), .Z(o[7201]) );
  AND U9329 ( .A(p_input[27201]), .B(p_input[17201]), .Z(n6220) );
  AND U9330 ( .A(p_input[7201]), .B(p_input[37201]), .Z(n6219) );
  AND U9331 ( .A(n6221), .B(n6222), .Z(o[7200]) );
  AND U9332 ( .A(p_input[27200]), .B(p_input[17200]), .Z(n6222) );
  AND U9333 ( .A(p_input[7200]), .B(p_input[37200]), .Z(n6221) );
  AND U9334 ( .A(n6223), .B(n6224), .Z(o[71]) );
  AND U9335 ( .A(p_input[20071]), .B(p_input[10071]), .Z(n6224) );
  AND U9336 ( .A(p_input[71]), .B(p_input[30071]), .Z(n6223) );
  AND U9337 ( .A(n6225), .B(n6226), .Z(o[719]) );
  AND U9338 ( .A(p_input[20719]), .B(p_input[10719]), .Z(n6226) );
  AND U9339 ( .A(p_input[719]), .B(p_input[30719]), .Z(n6225) );
  AND U9340 ( .A(n6227), .B(n6228), .Z(o[7199]) );
  AND U9341 ( .A(p_input[27199]), .B(p_input[17199]), .Z(n6228) );
  AND U9342 ( .A(p_input[7199]), .B(p_input[37199]), .Z(n6227) );
  AND U9343 ( .A(n6229), .B(n6230), .Z(o[7198]) );
  AND U9344 ( .A(p_input[27198]), .B(p_input[17198]), .Z(n6230) );
  AND U9345 ( .A(p_input[7198]), .B(p_input[37198]), .Z(n6229) );
  AND U9346 ( .A(n6231), .B(n6232), .Z(o[7197]) );
  AND U9347 ( .A(p_input[27197]), .B(p_input[17197]), .Z(n6232) );
  AND U9348 ( .A(p_input[7197]), .B(p_input[37197]), .Z(n6231) );
  AND U9349 ( .A(n6233), .B(n6234), .Z(o[7196]) );
  AND U9350 ( .A(p_input[27196]), .B(p_input[17196]), .Z(n6234) );
  AND U9351 ( .A(p_input[7196]), .B(p_input[37196]), .Z(n6233) );
  AND U9352 ( .A(n6235), .B(n6236), .Z(o[7195]) );
  AND U9353 ( .A(p_input[27195]), .B(p_input[17195]), .Z(n6236) );
  AND U9354 ( .A(p_input[7195]), .B(p_input[37195]), .Z(n6235) );
  AND U9355 ( .A(n6237), .B(n6238), .Z(o[7194]) );
  AND U9356 ( .A(p_input[27194]), .B(p_input[17194]), .Z(n6238) );
  AND U9357 ( .A(p_input[7194]), .B(p_input[37194]), .Z(n6237) );
  AND U9358 ( .A(n6239), .B(n6240), .Z(o[7193]) );
  AND U9359 ( .A(p_input[27193]), .B(p_input[17193]), .Z(n6240) );
  AND U9360 ( .A(p_input[7193]), .B(p_input[37193]), .Z(n6239) );
  AND U9361 ( .A(n6241), .B(n6242), .Z(o[7192]) );
  AND U9362 ( .A(p_input[27192]), .B(p_input[17192]), .Z(n6242) );
  AND U9363 ( .A(p_input[7192]), .B(p_input[37192]), .Z(n6241) );
  AND U9364 ( .A(n6243), .B(n6244), .Z(o[7191]) );
  AND U9365 ( .A(p_input[27191]), .B(p_input[17191]), .Z(n6244) );
  AND U9366 ( .A(p_input[7191]), .B(p_input[37191]), .Z(n6243) );
  AND U9367 ( .A(n6245), .B(n6246), .Z(o[7190]) );
  AND U9368 ( .A(p_input[27190]), .B(p_input[17190]), .Z(n6246) );
  AND U9369 ( .A(p_input[7190]), .B(p_input[37190]), .Z(n6245) );
  AND U9370 ( .A(n6247), .B(n6248), .Z(o[718]) );
  AND U9371 ( .A(p_input[20718]), .B(p_input[10718]), .Z(n6248) );
  AND U9372 ( .A(p_input[718]), .B(p_input[30718]), .Z(n6247) );
  AND U9373 ( .A(n6249), .B(n6250), .Z(o[7189]) );
  AND U9374 ( .A(p_input[27189]), .B(p_input[17189]), .Z(n6250) );
  AND U9375 ( .A(p_input[7189]), .B(p_input[37189]), .Z(n6249) );
  AND U9376 ( .A(n6251), .B(n6252), .Z(o[7188]) );
  AND U9377 ( .A(p_input[27188]), .B(p_input[17188]), .Z(n6252) );
  AND U9378 ( .A(p_input[7188]), .B(p_input[37188]), .Z(n6251) );
  AND U9379 ( .A(n6253), .B(n6254), .Z(o[7187]) );
  AND U9380 ( .A(p_input[27187]), .B(p_input[17187]), .Z(n6254) );
  AND U9381 ( .A(p_input[7187]), .B(p_input[37187]), .Z(n6253) );
  AND U9382 ( .A(n6255), .B(n6256), .Z(o[7186]) );
  AND U9383 ( .A(p_input[27186]), .B(p_input[17186]), .Z(n6256) );
  AND U9384 ( .A(p_input[7186]), .B(p_input[37186]), .Z(n6255) );
  AND U9385 ( .A(n6257), .B(n6258), .Z(o[7185]) );
  AND U9386 ( .A(p_input[27185]), .B(p_input[17185]), .Z(n6258) );
  AND U9387 ( .A(p_input[7185]), .B(p_input[37185]), .Z(n6257) );
  AND U9388 ( .A(n6259), .B(n6260), .Z(o[7184]) );
  AND U9389 ( .A(p_input[27184]), .B(p_input[17184]), .Z(n6260) );
  AND U9390 ( .A(p_input[7184]), .B(p_input[37184]), .Z(n6259) );
  AND U9391 ( .A(n6261), .B(n6262), .Z(o[7183]) );
  AND U9392 ( .A(p_input[27183]), .B(p_input[17183]), .Z(n6262) );
  AND U9393 ( .A(p_input[7183]), .B(p_input[37183]), .Z(n6261) );
  AND U9394 ( .A(n6263), .B(n6264), .Z(o[7182]) );
  AND U9395 ( .A(p_input[27182]), .B(p_input[17182]), .Z(n6264) );
  AND U9396 ( .A(p_input[7182]), .B(p_input[37182]), .Z(n6263) );
  AND U9397 ( .A(n6265), .B(n6266), .Z(o[7181]) );
  AND U9398 ( .A(p_input[27181]), .B(p_input[17181]), .Z(n6266) );
  AND U9399 ( .A(p_input[7181]), .B(p_input[37181]), .Z(n6265) );
  AND U9400 ( .A(n6267), .B(n6268), .Z(o[7180]) );
  AND U9401 ( .A(p_input[27180]), .B(p_input[17180]), .Z(n6268) );
  AND U9402 ( .A(p_input[7180]), .B(p_input[37180]), .Z(n6267) );
  AND U9403 ( .A(n6269), .B(n6270), .Z(o[717]) );
  AND U9404 ( .A(p_input[20717]), .B(p_input[10717]), .Z(n6270) );
  AND U9405 ( .A(p_input[717]), .B(p_input[30717]), .Z(n6269) );
  AND U9406 ( .A(n6271), .B(n6272), .Z(o[7179]) );
  AND U9407 ( .A(p_input[27179]), .B(p_input[17179]), .Z(n6272) );
  AND U9408 ( .A(p_input[7179]), .B(p_input[37179]), .Z(n6271) );
  AND U9409 ( .A(n6273), .B(n6274), .Z(o[7178]) );
  AND U9410 ( .A(p_input[27178]), .B(p_input[17178]), .Z(n6274) );
  AND U9411 ( .A(p_input[7178]), .B(p_input[37178]), .Z(n6273) );
  AND U9412 ( .A(n6275), .B(n6276), .Z(o[7177]) );
  AND U9413 ( .A(p_input[27177]), .B(p_input[17177]), .Z(n6276) );
  AND U9414 ( .A(p_input[7177]), .B(p_input[37177]), .Z(n6275) );
  AND U9415 ( .A(n6277), .B(n6278), .Z(o[7176]) );
  AND U9416 ( .A(p_input[27176]), .B(p_input[17176]), .Z(n6278) );
  AND U9417 ( .A(p_input[7176]), .B(p_input[37176]), .Z(n6277) );
  AND U9418 ( .A(n6279), .B(n6280), .Z(o[7175]) );
  AND U9419 ( .A(p_input[27175]), .B(p_input[17175]), .Z(n6280) );
  AND U9420 ( .A(p_input[7175]), .B(p_input[37175]), .Z(n6279) );
  AND U9421 ( .A(n6281), .B(n6282), .Z(o[7174]) );
  AND U9422 ( .A(p_input[27174]), .B(p_input[17174]), .Z(n6282) );
  AND U9423 ( .A(p_input[7174]), .B(p_input[37174]), .Z(n6281) );
  AND U9424 ( .A(n6283), .B(n6284), .Z(o[7173]) );
  AND U9425 ( .A(p_input[27173]), .B(p_input[17173]), .Z(n6284) );
  AND U9426 ( .A(p_input[7173]), .B(p_input[37173]), .Z(n6283) );
  AND U9427 ( .A(n6285), .B(n6286), .Z(o[7172]) );
  AND U9428 ( .A(p_input[27172]), .B(p_input[17172]), .Z(n6286) );
  AND U9429 ( .A(p_input[7172]), .B(p_input[37172]), .Z(n6285) );
  AND U9430 ( .A(n6287), .B(n6288), .Z(o[7171]) );
  AND U9431 ( .A(p_input[27171]), .B(p_input[17171]), .Z(n6288) );
  AND U9432 ( .A(p_input[7171]), .B(p_input[37171]), .Z(n6287) );
  AND U9433 ( .A(n6289), .B(n6290), .Z(o[7170]) );
  AND U9434 ( .A(p_input[27170]), .B(p_input[17170]), .Z(n6290) );
  AND U9435 ( .A(p_input[7170]), .B(p_input[37170]), .Z(n6289) );
  AND U9436 ( .A(n6291), .B(n6292), .Z(o[716]) );
  AND U9437 ( .A(p_input[20716]), .B(p_input[10716]), .Z(n6292) );
  AND U9438 ( .A(p_input[716]), .B(p_input[30716]), .Z(n6291) );
  AND U9439 ( .A(n6293), .B(n6294), .Z(o[7169]) );
  AND U9440 ( .A(p_input[27169]), .B(p_input[17169]), .Z(n6294) );
  AND U9441 ( .A(p_input[7169]), .B(p_input[37169]), .Z(n6293) );
  AND U9442 ( .A(n6295), .B(n6296), .Z(o[7168]) );
  AND U9443 ( .A(p_input[27168]), .B(p_input[17168]), .Z(n6296) );
  AND U9444 ( .A(p_input[7168]), .B(p_input[37168]), .Z(n6295) );
  AND U9445 ( .A(n6297), .B(n6298), .Z(o[7167]) );
  AND U9446 ( .A(p_input[27167]), .B(p_input[17167]), .Z(n6298) );
  AND U9447 ( .A(p_input[7167]), .B(p_input[37167]), .Z(n6297) );
  AND U9448 ( .A(n6299), .B(n6300), .Z(o[7166]) );
  AND U9449 ( .A(p_input[27166]), .B(p_input[17166]), .Z(n6300) );
  AND U9450 ( .A(p_input[7166]), .B(p_input[37166]), .Z(n6299) );
  AND U9451 ( .A(n6301), .B(n6302), .Z(o[7165]) );
  AND U9452 ( .A(p_input[27165]), .B(p_input[17165]), .Z(n6302) );
  AND U9453 ( .A(p_input[7165]), .B(p_input[37165]), .Z(n6301) );
  AND U9454 ( .A(n6303), .B(n6304), .Z(o[7164]) );
  AND U9455 ( .A(p_input[27164]), .B(p_input[17164]), .Z(n6304) );
  AND U9456 ( .A(p_input[7164]), .B(p_input[37164]), .Z(n6303) );
  AND U9457 ( .A(n6305), .B(n6306), .Z(o[7163]) );
  AND U9458 ( .A(p_input[27163]), .B(p_input[17163]), .Z(n6306) );
  AND U9459 ( .A(p_input[7163]), .B(p_input[37163]), .Z(n6305) );
  AND U9460 ( .A(n6307), .B(n6308), .Z(o[7162]) );
  AND U9461 ( .A(p_input[27162]), .B(p_input[17162]), .Z(n6308) );
  AND U9462 ( .A(p_input[7162]), .B(p_input[37162]), .Z(n6307) );
  AND U9463 ( .A(n6309), .B(n6310), .Z(o[7161]) );
  AND U9464 ( .A(p_input[27161]), .B(p_input[17161]), .Z(n6310) );
  AND U9465 ( .A(p_input[7161]), .B(p_input[37161]), .Z(n6309) );
  AND U9466 ( .A(n6311), .B(n6312), .Z(o[7160]) );
  AND U9467 ( .A(p_input[27160]), .B(p_input[17160]), .Z(n6312) );
  AND U9468 ( .A(p_input[7160]), .B(p_input[37160]), .Z(n6311) );
  AND U9469 ( .A(n6313), .B(n6314), .Z(o[715]) );
  AND U9470 ( .A(p_input[20715]), .B(p_input[10715]), .Z(n6314) );
  AND U9471 ( .A(p_input[715]), .B(p_input[30715]), .Z(n6313) );
  AND U9472 ( .A(n6315), .B(n6316), .Z(o[7159]) );
  AND U9473 ( .A(p_input[27159]), .B(p_input[17159]), .Z(n6316) );
  AND U9474 ( .A(p_input[7159]), .B(p_input[37159]), .Z(n6315) );
  AND U9475 ( .A(n6317), .B(n6318), .Z(o[7158]) );
  AND U9476 ( .A(p_input[27158]), .B(p_input[17158]), .Z(n6318) );
  AND U9477 ( .A(p_input[7158]), .B(p_input[37158]), .Z(n6317) );
  AND U9478 ( .A(n6319), .B(n6320), .Z(o[7157]) );
  AND U9479 ( .A(p_input[27157]), .B(p_input[17157]), .Z(n6320) );
  AND U9480 ( .A(p_input[7157]), .B(p_input[37157]), .Z(n6319) );
  AND U9481 ( .A(n6321), .B(n6322), .Z(o[7156]) );
  AND U9482 ( .A(p_input[27156]), .B(p_input[17156]), .Z(n6322) );
  AND U9483 ( .A(p_input[7156]), .B(p_input[37156]), .Z(n6321) );
  AND U9484 ( .A(n6323), .B(n6324), .Z(o[7155]) );
  AND U9485 ( .A(p_input[27155]), .B(p_input[17155]), .Z(n6324) );
  AND U9486 ( .A(p_input[7155]), .B(p_input[37155]), .Z(n6323) );
  AND U9487 ( .A(n6325), .B(n6326), .Z(o[7154]) );
  AND U9488 ( .A(p_input[27154]), .B(p_input[17154]), .Z(n6326) );
  AND U9489 ( .A(p_input[7154]), .B(p_input[37154]), .Z(n6325) );
  AND U9490 ( .A(n6327), .B(n6328), .Z(o[7153]) );
  AND U9491 ( .A(p_input[27153]), .B(p_input[17153]), .Z(n6328) );
  AND U9492 ( .A(p_input[7153]), .B(p_input[37153]), .Z(n6327) );
  AND U9493 ( .A(n6329), .B(n6330), .Z(o[7152]) );
  AND U9494 ( .A(p_input[27152]), .B(p_input[17152]), .Z(n6330) );
  AND U9495 ( .A(p_input[7152]), .B(p_input[37152]), .Z(n6329) );
  AND U9496 ( .A(n6331), .B(n6332), .Z(o[7151]) );
  AND U9497 ( .A(p_input[27151]), .B(p_input[17151]), .Z(n6332) );
  AND U9498 ( .A(p_input[7151]), .B(p_input[37151]), .Z(n6331) );
  AND U9499 ( .A(n6333), .B(n6334), .Z(o[7150]) );
  AND U9500 ( .A(p_input[27150]), .B(p_input[17150]), .Z(n6334) );
  AND U9501 ( .A(p_input[7150]), .B(p_input[37150]), .Z(n6333) );
  AND U9502 ( .A(n6335), .B(n6336), .Z(o[714]) );
  AND U9503 ( .A(p_input[20714]), .B(p_input[10714]), .Z(n6336) );
  AND U9504 ( .A(p_input[714]), .B(p_input[30714]), .Z(n6335) );
  AND U9505 ( .A(n6337), .B(n6338), .Z(o[7149]) );
  AND U9506 ( .A(p_input[27149]), .B(p_input[17149]), .Z(n6338) );
  AND U9507 ( .A(p_input[7149]), .B(p_input[37149]), .Z(n6337) );
  AND U9508 ( .A(n6339), .B(n6340), .Z(o[7148]) );
  AND U9509 ( .A(p_input[27148]), .B(p_input[17148]), .Z(n6340) );
  AND U9510 ( .A(p_input[7148]), .B(p_input[37148]), .Z(n6339) );
  AND U9511 ( .A(n6341), .B(n6342), .Z(o[7147]) );
  AND U9512 ( .A(p_input[27147]), .B(p_input[17147]), .Z(n6342) );
  AND U9513 ( .A(p_input[7147]), .B(p_input[37147]), .Z(n6341) );
  AND U9514 ( .A(n6343), .B(n6344), .Z(o[7146]) );
  AND U9515 ( .A(p_input[27146]), .B(p_input[17146]), .Z(n6344) );
  AND U9516 ( .A(p_input[7146]), .B(p_input[37146]), .Z(n6343) );
  AND U9517 ( .A(n6345), .B(n6346), .Z(o[7145]) );
  AND U9518 ( .A(p_input[27145]), .B(p_input[17145]), .Z(n6346) );
  AND U9519 ( .A(p_input[7145]), .B(p_input[37145]), .Z(n6345) );
  AND U9520 ( .A(n6347), .B(n6348), .Z(o[7144]) );
  AND U9521 ( .A(p_input[27144]), .B(p_input[17144]), .Z(n6348) );
  AND U9522 ( .A(p_input[7144]), .B(p_input[37144]), .Z(n6347) );
  AND U9523 ( .A(n6349), .B(n6350), .Z(o[7143]) );
  AND U9524 ( .A(p_input[27143]), .B(p_input[17143]), .Z(n6350) );
  AND U9525 ( .A(p_input[7143]), .B(p_input[37143]), .Z(n6349) );
  AND U9526 ( .A(n6351), .B(n6352), .Z(o[7142]) );
  AND U9527 ( .A(p_input[27142]), .B(p_input[17142]), .Z(n6352) );
  AND U9528 ( .A(p_input[7142]), .B(p_input[37142]), .Z(n6351) );
  AND U9529 ( .A(n6353), .B(n6354), .Z(o[7141]) );
  AND U9530 ( .A(p_input[27141]), .B(p_input[17141]), .Z(n6354) );
  AND U9531 ( .A(p_input[7141]), .B(p_input[37141]), .Z(n6353) );
  AND U9532 ( .A(n6355), .B(n6356), .Z(o[7140]) );
  AND U9533 ( .A(p_input[27140]), .B(p_input[17140]), .Z(n6356) );
  AND U9534 ( .A(p_input[7140]), .B(p_input[37140]), .Z(n6355) );
  AND U9535 ( .A(n6357), .B(n6358), .Z(o[713]) );
  AND U9536 ( .A(p_input[20713]), .B(p_input[10713]), .Z(n6358) );
  AND U9537 ( .A(p_input[713]), .B(p_input[30713]), .Z(n6357) );
  AND U9538 ( .A(n6359), .B(n6360), .Z(o[7139]) );
  AND U9539 ( .A(p_input[27139]), .B(p_input[17139]), .Z(n6360) );
  AND U9540 ( .A(p_input[7139]), .B(p_input[37139]), .Z(n6359) );
  AND U9541 ( .A(n6361), .B(n6362), .Z(o[7138]) );
  AND U9542 ( .A(p_input[27138]), .B(p_input[17138]), .Z(n6362) );
  AND U9543 ( .A(p_input[7138]), .B(p_input[37138]), .Z(n6361) );
  AND U9544 ( .A(n6363), .B(n6364), .Z(o[7137]) );
  AND U9545 ( .A(p_input[27137]), .B(p_input[17137]), .Z(n6364) );
  AND U9546 ( .A(p_input[7137]), .B(p_input[37137]), .Z(n6363) );
  AND U9547 ( .A(n6365), .B(n6366), .Z(o[7136]) );
  AND U9548 ( .A(p_input[27136]), .B(p_input[17136]), .Z(n6366) );
  AND U9549 ( .A(p_input[7136]), .B(p_input[37136]), .Z(n6365) );
  AND U9550 ( .A(n6367), .B(n6368), .Z(o[7135]) );
  AND U9551 ( .A(p_input[27135]), .B(p_input[17135]), .Z(n6368) );
  AND U9552 ( .A(p_input[7135]), .B(p_input[37135]), .Z(n6367) );
  AND U9553 ( .A(n6369), .B(n6370), .Z(o[7134]) );
  AND U9554 ( .A(p_input[27134]), .B(p_input[17134]), .Z(n6370) );
  AND U9555 ( .A(p_input[7134]), .B(p_input[37134]), .Z(n6369) );
  AND U9556 ( .A(n6371), .B(n6372), .Z(o[7133]) );
  AND U9557 ( .A(p_input[27133]), .B(p_input[17133]), .Z(n6372) );
  AND U9558 ( .A(p_input[7133]), .B(p_input[37133]), .Z(n6371) );
  AND U9559 ( .A(n6373), .B(n6374), .Z(o[7132]) );
  AND U9560 ( .A(p_input[27132]), .B(p_input[17132]), .Z(n6374) );
  AND U9561 ( .A(p_input[7132]), .B(p_input[37132]), .Z(n6373) );
  AND U9562 ( .A(n6375), .B(n6376), .Z(o[7131]) );
  AND U9563 ( .A(p_input[27131]), .B(p_input[17131]), .Z(n6376) );
  AND U9564 ( .A(p_input[7131]), .B(p_input[37131]), .Z(n6375) );
  AND U9565 ( .A(n6377), .B(n6378), .Z(o[7130]) );
  AND U9566 ( .A(p_input[27130]), .B(p_input[17130]), .Z(n6378) );
  AND U9567 ( .A(p_input[7130]), .B(p_input[37130]), .Z(n6377) );
  AND U9568 ( .A(n6379), .B(n6380), .Z(o[712]) );
  AND U9569 ( .A(p_input[20712]), .B(p_input[10712]), .Z(n6380) );
  AND U9570 ( .A(p_input[712]), .B(p_input[30712]), .Z(n6379) );
  AND U9571 ( .A(n6381), .B(n6382), .Z(o[7129]) );
  AND U9572 ( .A(p_input[27129]), .B(p_input[17129]), .Z(n6382) );
  AND U9573 ( .A(p_input[7129]), .B(p_input[37129]), .Z(n6381) );
  AND U9574 ( .A(n6383), .B(n6384), .Z(o[7128]) );
  AND U9575 ( .A(p_input[27128]), .B(p_input[17128]), .Z(n6384) );
  AND U9576 ( .A(p_input[7128]), .B(p_input[37128]), .Z(n6383) );
  AND U9577 ( .A(n6385), .B(n6386), .Z(o[7127]) );
  AND U9578 ( .A(p_input[27127]), .B(p_input[17127]), .Z(n6386) );
  AND U9579 ( .A(p_input[7127]), .B(p_input[37127]), .Z(n6385) );
  AND U9580 ( .A(n6387), .B(n6388), .Z(o[7126]) );
  AND U9581 ( .A(p_input[27126]), .B(p_input[17126]), .Z(n6388) );
  AND U9582 ( .A(p_input[7126]), .B(p_input[37126]), .Z(n6387) );
  AND U9583 ( .A(n6389), .B(n6390), .Z(o[7125]) );
  AND U9584 ( .A(p_input[27125]), .B(p_input[17125]), .Z(n6390) );
  AND U9585 ( .A(p_input[7125]), .B(p_input[37125]), .Z(n6389) );
  AND U9586 ( .A(n6391), .B(n6392), .Z(o[7124]) );
  AND U9587 ( .A(p_input[27124]), .B(p_input[17124]), .Z(n6392) );
  AND U9588 ( .A(p_input[7124]), .B(p_input[37124]), .Z(n6391) );
  AND U9589 ( .A(n6393), .B(n6394), .Z(o[7123]) );
  AND U9590 ( .A(p_input[27123]), .B(p_input[17123]), .Z(n6394) );
  AND U9591 ( .A(p_input[7123]), .B(p_input[37123]), .Z(n6393) );
  AND U9592 ( .A(n6395), .B(n6396), .Z(o[7122]) );
  AND U9593 ( .A(p_input[27122]), .B(p_input[17122]), .Z(n6396) );
  AND U9594 ( .A(p_input[7122]), .B(p_input[37122]), .Z(n6395) );
  AND U9595 ( .A(n6397), .B(n6398), .Z(o[7121]) );
  AND U9596 ( .A(p_input[27121]), .B(p_input[17121]), .Z(n6398) );
  AND U9597 ( .A(p_input[7121]), .B(p_input[37121]), .Z(n6397) );
  AND U9598 ( .A(n6399), .B(n6400), .Z(o[7120]) );
  AND U9599 ( .A(p_input[27120]), .B(p_input[17120]), .Z(n6400) );
  AND U9600 ( .A(p_input[7120]), .B(p_input[37120]), .Z(n6399) );
  AND U9601 ( .A(n6401), .B(n6402), .Z(o[711]) );
  AND U9602 ( .A(p_input[20711]), .B(p_input[10711]), .Z(n6402) );
  AND U9603 ( .A(p_input[711]), .B(p_input[30711]), .Z(n6401) );
  AND U9604 ( .A(n6403), .B(n6404), .Z(o[7119]) );
  AND U9605 ( .A(p_input[27119]), .B(p_input[17119]), .Z(n6404) );
  AND U9606 ( .A(p_input[7119]), .B(p_input[37119]), .Z(n6403) );
  AND U9607 ( .A(n6405), .B(n6406), .Z(o[7118]) );
  AND U9608 ( .A(p_input[27118]), .B(p_input[17118]), .Z(n6406) );
  AND U9609 ( .A(p_input[7118]), .B(p_input[37118]), .Z(n6405) );
  AND U9610 ( .A(n6407), .B(n6408), .Z(o[7117]) );
  AND U9611 ( .A(p_input[27117]), .B(p_input[17117]), .Z(n6408) );
  AND U9612 ( .A(p_input[7117]), .B(p_input[37117]), .Z(n6407) );
  AND U9613 ( .A(n6409), .B(n6410), .Z(o[7116]) );
  AND U9614 ( .A(p_input[27116]), .B(p_input[17116]), .Z(n6410) );
  AND U9615 ( .A(p_input[7116]), .B(p_input[37116]), .Z(n6409) );
  AND U9616 ( .A(n6411), .B(n6412), .Z(o[7115]) );
  AND U9617 ( .A(p_input[27115]), .B(p_input[17115]), .Z(n6412) );
  AND U9618 ( .A(p_input[7115]), .B(p_input[37115]), .Z(n6411) );
  AND U9619 ( .A(n6413), .B(n6414), .Z(o[7114]) );
  AND U9620 ( .A(p_input[27114]), .B(p_input[17114]), .Z(n6414) );
  AND U9621 ( .A(p_input[7114]), .B(p_input[37114]), .Z(n6413) );
  AND U9622 ( .A(n6415), .B(n6416), .Z(o[7113]) );
  AND U9623 ( .A(p_input[27113]), .B(p_input[17113]), .Z(n6416) );
  AND U9624 ( .A(p_input[7113]), .B(p_input[37113]), .Z(n6415) );
  AND U9625 ( .A(n6417), .B(n6418), .Z(o[7112]) );
  AND U9626 ( .A(p_input[27112]), .B(p_input[17112]), .Z(n6418) );
  AND U9627 ( .A(p_input[7112]), .B(p_input[37112]), .Z(n6417) );
  AND U9628 ( .A(n6419), .B(n6420), .Z(o[7111]) );
  AND U9629 ( .A(p_input[27111]), .B(p_input[17111]), .Z(n6420) );
  AND U9630 ( .A(p_input[7111]), .B(p_input[37111]), .Z(n6419) );
  AND U9631 ( .A(n6421), .B(n6422), .Z(o[7110]) );
  AND U9632 ( .A(p_input[27110]), .B(p_input[17110]), .Z(n6422) );
  AND U9633 ( .A(p_input[7110]), .B(p_input[37110]), .Z(n6421) );
  AND U9634 ( .A(n6423), .B(n6424), .Z(o[710]) );
  AND U9635 ( .A(p_input[20710]), .B(p_input[10710]), .Z(n6424) );
  AND U9636 ( .A(p_input[710]), .B(p_input[30710]), .Z(n6423) );
  AND U9637 ( .A(n6425), .B(n6426), .Z(o[7109]) );
  AND U9638 ( .A(p_input[27109]), .B(p_input[17109]), .Z(n6426) );
  AND U9639 ( .A(p_input[7109]), .B(p_input[37109]), .Z(n6425) );
  AND U9640 ( .A(n6427), .B(n6428), .Z(o[7108]) );
  AND U9641 ( .A(p_input[27108]), .B(p_input[17108]), .Z(n6428) );
  AND U9642 ( .A(p_input[7108]), .B(p_input[37108]), .Z(n6427) );
  AND U9643 ( .A(n6429), .B(n6430), .Z(o[7107]) );
  AND U9644 ( .A(p_input[27107]), .B(p_input[17107]), .Z(n6430) );
  AND U9645 ( .A(p_input[7107]), .B(p_input[37107]), .Z(n6429) );
  AND U9646 ( .A(n6431), .B(n6432), .Z(o[7106]) );
  AND U9647 ( .A(p_input[27106]), .B(p_input[17106]), .Z(n6432) );
  AND U9648 ( .A(p_input[7106]), .B(p_input[37106]), .Z(n6431) );
  AND U9649 ( .A(n6433), .B(n6434), .Z(o[7105]) );
  AND U9650 ( .A(p_input[27105]), .B(p_input[17105]), .Z(n6434) );
  AND U9651 ( .A(p_input[7105]), .B(p_input[37105]), .Z(n6433) );
  AND U9652 ( .A(n6435), .B(n6436), .Z(o[7104]) );
  AND U9653 ( .A(p_input[27104]), .B(p_input[17104]), .Z(n6436) );
  AND U9654 ( .A(p_input[7104]), .B(p_input[37104]), .Z(n6435) );
  AND U9655 ( .A(n6437), .B(n6438), .Z(o[7103]) );
  AND U9656 ( .A(p_input[27103]), .B(p_input[17103]), .Z(n6438) );
  AND U9657 ( .A(p_input[7103]), .B(p_input[37103]), .Z(n6437) );
  AND U9658 ( .A(n6439), .B(n6440), .Z(o[7102]) );
  AND U9659 ( .A(p_input[27102]), .B(p_input[17102]), .Z(n6440) );
  AND U9660 ( .A(p_input[7102]), .B(p_input[37102]), .Z(n6439) );
  AND U9661 ( .A(n6441), .B(n6442), .Z(o[7101]) );
  AND U9662 ( .A(p_input[27101]), .B(p_input[17101]), .Z(n6442) );
  AND U9663 ( .A(p_input[7101]), .B(p_input[37101]), .Z(n6441) );
  AND U9664 ( .A(n6443), .B(n6444), .Z(o[7100]) );
  AND U9665 ( .A(p_input[27100]), .B(p_input[17100]), .Z(n6444) );
  AND U9666 ( .A(p_input[7100]), .B(p_input[37100]), .Z(n6443) );
  AND U9667 ( .A(n6445), .B(n6446), .Z(o[70]) );
  AND U9668 ( .A(p_input[20070]), .B(p_input[10070]), .Z(n6446) );
  AND U9669 ( .A(p_input[70]), .B(p_input[30070]), .Z(n6445) );
  AND U9670 ( .A(n6447), .B(n6448), .Z(o[709]) );
  AND U9671 ( .A(p_input[20709]), .B(p_input[10709]), .Z(n6448) );
  AND U9672 ( .A(p_input[709]), .B(p_input[30709]), .Z(n6447) );
  AND U9673 ( .A(n6449), .B(n6450), .Z(o[7099]) );
  AND U9674 ( .A(p_input[27099]), .B(p_input[17099]), .Z(n6450) );
  AND U9675 ( .A(p_input[7099]), .B(p_input[37099]), .Z(n6449) );
  AND U9676 ( .A(n6451), .B(n6452), .Z(o[7098]) );
  AND U9677 ( .A(p_input[27098]), .B(p_input[17098]), .Z(n6452) );
  AND U9678 ( .A(p_input[7098]), .B(p_input[37098]), .Z(n6451) );
  AND U9679 ( .A(n6453), .B(n6454), .Z(o[7097]) );
  AND U9680 ( .A(p_input[27097]), .B(p_input[17097]), .Z(n6454) );
  AND U9681 ( .A(p_input[7097]), .B(p_input[37097]), .Z(n6453) );
  AND U9682 ( .A(n6455), .B(n6456), .Z(o[7096]) );
  AND U9683 ( .A(p_input[27096]), .B(p_input[17096]), .Z(n6456) );
  AND U9684 ( .A(p_input[7096]), .B(p_input[37096]), .Z(n6455) );
  AND U9685 ( .A(n6457), .B(n6458), .Z(o[7095]) );
  AND U9686 ( .A(p_input[27095]), .B(p_input[17095]), .Z(n6458) );
  AND U9687 ( .A(p_input[7095]), .B(p_input[37095]), .Z(n6457) );
  AND U9688 ( .A(n6459), .B(n6460), .Z(o[7094]) );
  AND U9689 ( .A(p_input[27094]), .B(p_input[17094]), .Z(n6460) );
  AND U9690 ( .A(p_input[7094]), .B(p_input[37094]), .Z(n6459) );
  AND U9691 ( .A(n6461), .B(n6462), .Z(o[7093]) );
  AND U9692 ( .A(p_input[27093]), .B(p_input[17093]), .Z(n6462) );
  AND U9693 ( .A(p_input[7093]), .B(p_input[37093]), .Z(n6461) );
  AND U9694 ( .A(n6463), .B(n6464), .Z(o[7092]) );
  AND U9695 ( .A(p_input[27092]), .B(p_input[17092]), .Z(n6464) );
  AND U9696 ( .A(p_input[7092]), .B(p_input[37092]), .Z(n6463) );
  AND U9697 ( .A(n6465), .B(n6466), .Z(o[7091]) );
  AND U9698 ( .A(p_input[27091]), .B(p_input[17091]), .Z(n6466) );
  AND U9699 ( .A(p_input[7091]), .B(p_input[37091]), .Z(n6465) );
  AND U9700 ( .A(n6467), .B(n6468), .Z(o[7090]) );
  AND U9701 ( .A(p_input[27090]), .B(p_input[17090]), .Z(n6468) );
  AND U9702 ( .A(p_input[7090]), .B(p_input[37090]), .Z(n6467) );
  AND U9703 ( .A(n6469), .B(n6470), .Z(o[708]) );
  AND U9704 ( .A(p_input[20708]), .B(p_input[10708]), .Z(n6470) );
  AND U9705 ( .A(p_input[708]), .B(p_input[30708]), .Z(n6469) );
  AND U9706 ( .A(n6471), .B(n6472), .Z(o[7089]) );
  AND U9707 ( .A(p_input[27089]), .B(p_input[17089]), .Z(n6472) );
  AND U9708 ( .A(p_input[7089]), .B(p_input[37089]), .Z(n6471) );
  AND U9709 ( .A(n6473), .B(n6474), .Z(o[7088]) );
  AND U9710 ( .A(p_input[27088]), .B(p_input[17088]), .Z(n6474) );
  AND U9711 ( .A(p_input[7088]), .B(p_input[37088]), .Z(n6473) );
  AND U9712 ( .A(n6475), .B(n6476), .Z(o[7087]) );
  AND U9713 ( .A(p_input[27087]), .B(p_input[17087]), .Z(n6476) );
  AND U9714 ( .A(p_input[7087]), .B(p_input[37087]), .Z(n6475) );
  AND U9715 ( .A(n6477), .B(n6478), .Z(o[7086]) );
  AND U9716 ( .A(p_input[27086]), .B(p_input[17086]), .Z(n6478) );
  AND U9717 ( .A(p_input[7086]), .B(p_input[37086]), .Z(n6477) );
  AND U9718 ( .A(n6479), .B(n6480), .Z(o[7085]) );
  AND U9719 ( .A(p_input[27085]), .B(p_input[17085]), .Z(n6480) );
  AND U9720 ( .A(p_input[7085]), .B(p_input[37085]), .Z(n6479) );
  AND U9721 ( .A(n6481), .B(n6482), .Z(o[7084]) );
  AND U9722 ( .A(p_input[27084]), .B(p_input[17084]), .Z(n6482) );
  AND U9723 ( .A(p_input[7084]), .B(p_input[37084]), .Z(n6481) );
  AND U9724 ( .A(n6483), .B(n6484), .Z(o[7083]) );
  AND U9725 ( .A(p_input[27083]), .B(p_input[17083]), .Z(n6484) );
  AND U9726 ( .A(p_input[7083]), .B(p_input[37083]), .Z(n6483) );
  AND U9727 ( .A(n6485), .B(n6486), .Z(o[7082]) );
  AND U9728 ( .A(p_input[27082]), .B(p_input[17082]), .Z(n6486) );
  AND U9729 ( .A(p_input[7082]), .B(p_input[37082]), .Z(n6485) );
  AND U9730 ( .A(n6487), .B(n6488), .Z(o[7081]) );
  AND U9731 ( .A(p_input[27081]), .B(p_input[17081]), .Z(n6488) );
  AND U9732 ( .A(p_input[7081]), .B(p_input[37081]), .Z(n6487) );
  AND U9733 ( .A(n6489), .B(n6490), .Z(o[7080]) );
  AND U9734 ( .A(p_input[27080]), .B(p_input[17080]), .Z(n6490) );
  AND U9735 ( .A(p_input[7080]), .B(p_input[37080]), .Z(n6489) );
  AND U9736 ( .A(n6491), .B(n6492), .Z(o[707]) );
  AND U9737 ( .A(p_input[20707]), .B(p_input[10707]), .Z(n6492) );
  AND U9738 ( .A(p_input[707]), .B(p_input[30707]), .Z(n6491) );
  AND U9739 ( .A(n6493), .B(n6494), .Z(o[7079]) );
  AND U9740 ( .A(p_input[27079]), .B(p_input[17079]), .Z(n6494) );
  AND U9741 ( .A(p_input[7079]), .B(p_input[37079]), .Z(n6493) );
  AND U9742 ( .A(n6495), .B(n6496), .Z(o[7078]) );
  AND U9743 ( .A(p_input[27078]), .B(p_input[17078]), .Z(n6496) );
  AND U9744 ( .A(p_input[7078]), .B(p_input[37078]), .Z(n6495) );
  AND U9745 ( .A(n6497), .B(n6498), .Z(o[7077]) );
  AND U9746 ( .A(p_input[27077]), .B(p_input[17077]), .Z(n6498) );
  AND U9747 ( .A(p_input[7077]), .B(p_input[37077]), .Z(n6497) );
  AND U9748 ( .A(n6499), .B(n6500), .Z(o[7076]) );
  AND U9749 ( .A(p_input[27076]), .B(p_input[17076]), .Z(n6500) );
  AND U9750 ( .A(p_input[7076]), .B(p_input[37076]), .Z(n6499) );
  AND U9751 ( .A(n6501), .B(n6502), .Z(o[7075]) );
  AND U9752 ( .A(p_input[27075]), .B(p_input[17075]), .Z(n6502) );
  AND U9753 ( .A(p_input[7075]), .B(p_input[37075]), .Z(n6501) );
  AND U9754 ( .A(n6503), .B(n6504), .Z(o[7074]) );
  AND U9755 ( .A(p_input[27074]), .B(p_input[17074]), .Z(n6504) );
  AND U9756 ( .A(p_input[7074]), .B(p_input[37074]), .Z(n6503) );
  AND U9757 ( .A(n6505), .B(n6506), .Z(o[7073]) );
  AND U9758 ( .A(p_input[27073]), .B(p_input[17073]), .Z(n6506) );
  AND U9759 ( .A(p_input[7073]), .B(p_input[37073]), .Z(n6505) );
  AND U9760 ( .A(n6507), .B(n6508), .Z(o[7072]) );
  AND U9761 ( .A(p_input[27072]), .B(p_input[17072]), .Z(n6508) );
  AND U9762 ( .A(p_input[7072]), .B(p_input[37072]), .Z(n6507) );
  AND U9763 ( .A(n6509), .B(n6510), .Z(o[7071]) );
  AND U9764 ( .A(p_input[27071]), .B(p_input[17071]), .Z(n6510) );
  AND U9765 ( .A(p_input[7071]), .B(p_input[37071]), .Z(n6509) );
  AND U9766 ( .A(n6511), .B(n6512), .Z(o[7070]) );
  AND U9767 ( .A(p_input[27070]), .B(p_input[17070]), .Z(n6512) );
  AND U9768 ( .A(p_input[7070]), .B(p_input[37070]), .Z(n6511) );
  AND U9769 ( .A(n6513), .B(n6514), .Z(o[706]) );
  AND U9770 ( .A(p_input[20706]), .B(p_input[10706]), .Z(n6514) );
  AND U9771 ( .A(p_input[706]), .B(p_input[30706]), .Z(n6513) );
  AND U9772 ( .A(n6515), .B(n6516), .Z(o[7069]) );
  AND U9773 ( .A(p_input[27069]), .B(p_input[17069]), .Z(n6516) );
  AND U9774 ( .A(p_input[7069]), .B(p_input[37069]), .Z(n6515) );
  AND U9775 ( .A(n6517), .B(n6518), .Z(o[7068]) );
  AND U9776 ( .A(p_input[27068]), .B(p_input[17068]), .Z(n6518) );
  AND U9777 ( .A(p_input[7068]), .B(p_input[37068]), .Z(n6517) );
  AND U9778 ( .A(n6519), .B(n6520), .Z(o[7067]) );
  AND U9779 ( .A(p_input[27067]), .B(p_input[17067]), .Z(n6520) );
  AND U9780 ( .A(p_input[7067]), .B(p_input[37067]), .Z(n6519) );
  AND U9781 ( .A(n6521), .B(n6522), .Z(o[7066]) );
  AND U9782 ( .A(p_input[27066]), .B(p_input[17066]), .Z(n6522) );
  AND U9783 ( .A(p_input[7066]), .B(p_input[37066]), .Z(n6521) );
  AND U9784 ( .A(n6523), .B(n6524), .Z(o[7065]) );
  AND U9785 ( .A(p_input[27065]), .B(p_input[17065]), .Z(n6524) );
  AND U9786 ( .A(p_input[7065]), .B(p_input[37065]), .Z(n6523) );
  AND U9787 ( .A(n6525), .B(n6526), .Z(o[7064]) );
  AND U9788 ( .A(p_input[27064]), .B(p_input[17064]), .Z(n6526) );
  AND U9789 ( .A(p_input[7064]), .B(p_input[37064]), .Z(n6525) );
  AND U9790 ( .A(n6527), .B(n6528), .Z(o[7063]) );
  AND U9791 ( .A(p_input[27063]), .B(p_input[17063]), .Z(n6528) );
  AND U9792 ( .A(p_input[7063]), .B(p_input[37063]), .Z(n6527) );
  AND U9793 ( .A(n6529), .B(n6530), .Z(o[7062]) );
  AND U9794 ( .A(p_input[27062]), .B(p_input[17062]), .Z(n6530) );
  AND U9795 ( .A(p_input[7062]), .B(p_input[37062]), .Z(n6529) );
  AND U9796 ( .A(n6531), .B(n6532), .Z(o[7061]) );
  AND U9797 ( .A(p_input[27061]), .B(p_input[17061]), .Z(n6532) );
  AND U9798 ( .A(p_input[7061]), .B(p_input[37061]), .Z(n6531) );
  AND U9799 ( .A(n6533), .B(n6534), .Z(o[7060]) );
  AND U9800 ( .A(p_input[27060]), .B(p_input[17060]), .Z(n6534) );
  AND U9801 ( .A(p_input[7060]), .B(p_input[37060]), .Z(n6533) );
  AND U9802 ( .A(n6535), .B(n6536), .Z(o[705]) );
  AND U9803 ( .A(p_input[20705]), .B(p_input[10705]), .Z(n6536) );
  AND U9804 ( .A(p_input[705]), .B(p_input[30705]), .Z(n6535) );
  AND U9805 ( .A(n6537), .B(n6538), .Z(o[7059]) );
  AND U9806 ( .A(p_input[27059]), .B(p_input[17059]), .Z(n6538) );
  AND U9807 ( .A(p_input[7059]), .B(p_input[37059]), .Z(n6537) );
  AND U9808 ( .A(n6539), .B(n6540), .Z(o[7058]) );
  AND U9809 ( .A(p_input[27058]), .B(p_input[17058]), .Z(n6540) );
  AND U9810 ( .A(p_input[7058]), .B(p_input[37058]), .Z(n6539) );
  AND U9811 ( .A(n6541), .B(n6542), .Z(o[7057]) );
  AND U9812 ( .A(p_input[27057]), .B(p_input[17057]), .Z(n6542) );
  AND U9813 ( .A(p_input[7057]), .B(p_input[37057]), .Z(n6541) );
  AND U9814 ( .A(n6543), .B(n6544), .Z(o[7056]) );
  AND U9815 ( .A(p_input[27056]), .B(p_input[17056]), .Z(n6544) );
  AND U9816 ( .A(p_input[7056]), .B(p_input[37056]), .Z(n6543) );
  AND U9817 ( .A(n6545), .B(n6546), .Z(o[7055]) );
  AND U9818 ( .A(p_input[27055]), .B(p_input[17055]), .Z(n6546) );
  AND U9819 ( .A(p_input[7055]), .B(p_input[37055]), .Z(n6545) );
  AND U9820 ( .A(n6547), .B(n6548), .Z(o[7054]) );
  AND U9821 ( .A(p_input[27054]), .B(p_input[17054]), .Z(n6548) );
  AND U9822 ( .A(p_input[7054]), .B(p_input[37054]), .Z(n6547) );
  AND U9823 ( .A(n6549), .B(n6550), .Z(o[7053]) );
  AND U9824 ( .A(p_input[27053]), .B(p_input[17053]), .Z(n6550) );
  AND U9825 ( .A(p_input[7053]), .B(p_input[37053]), .Z(n6549) );
  AND U9826 ( .A(n6551), .B(n6552), .Z(o[7052]) );
  AND U9827 ( .A(p_input[27052]), .B(p_input[17052]), .Z(n6552) );
  AND U9828 ( .A(p_input[7052]), .B(p_input[37052]), .Z(n6551) );
  AND U9829 ( .A(n6553), .B(n6554), .Z(o[7051]) );
  AND U9830 ( .A(p_input[27051]), .B(p_input[17051]), .Z(n6554) );
  AND U9831 ( .A(p_input[7051]), .B(p_input[37051]), .Z(n6553) );
  AND U9832 ( .A(n6555), .B(n6556), .Z(o[7050]) );
  AND U9833 ( .A(p_input[27050]), .B(p_input[17050]), .Z(n6556) );
  AND U9834 ( .A(p_input[7050]), .B(p_input[37050]), .Z(n6555) );
  AND U9835 ( .A(n6557), .B(n6558), .Z(o[704]) );
  AND U9836 ( .A(p_input[20704]), .B(p_input[10704]), .Z(n6558) );
  AND U9837 ( .A(p_input[704]), .B(p_input[30704]), .Z(n6557) );
  AND U9838 ( .A(n6559), .B(n6560), .Z(o[7049]) );
  AND U9839 ( .A(p_input[27049]), .B(p_input[17049]), .Z(n6560) );
  AND U9840 ( .A(p_input[7049]), .B(p_input[37049]), .Z(n6559) );
  AND U9841 ( .A(n6561), .B(n6562), .Z(o[7048]) );
  AND U9842 ( .A(p_input[27048]), .B(p_input[17048]), .Z(n6562) );
  AND U9843 ( .A(p_input[7048]), .B(p_input[37048]), .Z(n6561) );
  AND U9844 ( .A(n6563), .B(n6564), .Z(o[7047]) );
  AND U9845 ( .A(p_input[27047]), .B(p_input[17047]), .Z(n6564) );
  AND U9846 ( .A(p_input[7047]), .B(p_input[37047]), .Z(n6563) );
  AND U9847 ( .A(n6565), .B(n6566), .Z(o[7046]) );
  AND U9848 ( .A(p_input[27046]), .B(p_input[17046]), .Z(n6566) );
  AND U9849 ( .A(p_input[7046]), .B(p_input[37046]), .Z(n6565) );
  AND U9850 ( .A(n6567), .B(n6568), .Z(o[7045]) );
  AND U9851 ( .A(p_input[27045]), .B(p_input[17045]), .Z(n6568) );
  AND U9852 ( .A(p_input[7045]), .B(p_input[37045]), .Z(n6567) );
  AND U9853 ( .A(n6569), .B(n6570), .Z(o[7044]) );
  AND U9854 ( .A(p_input[27044]), .B(p_input[17044]), .Z(n6570) );
  AND U9855 ( .A(p_input[7044]), .B(p_input[37044]), .Z(n6569) );
  AND U9856 ( .A(n6571), .B(n6572), .Z(o[7043]) );
  AND U9857 ( .A(p_input[27043]), .B(p_input[17043]), .Z(n6572) );
  AND U9858 ( .A(p_input[7043]), .B(p_input[37043]), .Z(n6571) );
  AND U9859 ( .A(n6573), .B(n6574), .Z(o[7042]) );
  AND U9860 ( .A(p_input[27042]), .B(p_input[17042]), .Z(n6574) );
  AND U9861 ( .A(p_input[7042]), .B(p_input[37042]), .Z(n6573) );
  AND U9862 ( .A(n6575), .B(n6576), .Z(o[7041]) );
  AND U9863 ( .A(p_input[27041]), .B(p_input[17041]), .Z(n6576) );
  AND U9864 ( .A(p_input[7041]), .B(p_input[37041]), .Z(n6575) );
  AND U9865 ( .A(n6577), .B(n6578), .Z(o[7040]) );
  AND U9866 ( .A(p_input[27040]), .B(p_input[17040]), .Z(n6578) );
  AND U9867 ( .A(p_input[7040]), .B(p_input[37040]), .Z(n6577) );
  AND U9868 ( .A(n6579), .B(n6580), .Z(o[703]) );
  AND U9869 ( .A(p_input[20703]), .B(p_input[10703]), .Z(n6580) );
  AND U9870 ( .A(p_input[703]), .B(p_input[30703]), .Z(n6579) );
  AND U9871 ( .A(n6581), .B(n6582), .Z(o[7039]) );
  AND U9872 ( .A(p_input[27039]), .B(p_input[17039]), .Z(n6582) );
  AND U9873 ( .A(p_input[7039]), .B(p_input[37039]), .Z(n6581) );
  AND U9874 ( .A(n6583), .B(n6584), .Z(o[7038]) );
  AND U9875 ( .A(p_input[27038]), .B(p_input[17038]), .Z(n6584) );
  AND U9876 ( .A(p_input[7038]), .B(p_input[37038]), .Z(n6583) );
  AND U9877 ( .A(n6585), .B(n6586), .Z(o[7037]) );
  AND U9878 ( .A(p_input[27037]), .B(p_input[17037]), .Z(n6586) );
  AND U9879 ( .A(p_input[7037]), .B(p_input[37037]), .Z(n6585) );
  AND U9880 ( .A(n6587), .B(n6588), .Z(o[7036]) );
  AND U9881 ( .A(p_input[27036]), .B(p_input[17036]), .Z(n6588) );
  AND U9882 ( .A(p_input[7036]), .B(p_input[37036]), .Z(n6587) );
  AND U9883 ( .A(n6589), .B(n6590), .Z(o[7035]) );
  AND U9884 ( .A(p_input[27035]), .B(p_input[17035]), .Z(n6590) );
  AND U9885 ( .A(p_input[7035]), .B(p_input[37035]), .Z(n6589) );
  AND U9886 ( .A(n6591), .B(n6592), .Z(o[7034]) );
  AND U9887 ( .A(p_input[27034]), .B(p_input[17034]), .Z(n6592) );
  AND U9888 ( .A(p_input[7034]), .B(p_input[37034]), .Z(n6591) );
  AND U9889 ( .A(n6593), .B(n6594), .Z(o[7033]) );
  AND U9890 ( .A(p_input[27033]), .B(p_input[17033]), .Z(n6594) );
  AND U9891 ( .A(p_input[7033]), .B(p_input[37033]), .Z(n6593) );
  AND U9892 ( .A(n6595), .B(n6596), .Z(o[7032]) );
  AND U9893 ( .A(p_input[27032]), .B(p_input[17032]), .Z(n6596) );
  AND U9894 ( .A(p_input[7032]), .B(p_input[37032]), .Z(n6595) );
  AND U9895 ( .A(n6597), .B(n6598), .Z(o[7031]) );
  AND U9896 ( .A(p_input[27031]), .B(p_input[17031]), .Z(n6598) );
  AND U9897 ( .A(p_input[7031]), .B(p_input[37031]), .Z(n6597) );
  AND U9898 ( .A(n6599), .B(n6600), .Z(o[7030]) );
  AND U9899 ( .A(p_input[27030]), .B(p_input[17030]), .Z(n6600) );
  AND U9900 ( .A(p_input[7030]), .B(p_input[37030]), .Z(n6599) );
  AND U9901 ( .A(n6601), .B(n6602), .Z(o[702]) );
  AND U9902 ( .A(p_input[20702]), .B(p_input[10702]), .Z(n6602) );
  AND U9903 ( .A(p_input[702]), .B(p_input[30702]), .Z(n6601) );
  AND U9904 ( .A(n6603), .B(n6604), .Z(o[7029]) );
  AND U9905 ( .A(p_input[27029]), .B(p_input[17029]), .Z(n6604) );
  AND U9906 ( .A(p_input[7029]), .B(p_input[37029]), .Z(n6603) );
  AND U9907 ( .A(n6605), .B(n6606), .Z(o[7028]) );
  AND U9908 ( .A(p_input[27028]), .B(p_input[17028]), .Z(n6606) );
  AND U9909 ( .A(p_input[7028]), .B(p_input[37028]), .Z(n6605) );
  AND U9910 ( .A(n6607), .B(n6608), .Z(o[7027]) );
  AND U9911 ( .A(p_input[27027]), .B(p_input[17027]), .Z(n6608) );
  AND U9912 ( .A(p_input[7027]), .B(p_input[37027]), .Z(n6607) );
  AND U9913 ( .A(n6609), .B(n6610), .Z(o[7026]) );
  AND U9914 ( .A(p_input[27026]), .B(p_input[17026]), .Z(n6610) );
  AND U9915 ( .A(p_input[7026]), .B(p_input[37026]), .Z(n6609) );
  AND U9916 ( .A(n6611), .B(n6612), .Z(o[7025]) );
  AND U9917 ( .A(p_input[27025]), .B(p_input[17025]), .Z(n6612) );
  AND U9918 ( .A(p_input[7025]), .B(p_input[37025]), .Z(n6611) );
  AND U9919 ( .A(n6613), .B(n6614), .Z(o[7024]) );
  AND U9920 ( .A(p_input[27024]), .B(p_input[17024]), .Z(n6614) );
  AND U9921 ( .A(p_input[7024]), .B(p_input[37024]), .Z(n6613) );
  AND U9922 ( .A(n6615), .B(n6616), .Z(o[7023]) );
  AND U9923 ( .A(p_input[27023]), .B(p_input[17023]), .Z(n6616) );
  AND U9924 ( .A(p_input[7023]), .B(p_input[37023]), .Z(n6615) );
  AND U9925 ( .A(n6617), .B(n6618), .Z(o[7022]) );
  AND U9926 ( .A(p_input[27022]), .B(p_input[17022]), .Z(n6618) );
  AND U9927 ( .A(p_input[7022]), .B(p_input[37022]), .Z(n6617) );
  AND U9928 ( .A(n6619), .B(n6620), .Z(o[7021]) );
  AND U9929 ( .A(p_input[27021]), .B(p_input[17021]), .Z(n6620) );
  AND U9930 ( .A(p_input[7021]), .B(p_input[37021]), .Z(n6619) );
  AND U9931 ( .A(n6621), .B(n6622), .Z(o[7020]) );
  AND U9932 ( .A(p_input[27020]), .B(p_input[17020]), .Z(n6622) );
  AND U9933 ( .A(p_input[7020]), .B(p_input[37020]), .Z(n6621) );
  AND U9934 ( .A(n6623), .B(n6624), .Z(o[701]) );
  AND U9935 ( .A(p_input[20701]), .B(p_input[10701]), .Z(n6624) );
  AND U9936 ( .A(p_input[701]), .B(p_input[30701]), .Z(n6623) );
  AND U9937 ( .A(n6625), .B(n6626), .Z(o[7019]) );
  AND U9938 ( .A(p_input[27019]), .B(p_input[17019]), .Z(n6626) );
  AND U9939 ( .A(p_input[7019]), .B(p_input[37019]), .Z(n6625) );
  AND U9940 ( .A(n6627), .B(n6628), .Z(o[7018]) );
  AND U9941 ( .A(p_input[27018]), .B(p_input[17018]), .Z(n6628) );
  AND U9942 ( .A(p_input[7018]), .B(p_input[37018]), .Z(n6627) );
  AND U9943 ( .A(n6629), .B(n6630), .Z(o[7017]) );
  AND U9944 ( .A(p_input[27017]), .B(p_input[17017]), .Z(n6630) );
  AND U9945 ( .A(p_input[7017]), .B(p_input[37017]), .Z(n6629) );
  AND U9946 ( .A(n6631), .B(n6632), .Z(o[7016]) );
  AND U9947 ( .A(p_input[27016]), .B(p_input[17016]), .Z(n6632) );
  AND U9948 ( .A(p_input[7016]), .B(p_input[37016]), .Z(n6631) );
  AND U9949 ( .A(n6633), .B(n6634), .Z(o[7015]) );
  AND U9950 ( .A(p_input[27015]), .B(p_input[17015]), .Z(n6634) );
  AND U9951 ( .A(p_input[7015]), .B(p_input[37015]), .Z(n6633) );
  AND U9952 ( .A(n6635), .B(n6636), .Z(o[7014]) );
  AND U9953 ( .A(p_input[27014]), .B(p_input[17014]), .Z(n6636) );
  AND U9954 ( .A(p_input[7014]), .B(p_input[37014]), .Z(n6635) );
  AND U9955 ( .A(n6637), .B(n6638), .Z(o[7013]) );
  AND U9956 ( .A(p_input[27013]), .B(p_input[17013]), .Z(n6638) );
  AND U9957 ( .A(p_input[7013]), .B(p_input[37013]), .Z(n6637) );
  AND U9958 ( .A(n6639), .B(n6640), .Z(o[7012]) );
  AND U9959 ( .A(p_input[27012]), .B(p_input[17012]), .Z(n6640) );
  AND U9960 ( .A(p_input[7012]), .B(p_input[37012]), .Z(n6639) );
  AND U9961 ( .A(n6641), .B(n6642), .Z(o[7011]) );
  AND U9962 ( .A(p_input[27011]), .B(p_input[17011]), .Z(n6642) );
  AND U9963 ( .A(p_input[7011]), .B(p_input[37011]), .Z(n6641) );
  AND U9964 ( .A(n6643), .B(n6644), .Z(o[7010]) );
  AND U9965 ( .A(p_input[27010]), .B(p_input[17010]), .Z(n6644) );
  AND U9966 ( .A(p_input[7010]), .B(p_input[37010]), .Z(n6643) );
  AND U9967 ( .A(n6645), .B(n6646), .Z(o[700]) );
  AND U9968 ( .A(p_input[20700]), .B(p_input[10700]), .Z(n6646) );
  AND U9969 ( .A(p_input[700]), .B(p_input[30700]), .Z(n6645) );
  AND U9970 ( .A(n6647), .B(n6648), .Z(o[7009]) );
  AND U9971 ( .A(p_input[27009]), .B(p_input[17009]), .Z(n6648) );
  AND U9972 ( .A(p_input[7009]), .B(p_input[37009]), .Z(n6647) );
  AND U9973 ( .A(n6649), .B(n6650), .Z(o[7008]) );
  AND U9974 ( .A(p_input[27008]), .B(p_input[17008]), .Z(n6650) );
  AND U9975 ( .A(p_input[7008]), .B(p_input[37008]), .Z(n6649) );
  AND U9976 ( .A(n6651), .B(n6652), .Z(o[7007]) );
  AND U9977 ( .A(p_input[27007]), .B(p_input[17007]), .Z(n6652) );
  AND U9978 ( .A(p_input[7007]), .B(p_input[37007]), .Z(n6651) );
  AND U9979 ( .A(n6653), .B(n6654), .Z(o[7006]) );
  AND U9980 ( .A(p_input[27006]), .B(p_input[17006]), .Z(n6654) );
  AND U9981 ( .A(p_input[7006]), .B(p_input[37006]), .Z(n6653) );
  AND U9982 ( .A(n6655), .B(n6656), .Z(o[7005]) );
  AND U9983 ( .A(p_input[27005]), .B(p_input[17005]), .Z(n6656) );
  AND U9984 ( .A(p_input[7005]), .B(p_input[37005]), .Z(n6655) );
  AND U9985 ( .A(n6657), .B(n6658), .Z(o[7004]) );
  AND U9986 ( .A(p_input[27004]), .B(p_input[17004]), .Z(n6658) );
  AND U9987 ( .A(p_input[7004]), .B(p_input[37004]), .Z(n6657) );
  AND U9988 ( .A(n6659), .B(n6660), .Z(o[7003]) );
  AND U9989 ( .A(p_input[27003]), .B(p_input[17003]), .Z(n6660) );
  AND U9990 ( .A(p_input[7003]), .B(p_input[37003]), .Z(n6659) );
  AND U9991 ( .A(n6661), .B(n6662), .Z(o[7002]) );
  AND U9992 ( .A(p_input[27002]), .B(p_input[17002]), .Z(n6662) );
  AND U9993 ( .A(p_input[7002]), .B(p_input[37002]), .Z(n6661) );
  AND U9994 ( .A(n6663), .B(n6664), .Z(o[7001]) );
  AND U9995 ( .A(p_input[27001]), .B(p_input[17001]), .Z(n6664) );
  AND U9996 ( .A(p_input[7001]), .B(p_input[37001]), .Z(n6663) );
  AND U9997 ( .A(n6665), .B(n6666), .Z(o[7000]) );
  AND U9998 ( .A(p_input[27000]), .B(p_input[17000]), .Z(n6666) );
  AND U9999 ( .A(p_input[7000]), .B(p_input[37000]), .Z(n6665) );
  AND U10000 ( .A(n6667), .B(n6668), .Z(o[6]) );
  AND U10001 ( .A(p_input[20006]), .B(p_input[10006]), .Z(n6668) );
  AND U10002 ( .A(p_input[6]), .B(p_input[30006]), .Z(n6667) );
  AND U10003 ( .A(n6669), .B(n6670), .Z(o[69]) );
  AND U10004 ( .A(p_input[20069]), .B(p_input[10069]), .Z(n6670) );
  AND U10005 ( .A(p_input[69]), .B(p_input[30069]), .Z(n6669) );
  AND U10006 ( .A(n6671), .B(n6672), .Z(o[699]) );
  AND U10007 ( .A(p_input[20699]), .B(p_input[10699]), .Z(n6672) );
  AND U10008 ( .A(p_input[699]), .B(p_input[30699]), .Z(n6671) );
  AND U10009 ( .A(n6673), .B(n6674), .Z(o[6999]) );
  AND U10010 ( .A(p_input[26999]), .B(p_input[16999]), .Z(n6674) );
  AND U10011 ( .A(p_input[6999]), .B(p_input[36999]), .Z(n6673) );
  AND U10012 ( .A(n6675), .B(n6676), .Z(o[6998]) );
  AND U10013 ( .A(p_input[26998]), .B(p_input[16998]), .Z(n6676) );
  AND U10014 ( .A(p_input[6998]), .B(p_input[36998]), .Z(n6675) );
  AND U10015 ( .A(n6677), .B(n6678), .Z(o[6997]) );
  AND U10016 ( .A(p_input[26997]), .B(p_input[16997]), .Z(n6678) );
  AND U10017 ( .A(p_input[6997]), .B(p_input[36997]), .Z(n6677) );
  AND U10018 ( .A(n6679), .B(n6680), .Z(o[6996]) );
  AND U10019 ( .A(p_input[26996]), .B(p_input[16996]), .Z(n6680) );
  AND U10020 ( .A(p_input[6996]), .B(p_input[36996]), .Z(n6679) );
  AND U10021 ( .A(n6681), .B(n6682), .Z(o[6995]) );
  AND U10022 ( .A(p_input[26995]), .B(p_input[16995]), .Z(n6682) );
  AND U10023 ( .A(p_input[6995]), .B(p_input[36995]), .Z(n6681) );
  AND U10024 ( .A(n6683), .B(n6684), .Z(o[6994]) );
  AND U10025 ( .A(p_input[26994]), .B(p_input[16994]), .Z(n6684) );
  AND U10026 ( .A(p_input[6994]), .B(p_input[36994]), .Z(n6683) );
  AND U10027 ( .A(n6685), .B(n6686), .Z(o[6993]) );
  AND U10028 ( .A(p_input[26993]), .B(p_input[16993]), .Z(n6686) );
  AND U10029 ( .A(p_input[6993]), .B(p_input[36993]), .Z(n6685) );
  AND U10030 ( .A(n6687), .B(n6688), .Z(o[6992]) );
  AND U10031 ( .A(p_input[26992]), .B(p_input[16992]), .Z(n6688) );
  AND U10032 ( .A(p_input[6992]), .B(p_input[36992]), .Z(n6687) );
  AND U10033 ( .A(n6689), .B(n6690), .Z(o[6991]) );
  AND U10034 ( .A(p_input[26991]), .B(p_input[16991]), .Z(n6690) );
  AND U10035 ( .A(p_input[6991]), .B(p_input[36991]), .Z(n6689) );
  AND U10036 ( .A(n6691), .B(n6692), .Z(o[6990]) );
  AND U10037 ( .A(p_input[26990]), .B(p_input[16990]), .Z(n6692) );
  AND U10038 ( .A(p_input[6990]), .B(p_input[36990]), .Z(n6691) );
  AND U10039 ( .A(n6693), .B(n6694), .Z(o[698]) );
  AND U10040 ( .A(p_input[20698]), .B(p_input[10698]), .Z(n6694) );
  AND U10041 ( .A(p_input[698]), .B(p_input[30698]), .Z(n6693) );
  AND U10042 ( .A(n6695), .B(n6696), .Z(o[6989]) );
  AND U10043 ( .A(p_input[26989]), .B(p_input[16989]), .Z(n6696) );
  AND U10044 ( .A(p_input[6989]), .B(p_input[36989]), .Z(n6695) );
  AND U10045 ( .A(n6697), .B(n6698), .Z(o[6988]) );
  AND U10046 ( .A(p_input[26988]), .B(p_input[16988]), .Z(n6698) );
  AND U10047 ( .A(p_input[6988]), .B(p_input[36988]), .Z(n6697) );
  AND U10048 ( .A(n6699), .B(n6700), .Z(o[6987]) );
  AND U10049 ( .A(p_input[26987]), .B(p_input[16987]), .Z(n6700) );
  AND U10050 ( .A(p_input[6987]), .B(p_input[36987]), .Z(n6699) );
  AND U10051 ( .A(n6701), .B(n6702), .Z(o[6986]) );
  AND U10052 ( .A(p_input[26986]), .B(p_input[16986]), .Z(n6702) );
  AND U10053 ( .A(p_input[6986]), .B(p_input[36986]), .Z(n6701) );
  AND U10054 ( .A(n6703), .B(n6704), .Z(o[6985]) );
  AND U10055 ( .A(p_input[26985]), .B(p_input[16985]), .Z(n6704) );
  AND U10056 ( .A(p_input[6985]), .B(p_input[36985]), .Z(n6703) );
  AND U10057 ( .A(n6705), .B(n6706), .Z(o[6984]) );
  AND U10058 ( .A(p_input[26984]), .B(p_input[16984]), .Z(n6706) );
  AND U10059 ( .A(p_input[6984]), .B(p_input[36984]), .Z(n6705) );
  AND U10060 ( .A(n6707), .B(n6708), .Z(o[6983]) );
  AND U10061 ( .A(p_input[26983]), .B(p_input[16983]), .Z(n6708) );
  AND U10062 ( .A(p_input[6983]), .B(p_input[36983]), .Z(n6707) );
  AND U10063 ( .A(n6709), .B(n6710), .Z(o[6982]) );
  AND U10064 ( .A(p_input[26982]), .B(p_input[16982]), .Z(n6710) );
  AND U10065 ( .A(p_input[6982]), .B(p_input[36982]), .Z(n6709) );
  AND U10066 ( .A(n6711), .B(n6712), .Z(o[6981]) );
  AND U10067 ( .A(p_input[26981]), .B(p_input[16981]), .Z(n6712) );
  AND U10068 ( .A(p_input[6981]), .B(p_input[36981]), .Z(n6711) );
  AND U10069 ( .A(n6713), .B(n6714), .Z(o[6980]) );
  AND U10070 ( .A(p_input[26980]), .B(p_input[16980]), .Z(n6714) );
  AND U10071 ( .A(p_input[6980]), .B(p_input[36980]), .Z(n6713) );
  AND U10072 ( .A(n6715), .B(n6716), .Z(o[697]) );
  AND U10073 ( .A(p_input[20697]), .B(p_input[10697]), .Z(n6716) );
  AND U10074 ( .A(p_input[697]), .B(p_input[30697]), .Z(n6715) );
  AND U10075 ( .A(n6717), .B(n6718), .Z(o[6979]) );
  AND U10076 ( .A(p_input[26979]), .B(p_input[16979]), .Z(n6718) );
  AND U10077 ( .A(p_input[6979]), .B(p_input[36979]), .Z(n6717) );
  AND U10078 ( .A(n6719), .B(n6720), .Z(o[6978]) );
  AND U10079 ( .A(p_input[26978]), .B(p_input[16978]), .Z(n6720) );
  AND U10080 ( .A(p_input[6978]), .B(p_input[36978]), .Z(n6719) );
  AND U10081 ( .A(n6721), .B(n6722), .Z(o[6977]) );
  AND U10082 ( .A(p_input[26977]), .B(p_input[16977]), .Z(n6722) );
  AND U10083 ( .A(p_input[6977]), .B(p_input[36977]), .Z(n6721) );
  AND U10084 ( .A(n6723), .B(n6724), .Z(o[6976]) );
  AND U10085 ( .A(p_input[26976]), .B(p_input[16976]), .Z(n6724) );
  AND U10086 ( .A(p_input[6976]), .B(p_input[36976]), .Z(n6723) );
  AND U10087 ( .A(n6725), .B(n6726), .Z(o[6975]) );
  AND U10088 ( .A(p_input[26975]), .B(p_input[16975]), .Z(n6726) );
  AND U10089 ( .A(p_input[6975]), .B(p_input[36975]), .Z(n6725) );
  AND U10090 ( .A(n6727), .B(n6728), .Z(o[6974]) );
  AND U10091 ( .A(p_input[26974]), .B(p_input[16974]), .Z(n6728) );
  AND U10092 ( .A(p_input[6974]), .B(p_input[36974]), .Z(n6727) );
  AND U10093 ( .A(n6729), .B(n6730), .Z(o[6973]) );
  AND U10094 ( .A(p_input[26973]), .B(p_input[16973]), .Z(n6730) );
  AND U10095 ( .A(p_input[6973]), .B(p_input[36973]), .Z(n6729) );
  AND U10096 ( .A(n6731), .B(n6732), .Z(o[6972]) );
  AND U10097 ( .A(p_input[26972]), .B(p_input[16972]), .Z(n6732) );
  AND U10098 ( .A(p_input[6972]), .B(p_input[36972]), .Z(n6731) );
  AND U10099 ( .A(n6733), .B(n6734), .Z(o[6971]) );
  AND U10100 ( .A(p_input[26971]), .B(p_input[16971]), .Z(n6734) );
  AND U10101 ( .A(p_input[6971]), .B(p_input[36971]), .Z(n6733) );
  AND U10102 ( .A(n6735), .B(n6736), .Z(o[6970]) );
  AND U10103 ( .A(p_input[26970]), .B(p_input[16970]), .Z(n6736) );
  AND U10104 ( .A(p_input[6970]), .B(p_input[36970]), .Z(n6735) );
  AND U10105 ( .A(n6737), .B(n6738), .Z(o[696]) );
  AND U10106 ( .A(p_input[20696]), .B(p_input[10696]), .Z(n6738) );
  AND U10107 ( .A(p_input[696]), .B(p_input[30696]), .Z(n6737) );
  AND U10108 ( .A(n6739), .B(n6740), .Z(o[6969]) );
  AND U10109 ( .A(p_input[26969]), .B(p_input[16969]), .Z(n6740) );
  AND U10110 ( .A(p_input[6969]), .B(p_input[36969]), .Z(n6739) );
  AND U10111 ( .A(n6741), .B(n6742), .Z(o[6968]) );
  AND U10112 ( .A(p_input[26968]), .B(p_input[16968]), .Z(n6742) );
  AND U10113 ( .A(p_input[6968]), .B(p_input[36968]), .Z(n6741) );
  AND U10114 ( .A(n6743), .B(n6744), .Z(o[6967]) );
  AND U10115 ( .A(p_input[26967]), .B(p_input[16967]), .Z(n6744) );
  AND U10116 ( .A(p_input[6967]), .B(p_input[36967]), .Z(n6743) );
  AND U10117 ( .A(n6745), .B(n6746), .Z(o[6966]) );
  AND U10118 ( .A(p_input[26966]), .B(p_input[16966]), .Z(n6746) );
  AND U10119 ( .A(p_input[6966]), .B(p_input[36966]), .Z(n6745) );
  AND U10120 ( .A(n6747), .B(n6748), .Z(o[6965]) );
  AND U10121 ( .A(p_input[26965]), .B(p_input[16965]), .Z(n6748) );
  AND U10122 ( .A(p_input[6965]), .B(p_input[36965]), .Z(n6747) );
  AND U10123 ( .A(n6749), .B(n6750), .Z(o[6964]) );
  AND U10124 ( .A(p_input[26964]), .B(p_input[16964]), .Z(n6750) );
  AND U10125 ( .A(p_input[6964]), .B(p_input[36964]), .Z(n6749) );
  AND U10126 ( .A(n6751), .B(n6752), .Z(o[6963]) );
  AND U10127 ( .A(p_input[26963]), .B(p_input[16963]), .Z(n6752) );
  AND U10128 ( .A(p_input[6963]), .B(p_input[36963]), .Z(n6751) );
  AND U10129 ( .A(n6753), .B(n6754), .Z(o[6962]) );
  AND U10130 ( .A(p_input[26962]), .B(p_input[16962]), .Z(n6754) );
  AND U10131 ( .A(p_input[6962]), .B(p_input[36962]), .Z(n6753) );
  AND U10132 ( .A(n6755), .B(n6756), .Z(o[6961]) );
  AND U10133 ( .A(p_input[26961]), .B(p_input[16961]), .Z(n6756) );
  AND U10134 ( .A(p_input[6961]), .B(p_input[36961]), .Z(n6755) );
  AND U10135 ( .A(n6757), .B(n6758), .Z(o[6960]) );
  AND U10136 ( .A(p_input[26960]), .B(p_input[16960]), .Z(n6758) );
  AND U10137 ( .A(p_input[6960]), .B(p_input[36960]), .Z(n6757) );
  AND U10138 ( .A(n6759), .B(n6760), .Z(o[695]) );
  AND U10139 ( .A(p_input[20695]), .B(p_input[10695]), .Z(n6760) );
  AND U10140 ( .A(p_input[695]), .B(p_input[30695]), .Z(n6759) );
  AND U10141 ( .A(n6761), .B(n6762), .Z(o[6959]) );
  AND U10142 ( .A(p_input[26959]), .B(p_input[16959]), .Z(n6762) );
  AND U10143 ( .A(p_input[6959]), .B(p_input[36959]), .Z(n6761) );
  AND U10144 ( .A(n6763), .B(n6764), .Z(o[6958]) );
  AND U10145 ( .A(p_input[26958]), .B(p_input[16958]), .Z(n6764) );
  AND U10146 ( .A(p_input[6958]), .B(p_input[36958]), .Z(n6763) );
  AND U10147 ( .A(n6765), .B(n6766), .Z(o[6957]) );
  AND U10148 ( .A(p_input[26957]), .B(p_input[16957]), .Z(n6766) );
  AND U10149 ( .A(p_input[6957]), .B(p_input[36957]), .Z(n6765) );
  AND U10150 ( .A(n6767), .B(n6768), .Z(o[6956]) );
  AND U10151 ( .A(p_input[26956]), .B(p_input[16956]), .Z(n6768) );
  AND U10152 ( .A(p_input[6956]), .B(p_input[36956]), .Z(n6767) );
  AND U10153 ( .A(n6769), .B(n6770), .Z(o[6955]) );
  AND U10154 ( .A(p_input[26955]), .B(p_input[16955]), .Z(n6770) );
  AND U10155 ( .A(p_input[6955]), .B(p_input[36955]), .Z(n6769) );
  AND U10156 ( .A(n6771), .B(n6772), .Z(o[6954]) );
  AND U10157 ( .A(p_input[26954]), .B(p_input[16954]), .Z(n6772) );
  AND U10158 ( .A(p_input[6954]), .B(p_input[36954]), .Z(n6771) );
  AND U10159 ( .A(n6773), .B(n6774), .Z(o[6953]) );
  AND U10160 ( .A(p_input[26953]), .B(p_input[16953]), .Z(n6774) );
  AND U10161 ( .A(p_input[6953]), .B(p_input[36953]), .Z(n6773) );
  AND U10162 ( .A(n6775), .B(n6776), .Z(o[6952]) );
  AND U10163 ( .A(p_input[26952]), .B(p_input[16952]), .Z(n6776) );
  AND U10164 ( .A(p_input[6952]), .B(p_input[36952]), .Z(n6775) );
  AND U10165 ( .A(n6777), .B(n6778), .Z(o[6951]) );
  AND U10166 ( .A(p_input[26951]), .B(p_input[16951]), .Z(n6778) );
  AND U10167 ( .A(p_input[6951]), .B(p_input[36951]), .Z(n6777) );
  AND U10168 ( .A(n6779), .B(n6780), .Z(o[6950]) );
  AND U10169 ( .A(p_input[26950]), .B(p_input[16950]), .Z(n6780) );
  AND U10170 ( .A(p_input[6950]), .B(p_input[36950]), .Z(n6779) );
  AND U10171 ( .A(n6781), .B(n6782), .Z(o[694]) );
  AND U10172 ( .A(p_input[20694]), .B(p_input[10694]), .Z(n6782) );
  AND U10173 ( .A(p_input[694]), .B(p_input[30694]), .Z(n6781) );
  AND U10174 ( .A(n6783), .B(n6784), .Z(o[6949]) );
  AND U10175 ( .A(p_input[26949]), .B(p_input[16949]), .Z(n6784) );
  AND U10176 ( .A(p_input[6949]), .B(p_input[36949]), .Z(n6783) );
  AND U10177 ( .A(n6785), .B(n6786), .Z(o[6948]) );
  AND U10178 ( .A(p_input[26948]), .B(p_input[16948]), .Z(n6786) );
  AND U10179 ( .A(p_input[6948]), .B(p_input[36948]), .Z(n6785) );
  AND U10180 ( .A(n6787), .B(n6788), .Z(o[6947]) );
  AND U10181 ( .A(p_input[26947]), .B(p_input[16947]), .Z(n6788) );
  AND U10182 ( .A(p_input[6947]), .B(p_input[36947]), .Z(n6787) );
  AND U10183 ( .A(n6789), .B(n6790), .Z(o[6946]) );
  AND U10184 ( .A(p_input[26946]), .B(p_input[16946]), .Z(n6790) );
  AND U10185 ( .A(p_input[6946]), .B(p_input[36946]), .Z(n6789) );
  AND U10186 ( .A(n6791), .B(n6792), .Z(o[6945]) );
  AND U10187 ( .A(p_input[26945]), .B(p_input[16945]), .Z(n6792) );
  AND U10188 ( .A(p_input[6945]), .B(p_input[36945]), .Z(n6791) );
  AND U10189 ( .A(n6793), .B(n6794), .Z(o[6944]) );
  AND U10190 ( .A(p_input[26944]), .B(p_input[16944]), .Z(n6794) );
  AND U10191 ( .A(p_input[6944]), .B(p_input[36944]), .Z(n6793) );
  AND U10192 ( .A(n6795), .B(n6796), .Z(o[6943]) );
  AND U10193 ( .A(p_input[26943]), .B(p_input[16943]), .Z(n6796) );
  AND U10194 ( .A(p_input[6943]), .B(p_input[36943]), .Z(n6795) );
  AND U10195 ( .A(n6797), .B(n6798), .Z(o[6942]) );
  AND U10196 ( .A(p_input[26942]), .B(p_input[16942]), .Z(n6798) );
  AND U10197 ( .A(p_input[6942]), .B(p_input[36942]), .Z(n6797) );
  AND U10198 ( .A(n6799), .B(n6800), .Z(o[6941]) );
  AND U10199 ( .A(p_input[26941]), .B(p_input[16941]), .Z(n6800) );
  AND U10200 ( .A(p_input[6941]), .B(p_input[36941]), .Z(n6799) );
  AND U10201 ( .A(n6801), .B(n6802), .Z(o[6940]) );
  AND U10202 ( .A(p_input[26940]), .B(p_input[16940]), .Z(n6802) );
  AND U10203 ( .A(p_input[6940]), .B(p_input[36940]), .Z(n6801) );
  AND U10204 ( .A(n6803), .B(n6804), .Z(o[693]) );
  AND U10205 ( .A(p_input[20693]), .B(p_input[10693]), .Z(n6804) );
  AND U10206 ( .A(p_input[693]), .B(p_input[30693]), .Z(n6803) );
  AND U10207 ( .A(n6805), .B(n6806), .Z(o[6939]) );
  AND U10208 ( .A(p_input[26939]), .B(p_input[16939]), .Z(n6806) );
  AND U10209 ( .A(p_input[6939]), .B(p_input[36939]), .Z(n6805) );
  AND U10210 ( .A(n6807), .B(n6808), .Z(o[6938]) );
  AND U10211 ( .A(p_input[26938]), .B(p_input[16938]), .Z(n6808) );
  AND U10212 ( .A(p_input[6938]), .B(p_input[36938]), .Z(n6807) );
  AND U10213 ( .A(n6809), .B(n6810), .Z(o[6937]) );
  AND U10214 ( .A(p_input[26937]), .B(p_input[16937]), .Z(n6810) );
  AND U10215 ( .A(p_input[6937]), .B(p_input[36937]), .Z(n6809) );
  AND U10216 ( .A(n6811), .B(n6812), .Z(o[6936]) );
  AND U10217 ( .A(p_input[26936]), .B(p_input[16936]), .Z(n6812) );
  AND U10218 ( .A(p_input[6936]), .B(p_input[36936]), .Z(n6811) );
  AND U10219 ( .A(n6813), .B(n6814), .Z(o[6935]) );
  AND U10220 ( .A(p_input[26935]), .B(p_input[16935]), .Z(n6814) );
  AND U10221 ( .A(p_input[6935]), .B(p_input[36935]), .Z(n6813) );
  AND U10222 ( .A(n6815), .B(n6816), .Z(o[6934]) );
  AND U10223 ( .A(p_input[26934]), .B(p_input[16934]), .Z(n6816) );
  AND U10224 ( .A(p_input[6934]), .B(p_input[36934]), .Z(n6815) );
  AND U10225 ( .A(n6817), .B(n6818), .Z(o[6933]) );
  AND U10226 ( .A(p_input[26933]), .B(p_input[16933]), .Z(n6818) );
  AND U10227 ( .A(p_input[6933]), .B(p_input[36933]), .Z(n6817) );
  AND U10228 ( .A(n6819), .B(n6820), .Z(o[6932]) );
  AND U10229 ( .A(p_input[26932]), .B(p_input[16932]), .Z(n6820) );
  AND U10230 ( .A(p_input[6932]), .B(p_input[36932]), .Z(n6819) );
  AND U10231 ( .A(n6821), .B(n6822), .Z(o[6931]) );
  AND U10232 ( .A(p_input[26931]), .B(p_input[16931]), .Z(n6822) );
  AND U10233 ( .A(p_input[6931]), .B(p_input[36931]), .Z(n6821) );
  AND U10234 ( .A(n6823), .B(n6824), .Z(o[6930]) );
  AND U10235 ( .A(p_input[26930]), .B(p_input[16930]), .Z(n6824) );
  AND U10236 ( .A(p_input[6930]), .B(p_input[36930]), .Z(n6823) );
  AND U10237 ( .A(n6825), .B(n6826), .Z(o[692]) );
  AND U10238 ( .A(p_input[20692]), .B(p_input[10692]), .Z(n6826) );
  AND U10239 ( .A(p_input[692]), .B(p_input[30692]), .Z(n6825) );
  AND U10240 ( .A(n6827), .B(n6828), .Z(o[6929]) );
  AND U10241 ( .A(p_input[26929]), .B(p_input[16929]), .Z(n6828) );
  AND U10242 ( .A(p_input[6929]), .B(p_input[36929]), .Z(n6827) );
  AND U10243 ( .A(n6829), .B(n6830), .Z(o[6928]) );
  AND U10244 ( .A(p_input[26928]), .B(p_input[16928]), .Z(n6830) );
  AND U10245 ( .A(p_input[6928]), .B(p_input[36928]), .Z(n6829) );
  AND U10246 ( .A(n6831), .B(n6832), .Z(o[6927]) );
  AND U10247 ( .A(p_input[26927]), .B(p_input[16927]), .Z(n6832) );
  AND U10248 ( .A(p_input[6927]), .B(p_input[36927]), .Z(n6831) );
  AND U10249 ( .A(n6833), .B(n6834), .Z(o[6926]) );
  AND U10250 ( .A(p_input[26926]), .B(p_input[16926]), .Z(n6834) );
  AND U10251 ( .A(p_input[6926]), .B(p_input[36926]), .Z(n6833) );
  AND U10252 ( .A(n6835), .B(n6836), .Z(o[6925]) );
  AND U10253 ( .A(p_input[26925]), .B(p_input[16925]), .Z(n6836) );
  AND U10254 ( .A(p_input[6925]), .B(p_input[36925]), .Z(n6835) );
  AND U10255 ( .A(n6837), .B(n6838), .Z(o[6924]) );
  AND U10256 ( .A(p_input[26924]), .B(p_input[16924]), .Z(n6838) );
  AND U10257 ( .A(p_input[6924]), .B(p_input[36924]), .Z(n6837) );
  AND U10258 ( .A(n6839), .B(n6840), .Z(o[6923]) );
  AND U10259 ( .A(p_input[26923]), .B(p_input[16923]), .Z(n6840) );
  AND U10260 ( .A(p_input[6923]), .B(p_input[36923]), .Z(n6839) );
  AND U10261 ( .A(n6841), .B(n6842), .Z(o[6922]) );
  AND U10262 ( .A(p_input[26922]), .B(p_input[16922]), .Z(n6842) );
  AND U10263 ( .A(p_input[6922]), .B(p_input[36922]), .Z(n6841) );
  AND U10264 ( .A(n6843), .B(n6844), .Z(o[6921]) );
  AND U10265 ( .A(p_input[26921]), .B(p_input[16921]), .Z(n6844) );
  AND U10266 ( .A(p_input[6921]), .B(p_input[36921]), .Z(n6843) );
  AND U10267 ( .A(n6845), .B(n6846), .Z(o[6920]) );
  AND U10268 ( .A(p_input[26920]), .B(p_input[16920]), .Z(n6846) );
  AND U10269 ( .A(p_input[6920]), .B(p_input[36920]), .Z(n6845) );
  AND U10270 ( .A(n6847), .B(n6848), .Z(o[691]) );
  AND U10271 ( .A(p_input[20691]), .B(p_input[10691]), .Z(n6848) );
  AND U10272 ( .A(p_input[691]), .B(p_input[30691]), .Z(n6847) );
  AND U10273 ( .A(n6849), .B(n6850), .Z(o[6919]) );
  AND U10274 ( .A(p_input[26919]), .B(p_input[16919]), .Z(n6850) );
  AND U10275 ( .A(p_input[6919]), .B(p_input[36919]), .Z(n6849) );
  AND U10276 ( .A(n6851), .B(n6852), .Z(o[6918]) );
  AND U10277 ( .A(p_input[26918]), .B(p_input[16918]), .Z(n6852) );
  AND U10278 ( .A(p_input[6918]), .B(p_input[36918]), .Z(n6851) );
  AND U10279 ( .A(n6853), .B(n6854), .Z(o[6917]) );
  AND U10280 ( .A(p_input[26917]), .B(p_input[16917]), .Z(n6854) );
  AND U10281 ( .A(p_input[6917]), .B(p_input[36917]), .Z(n6853) );
  AND U10282 ( .A(n6855), .B(n6856), .Z(o[6916]) );
  AND U10283 ( .A(p_input[26916]), .B(p_input[16916]), .Z(n6856) );
  AND U10284 ( .A(p_input[6916]), .B(p_input[36916]), .Z(n6855) );
  AND U10285 ( .A(n6857), .B(n6858), .Z(o[6915]) );
  AND U10286 ( .A(p_input[26915]), .B(p_input[16915]), .Z(n6858) );
  AND U10287 ( .A(p_input[6915]), .B(p_input[36915]), .Z(n6857) );
  AND U10288 ( .A(n6859), .B(n6860), .Z(o[6914]) );
  AND U10289 ( .A(p_input[26914]), .B(p_input[16914]), .Z(n6860) );
  AND U10290 ( .A(p_input[6914]), .B(p_input[36914]), .Z(n6859) );
  AND U10291 ( .A(n6861), .B(n6862), .Z(o[6913]) );
  AND U10292 ( .A(p_input[26913]), .B(p_input[16913]), .Z(n6862) );
  AND U10293 ( .A(p_input[6913]), .B(p_input[36913]), .Z(n6861) );
  AND U10294 ( .A(n6863), .B(n6864), .Z(o[6912]) );
  AND U10295 ( .A(p_input[26912]), .B(p_input[16912]), .Z(n6864) );
  AND U10296 ( .A(p_input[6912]), .B(p_input[36912]), .Z(n6863) );
  AND U10297 ( .A(n6865), .B(n6866), .Z(o[6911]) );
  AND U10298 ( .A(p_input[26911]), .B(p_input[16911]), .Z(n6866) );
  AND U10299 ( .A(p_input[6911]), .B(p_input[36911]), .Z(n6865) );
  AND U10300 ( .A(n6867), .B(n6868), .Z(o[6910]) );
  AND U10301 ( .A(p_input[26910]), .B(p_input[16910]), .Z(n6868) );
  AND U10302 ( .A(p_input[6910]), .B(p_input[36910]), .Z(n6867) );
  AND U10303 ( .A(n6869), .B(n6870), .Z(o[690]) );
  AND U10304 ( .A(p_input[20690]), .B(p_input[10690]), .Z(n6870) );
  AND U10305 ( .A(p_input[690]), .B(p_input[30690]), .Z(n6869) );
  AND U10306 ( .A(n6871), .B(n6872), .Z(o[6909]) );
  AND U10307 ( .A(p_input[26909]), .B(p_input[16909]), .Z(n6872) );
  AND U10308 ( .A(p_input[6909]), .B(p_input[36909]), .Z(n6871) );
  AND U10309 ( .A(n6873), .B(n6874), .Z(o[6908]) );
  AND U10310 ( .A(p_input[26908]), .B(p_input[16908]), .Z(n6874) );
  AND U10311 ( .A(p_input[6908]), .B(p_input[36908]), .Z(n6873) );
  AND U10312 ( .A(n6875), .B(n6876), .Z(o[6907]) );
  AND U10313 ( .A(p_input[26907]), .B(p_input[16907]), .Z(n6876) );
  AND U10314 ( .A(p_input[6907]), .B(p_input[36907]), .Z(n6875) );
  AND U10315 ( .A(n6877), .B(n6878), .Z(o[6906]) );
  AND U10316 ( .A(p_input[26906]), .B(p_input[16906]), .Z(n6878) );
  AND U10317 ( .A(p_input[6906]), .B(p_input[36906]), .Z(n6877) );
  AND U10318 ( .A(n6879), .B(n6880), .Z(o[6905]) );
  AND U10319 ( .A(p_input[26905]), .B(p_input[16905]), .Z(n6880) );
  AND U10320 ( .A(p_input[6905]), .B(p_input[36905]), .Z(n6879) );
  AND U10321 ( .A(n6881), .B(n6882), .Z(o[6904]) );
  AND U10322 ( .A(p_input[26904]), .B(p_input[16904]), .Z(n6882) );
  AND U10323 ( .A(p_input[6904]), .B(p_input[36904]), .Z(n6881) );
  AND U10324 ( .A(n6883), .B(n6884), .Z(o[6903]) );
  AND U10325 ( .A(p_input[26903]), .B(p_input[16903]), .Z(n6884) );
  AND U10326 ( .A(p_input[6903]), .B(p_input[36903]), .Z(n6883) );
  AND U10327 ( .A(n6885), .B(n6886), .Z(o[6902]) );
  AND U10328 ( .A(p_input[26902]), .B(p_input[16902]), .Z(n6886) );
  AND U10329 ( .A(p_input[6902]), .B(p_input[36902]), .Z(n6885) );
  AND U10330 ( .A(n6887), .B(n6888), .Z(o[6901]) );
  AND U10331 ( .A(p_input[26901]), .B(p_input[16901]), .Z(n6888) );
  AND U10332 ( .A(p_input[6901]), .B(p_input[36901]), .Z(n6887) );
  AND U10333 ( .A(n6889), .B(n6890), .Z(o[6900]) );
  AND U10334 ( .A(p_input[26900]), .B(p_input[16900]), .Z(n6890) );
  AND U10335 ( .A(p_input[6900]), .B(p_input[36900]), .Z(n6889) );
  AND U10336 ( .A(n6891), .B(n6892), .Z(o[68]) );
  AND U10337 ( .A(p_input[20068]), .B(p_input[10068]), .Z(n6892) );
  AND U10338 ( .A(p_input[68]), .B(p_input[30068]), .Z(n6891) );
  AND U10339 ( .A(n6893), .B(n6894), .Z(o[689]) );
  AND U10340 ( .A(p_input[20689]), .B(p_input[10689]), .Z(n6894) );
  AND U10341 ( .A(p_input[689]), .B(p_input[30689]), .Z(n6893) );
  AND U10342 ( .A(n6895), .B(n6896), .Z(o[6899]) );
  AND U10343 ( .A(p_input[26899]), .B(p_input[16899]), .Z(n6896) );
  AND U10344 ( .A(p_input[6899]), .B(p_input[36899]), .Z(n6895) );
  AND U10345 ( .A(n6897), .B(n6898), .Z(o[6898]) );
  AND U10346 ( .A(p_input[26898]), .B(p_input[16898]), .Z(n6898) );
  AND U10347 ( .A(p_input[6898]), .B(p_input[36898]), .Z(n6897) );
  AND U10348 ( .A(n6899), .B(n6900), .Z(o[6897]) );
  AND U10349 ( .A(p_input[26897]), .B(p_input[16897]), .Z(n6900) );
  AND U10350 ( .A(p_input[6897]), .B(p_input[36897]), .Z(n6899) );
  AND U10351 ( .A(n6901), .B(n6902), .Z(o[6896]) );
  AND U10352 ( .A(p_input[26896]), .B(p_input[16896]), .Z(n6902) );
  AND U10353 ( .A(p_input[6896]), .B(p_input[36896]), .Z(n6901) );
  AND U10354 ( .A(n6903), .B(n6904), .Z(o[6895]) );
  AND U10355 ( .A(p_input[26895]), .B(p_input[16895]), .Z(n6904) );
  AND U10356 ( .A(p_input[6895]), .B(p_input[36895]), .Z(n6903) );
  AND U10357 ( .A(n6905), .B(n6906), .Z(o[6894]) );
  AND U10358 ( .A(p_input[26894]), .B(p_input[16894]), .Z(n6906) );
  AND U10359 ( .A(p_input[6894]), .B(p_input[36894]), .Z(n6905) );
  AND U10360 ( .A(n6907), .B(n6908), .Z(o[6893]) );
  AND U10361 ( .A(p_input[26893]), .B(p_input[16893]), .Z(n6908) );
  AND U10362 ( .A(p_input[6893]), .B(p_input[36893]), .Z(n6907) );
  AND U10363 ( .A(n6909), .B(n6910), .Z(o[6892]) );
  AND U10364 ( .A(p_input[26892]), .B(p_input[16892]), .Z(n6910) );
  AND U10365 ( .A(p_input[6892]), .B(p_input[36892]), .Z(n6909) );
  AND U10366 ( .A(n6911), .B(n6912), .Z(o[6891]) );
  AND U10367 ( .A(p_input[26891]), .B(p_input[16891]), .Z(n6912) );
  AND U10368 ( .A(p_input[6891]), .B(p_input[36891]), .Z(n6911) );
  AND U10369 ( .A(n6913), .B(n6914), .Z(o[6890]) );
  AND U10370 ( .A(p_input[26890]), .B(p_input[16890]), .Z(n6914) );
  AND U10371 ( .A(p_input[6890]), .B(p_input[36890]), .Z(n6913) );
  AND U10372 ( .A(n6915), .B(n6916), .Z(o[688]) );
  AND U10373 ( .A(p_input[20688]), .B(p_input[10688]), .Z(n6916) );
  AND U10374 ( .A(p_input[688]), .B(p_input[30688]), .Z(n6915) );
  AND U10375 ( .A(n6917), .B(n6918), .Z(o[6889]) );
  AND U10376 ( .A(p_input[26889]), .B(p_input[16889]), .Z(n6918) );
  AND U10377 ( .A(p_input[6889]), .B(p_input[36889]), .Z(n6917) );
  AND U10378 ( .A(n6919), .B(n6920), .Z(o[6888]) );
  AND U10379 ( .A(p_input[26888]), .B(p_input[16888]), .Z(n6920) );
  AND U10380 ( .A(p_input[6888]), .B(p_input[36888]), .Z(n6919) );
  AND U10381 ( .A(n6921), .B(n6922), .Z(o[6887]) );
  AND U10382 ( .A(p_input[26887]), .B(p_input[16887]), .Z(n6922) );
  AND U10383 ( .A(p_input[6887]), .B(p_input[36887]), .Z(n6921) );
  AND U10384 ( .A(n6923), .B(n6924), .Z(o[6886]) );
  AND U10385 ( .A(p_input[26886]), .B(p_input[16886]), .Z(n6924) );
  AND U10386 ( .A(p_input[6886]), .B(p_input[36886]), .Z(n6923) );
  AND U10387 ( .A(n6925), .B(n6926), .Z(o[6885]) );
  AND U10388 ( .A(p_input[26885]), .B(p_input[16885]), .Z(n6926) );
  AND U10389 ( .A(p_input[6885]), .B(p_input[36885]), .Z(n6925) );
  AND U10390 ( .A(n6927), .B(n6928), .Z(o[6884]) );
  AND U10391 ( .A(p_input[26884]), .B(p_input[16884]), .Z(n6928) );
  AND U10392 ( .A(p_input[6884]), .B(p_input[36884]), .Z(n6927) );
  AND U10393 ( .A(n6929), .B(n6930), .Z(o[6883]) );
  AND U10394 ( .A(p_input[26883]), .B(p_input[16883]), .Z(n6930) );
  AND U10395 ( .A(p_input[6883]), .B(p_input[36883]), .Z(n6929) );
  AND U10396 ( .A(n6931), .B(n6932), .Z(o[6882]) );
  AND U10397 ( .A(p_input[26882]), .B(p_input[16882]), .Z(n6932) );
  AND U10398 ( .A(p_input[6882]), .B(p_input[36882]), .Z(n6931) );
  AND U10399 ( .A(n6933), .B(n6934), .Z(o[6881]) );
  AND U10400 ( .A(p_input[26881]), .B(p_input[16881]), .Z(n6934) );
  AND U10401 ( .A(p_input[6881]), .B(p_input[36881]), .Z(n6933) );
  AND U10402 ( .A(n6935), .B(n6936), .Z(o[6880]) );
  AND U10403 ( .A(p_input[26880]), .B(p_input[16880]), .Z(n6936) );
  AND U10404 ( .A(p_input[6880]), .B(p_input[36880]), .Z(n6935) );
  AND U10405 ( .A(n6937), .B(n6938), .Z(o[687]) );
  AND U10406 ( .A(p_input[20687]), .B(p_input[10687]), .Z(n6938) );
  AND U10407 ( .A(p_input[687]), .B(p_input[30687]), .Z(n6937) );
  AND U10408 ( .A(n6939), .B(n6940), .Z(o[6879]) );
  AND U10409 ( .A(p_input[26879]), .B(p_input[16879]), .Z(n6940) );
  AND U10410 ( .A(p_input[6879]), .B(p_input[36879]), .Z(n6939) );
  AND U10411 ( .A(n6941), .B(n6942), .Z(o[6878]) );
  AND U10412 ( .A(p_input[26878]), .B(p_input[16878]), .Z(n6942) );
  AND U10413 ( .A(p_input[6878]), .B(p_input[36878]), .Z(n6941) );
  AND U10414 ( .A(n6943), .B(n6944), .Z(o[6877]) );
  AND U10415 ( .A(p_input[26877]), .B(p_input[16877]), .Z(n6944) );
  AND U10416 ( .A(p_input[6877]), .B(p_input[36877]), .Z(n6943) );
  AND U10417 ( .A(n6945), .B(n6946), .Z(o[6876]) );
  AND U10418 ( .A(p_input[26876]), .B(p_input[16876]), .Z(n6946) );
  AND U10419 ( .A(p_input[6876]), .B(p_input[36876]), .Z(n6945) );
  AND U10420 ( .A(n6947), .B(n6948), .Z(o[6875]) );
  AND U10421 ( .A(p_input[26875]), .B(p_input[16875]), .Z(n6948) );
  AND U10422 ( .A(p_input[6875]), .B(p_input[36875]), .Z(n6947) );
  AND U10423 ( .A(n6949), .B(n6950), .Z(o[6874]) );
  AND U10424 ( .A(p_input[26874]), .B(p_input[16874]), .Z(n6950) );
  AND U10425 ( .A(p_input[6874]), .B(p_input[36874]), .Z(n6949) );
  AND U10426 ( .A(n6951), .B(n6952), .Z(o[6873]) );
  AND U10427 ( .A(p_input[26873]), .B(p_input[16873]), .Z(n6952) );
  AND U10428 ( .A(p_input[6873]), .B(p_input[36873]), .Z(n6951) );
  AND U10429 ( .A(n6953), .B(n6954), .Z(o[6872]) );
  AND U10430 ( .A(p_input[26872]), .B(p_input[16872]), .Z(n6954) );
  AND U10431 ( .A(p_input[6872]), .B(p_input[36872]), .Z(n6953) );
  AND U10432 ( .A(n6955), .B(n6956), .Z(o[6871]) );
  AND U10433 ( .A(p_input[26871]), .B(p_input[16871]), .Z(n6956) );
  AND U10434 ( .A(p_input[6871]), .B(p_input[36871]), .Z(n6955) );
  AND U10435 ( .A(n6957), .B(n6958), .Z(o[6870]) );
  AND U10436 ( .A(p_input[26870]), .B(p_input[16870]), .Z(n6958) );
  AND U10437 ( .A(p_input[6870]), .B(p_input[36870]), .Z(n6957) );
  AND U10438 ( .A(n6959), .B(n6960), .Z(o[686]) );
  AND U10439 ( .A(p_input[20686]), .B(p_input[10686]), .Z(n6960) );
  AND U10440 ( .A(p_input[686]), .B(p_input[30686]), .Z(n6959) );
  AND U10441 ( .A(n6961), .B(n6962), .Z(o[6869]) );
  AND U10442 ( .A(p_input[26869]), .B(p_input[16869]), .Z(n6962) );
  AND U10443 ( .A(p_input[6869]), .B(p_input[36869]), .Z(n6961) );
  AND U10444 ( .A(n6963), .B(n6964), .Z(o[6868]) );
  AND U10445 ( .A(p_input[26868]), .B(p_input[16868]), .Z(n6964) );
  AND U10446 ( .A(p_input[6868]), .B(p_input[36868]), .Z(n6963) );
  AND U10447 ( .A(n6965), .B(n6966), .Z(o[6867]) );
  AND U10448 ( .A(p_input[26867]), .B(p_input[16867]), .Z(n6966) );
  AND U10449 ( .A(p_input[6867]), .B(p_input[36867]), .Z(n6965) );
  AND U10450 ( .A(n6967), .B(n6968), .Z(o[6866]) );
  AND U10451 ( .A(p_input[26866]), .B(p_input[16866]), .Z(n6968) );
  AND U10452 ( .A(p_input[6866]), .B(p_input[36866]), .Z(n6967) );
  AND U10453 ( .A(n6969), .B(n6970), .Z(o[6865]) );
  AND U10454 ( .A(p_input[26865]), .B(p_input[16865]), .Z(n6970) );
  AND U10455 ( .A(p_input[6865]), .B(p_input[36865]), .Z(n6969) );
  AND U10456 ( .A(n6971), .B(n6972), .Z(o[6864]) );
  AND U10457 ( .A(p_input[26864]), .B(p_input[16864]), .Z(n6972) );
  AND U10458 ( .A(p_input[6864]), .B(p_input[36864]), .Z(n6971) );
  AND U10459 ( .A(n6973), .B(n6974), .Z(o[6863]) );
  AND U10460 ( .A(p_input[26863]), .B(p_input[16863]), .Z(n6974) );
  AND U10461 ( .A(p_input[6863]), .B(p_input[36863]), .Z(n6973) );
  AND U10462 ( .A(n6975), .B(n6976), .Z(o[6862]) );
  AND U10463 ( .A(p_input[26862]), .B(p_input[16862]), .Z(n6976) );
  AND U10464 ( .A(p_input[6862]), .B(p_input[36862]), .Z(n6975) );
  AND U10465 ( .A(n6977), .B(n6978), .Z(o[6861]) );
  AND U10466 ( .A(p_input[26861]), .B(p_input[16861]), .Z(n6978) );
  AND U10467 ( .A(p_input[6861]), .B(p_input[36861]), .Z(n6977) );
  AND U10468 ( .A(n6979), .B(n6980), .Z(o[6860]) );
  AND U10469 ( .A(p_input[26860]), .B(p_input[16860]), .Z(n6980) );
  AND U10470 ( .A(p_input[6860]), .B(p_input[36860]), .Z(n6979) );
  AND U10471 ( .A(n6981), .B(n6982), .Z(o[685]) );
  AND U10472 ( .A(p_input[20685]), .B(p_input[10685]), .Z(n6982) );
  AND U10473 ( .A(p_input[685]), .B(p_input[30685]), .Z(n6981) );
  AND U10474 ( .A(n6983), .B(n6984), .Z(o[6859]) );
  AND U10475 ( .A(p_input[26859]), .B(p_input[16859]), .Z(n6984) );
  AND U10476 ( .A(p_input[6859]), .B(p_input[36859]), .Z(n6983) );
  AND U10477 ( .A(n6985), .B(n6986), .Z(o[6858]) );
  AND U10478 ( .A(p_input[26858]), .B(p_input[16858]), .Z(n6986) );
  AND U10479 ( .A(p_input[6858]), .B(p_input[36858]), .Z(n6985) );
  AND U10480 ( .A(n6987), .B(n6988), .Z(o[6857]) );
  AND U10481 ( .A(p_input[26857]), .B(p_input[16857]), .Z(n6988) );
  AND U10482 ( .A(p_input[6857]), .B(p_input[36857]), .Z(n6987) );
  AND U10483 ( .A(n6989), .B(n6990), .Z(o[6856]) );
  AND U10484 ( .A(p_input[26856]), .B(p_input[16856]), .Z(n6990) );
  AND U10485 ( .A(p_input[6856]), .B(p_input[36856]), .Z(n6989) );
  AND U10486 ( .A(n6991), .B(n6992), .Z(o[6855]) );
  AND U10487 ( .A(p_input[26855]), .B(p_input[16855]), .Z(n6992) );
  AND U10488 ( .A(p_input[6855]), .B(p_input[36855]), .Z(n6991) );
  AND U10489 ( .A(n6993), .B(n6994), .Z(o[6854]) );
  AND U10490 ( .A(p_input[26854]), .B(p_input[16854]), .Z(n6994) );
  AND U10491 ( .A(p_input[6854]), .B(p_input[36854]), .Z(n6993) );
  AND U10492 ( .A(n6995), .B(n6996), .Z(o[6853]) );
  AND U10493 ( .A(p_input[26853]), .B(p_input[16853]), .Z(n6996) );
  AND U10494 ( .A(p_input[6853]), .B(p_input[36853]), .Z(n6995) );
  AND U10495 ( .A(n6997), .B(n6998), .Z(o[6852]) );
  AND U10496 ( .A(p_input[26852]), .B(p_input[16852]), .Z(n6998) );
  AND U10497 ( .A(p_input[6852]), .B(p_input[36852]), .Z(n6997) );
  AND U10498 ( .A(n6999), .B(n7000), .Z(o[6851]) );
  AND U10499 ( .A(p_input[26851]), .B(p_input[16851]), .Z(n7000) );
  AND U10500 ( .A(p_input[6851]), .B(p_input[36851]), .Z(n6999) );
  AND U10501 ( .A(n7001), .B(n7002), .Z(o[6850]) );
  AND U10502 ( .A(p_input[26850]), .B(p_input[16850]), .Z(n7002) );
  AND U10503 ( .A(p_input[6850]), .B(p_input[36850]), .Z(n7001) );
  AND U10504 ( .A(n7003), .B(n7004), .Z(o[684]) );
  AND U10505 ( .A(p_input[20684]), .B(p_input[10684]), .Z(n7004) );
  AND U10506 ( .A(p_input[684]), .B(p_input[30684]), .Z(n7003) );
  AND U10507 ( .A(n7005), .B(n7006), .Z(o[6849]) );
  AND U10508 ( .A(p_input[26849]), .B(p_input[16849]), .Z(n7006) );
  AND U10509 ( .A(p_input[6849]), .B(p_input[36849]), .Z(n7005) );
  AND U10510 ( .A(n7007), .B(n7008), .Z(o[6848]) );
  AND U10511 ( .A(p_input[26848]), .B(p_input[16848]), .Z(n7008) );
  AND U10512 ( .A(p_input[6848]), .B(p_input[36848]), .Z(n7007) );
  AND U10513 ( .A(n7009), .B(n7010), .Z(o[6847]) );
  AND U10514 ( .A(p_input[26847]), .B(p_input[16847]), .Z(n7010) );
  AND U10515 ( .A(p_input[6847]), .B(p_input[36847]), .Z(n7009) );
  AND U10516 ( .A(n7011), .B(n7012), .Z(o[6846]) );
  AND U10517 ( .A(p_input[26846]), .B(p_input[16846]), .Z(n7012) );
  AND U10518 ( .A(p_input[6846]), .B(p_input[36846]), .Z(n7011) );
  AND U10519 ( .A(n7013), .B(n7014), .Z(o[6845]) );
  AND U10520 ( .A(p_input[26845]), .B(p_input[16845]), .Z(n7014) );
  AND U10521 ( .A(p_input[6845]), .B(p_input[36845]), .Z(n7013) );
  AND U10522 ( .A(n7015), .B(n7016), .Z(o[6844]) );
  AND U10523 ( .A(p_input[26844]), .B(p_input[16844]), .Z(n7016) );
  AND U10524 ( .A(p_input[6844]), .B(p_input[36844]), .Z(n7015) );
  AND U10525 ( .A(n7017), .B(n7018), .Z(o[6843]) );
  AND U10526 ( .A(p_input[26843]), .B(p_input[16843]), .Z(n7018) );
  AND U10527 ( .A(p_input[6843]), .B(p_input[36843]), .Z(n7017) );
  AND U10528 ( .A(n7019), .B(n7020), .Z(o[6842]) );
  AND U10529 ( .A(p_input[26842]), .B(p_input[16842]), .Z(n7020) );
  AND U10530 ( .A(p_input[6842]), .B(p_input[36842]), .Z(n7019) );
  AND U10531 ( .A(n7021), .B(n7022), .Z(o[6841]) );
  AND U10532 ( .A(p_input[26841]), .B(p_input[16841]), .Z(n7022) );
  AND U10533 ( .A(p_input[6841]), .B(p_input[36841]), .Z(n7021) );
  AND U10534 ( .A(n7023), .B(n7024), .Z(o[6840]) );
  AND U10535 ( .A(p_input[26840]), .B(p_input[16840]), .Z(n7024) );
  AND U10536 ( .A(p_input[6840]), .B(p_input[36840]), .Z(n7023) );
  AND U10537 ( .A(n7025), .B(n7026), .Z(o[683]) );
  AND U10538 ( .A(p_input[20683]), .B(p_input[10683]), .Z(n7026) );
  AND U10539 ( .A(p_input[683]), .B(p_input[30683]), .Z(n7025) );
  AND U10540 ( .A(n7027), .B(n7028), .Z(o[6839]) );
  AND U10541 ( .A(p_input[26839]), .B(p_input[16839]), .Z(n7028) );
  AND U10542 ( .A(p_input[6839]), .B(p_input[36839]), .Z(n7027) );
  AND U10543 ( .A(n7029), .B(n7030), .Z(o[6838]) );
  AND U10544 ( .A(p_input[26838]), .B(p_input[16838]), .Z(n7030) );
  AND U10545 ( .A(p_input[6838]), .B(p_input[36838]), .Z(n7029) );
  AND U10546 ( .A(n7031), .B(n7032), .Z(o[6837]) );
  AND U10547 ( .A(p_input[26837]), .B(p_input[16837]), .Z(n7032) );
  AND U10548 ( .A(p_input[6837]), .B(p_input[36837]), .Z(n7031) );
  AND U10549 ( .A(n7033), .B(n7034), .Z(o[6836]) );
  AND U10550 ( .A(p_input[26836]), .B(p_input[16836]), .Z(n7034) );
  AND U10551 ( .A(p_input[6836]), .B(p_input[36836]), .Z(n7033) );
  AND U10552 ( .A(n7035), .B(n7036), .Z(o[6835]) );
  AND U10553 ( .A(p_input[26835]), .B(p_input[16835]), .Z(n7036) );
  AND U10554 ( .A(p_input[6835]), .B(p_input[36835]), .Z(n7035) );
  AND U10555 ( .A(n7037), .B(n7038), .Z(o[6834]) );
  AND U10556 ( .A(p_input[26834]), .B(p_input[16834]), .Z(n7038) );
  AND U10557 ( .A(p_input[6834]), .B(p_input[36834]), .Z(n7037) );
  AND U10558 ( .A(n7039), .B(n7040), .Z(o[6833]) );
  AND U10559 ( .A(p_input[26833]), .B(p_input[16833]), .Z(n7040) );
  AND U10560 ( .A(p_input[6833]), .B(p_input[36833]), .Z(n7039) );
  AND U10561 ( .A(n7041), .B(n7042), .Z(o[6832]) );
  AND U10562 ( .A(p_input[26832]), .B(p_input[16832]), .Z(n7042) );
  AND U10563 ( .A(p_input[6832]), .B(p_input[36832]), .Z(n7041) );
  AND U10564 ( .A(n7043), .B(n7044), .Z(o[6831]) );
  AND U10565 ( .A(p_input[26831]), .B(p_input[16831]), .Z(n7044) );
  AND U10566 ( .A(p_input[6831]), .B(p_input[36831]), .Z(n7043) );
  AND U10567 ( .A(n7045), .B(n7046), .Z(o[6830]) );
  AND U10568 ( .A(p_input[26830]), .B(p_input[16830]), .Z(n7046) );
  AND U10569 ( .A(p_input[6830]), .B(p_input[36830]), .Z(n7045) );
  AND U10570 ( .A(n7047), .B(n7048), .Z(o[682]) );
  AND U10571 ( .A(p_input[20682]), .B(p_input[10682]), .Z(n7048) );
  AND U10572 ( .A(p_input[682]), .B(p_input[30682]), .Z(n7047) );
  AND U10573 ( .A(n7049), .B(n7050), .Z(o[6829]) );
  AND U10574 ( .A(p_input[26829]), .B(p_input[16829]), .Z(n7050) );
  AND U10575 ( .A(p_input[6829]), .B(p_input[36829]), .Z(n7049) );
  AND U10576 ( .A(n7051), .B(n7052), .Z(o[6828]) );
  AND U10577 ( .A(p_input[26828]), .B(p_input[16828]), .Z(n7052) );
  AND U10578 ( .A(p_input[6828]), .B(p_input[36828]), .Z(n7051) );
  AND U10579 ( .A(n7053), .B(n7054), .Z(o[6827]) );
  AND U10580 ( .A(p_input[26827]), .B(p_input[16827]), .Z(n7054) );
  AND U10581 ( .A(p_input[6827]), .B(p_input[36827]), .Z(n7053) );
  AND U10582 ( .A(n7055), .B(n7056), .Z(o[6826]) );
  AND U10583 ( .A(p_input[26826]), .B(p_input[16826]), .Z(n7056) );
  AND U10584 ( .A(p_input[6826]), .B(p_input[36826]), .Z(n7055) );
  AND U10585 ( .A(n7057), .B(n7058), .Z(o[6825]) );
  AND U10586 ( .A(p_input[26825]), .B(p_input[16825]), .Z(n7058) );
  AND U10587 ( .A(p_input[6825]), .B(p_input[36825]), .Z(n7057) );
  AND U10588 ( .A(n7059), .B(n7060), .Z(o[6824]) );
  AND U10589 ( .A(p_input[26824]), .B(p_input[16824]), .Z(n7060) );
  AND U10590 ( .A(p_input[6824]), .B(p_input[36824]), .Z(n7059) );
  AND U10591 ( .A(n7061), .B(n7062), .Z(o[6823]) );
  AND U10592 ( .A(p_input[26823]), .B(p_input[16823]), .Z(n7062) );
  AND U10593 ( .A(p_input[6823]), .B(p_input[36823]), .Z(n7061) );
  AND U10594 ( .A(n7063), .B(n7064), .Z(o[6822]) );
  AND U10595 ( .A(p_input[26822]), .B(p_input[16822]), .Z(n7064) );
  AND U10596 ( .A(p_input[6822]), .B(p_input[36822]), .Z(n7063) );
  AND U10597 ( .A(n7065), .B(n7066), .Z(o[6821]) );
  AND U10598 ( .A(p_input[26821]), .B(p_input[16821]), .Z(n7066) );
  AND U10599 ( .A(p_input[6821]), .B(p_input[36821]), .Z(n7065) );
  AND U10600 ( .A(n7067), .B(n7068), .Z(o[6820]) );
  AND U10601 ( .A(p_input[26820]), .B(p_input[16820]), .Z(n7068) );
  AND U10602 ( .A(p_input[6820]), .B(p_input[36820]), .Z(n7067) );
  AND U10603 ( .A(n7069), .B(n7070), .Z(o[681]) );
  AND U10604 ( .A(p_input[20681]), .B(p_input[10681]), .Z(n7070) );
  AND U10605 ( .A(p_input[681]), .B(p_input[30681]), .Z(n7069) );
  AND U10606 ( .A(n7071), .B(n7072), .Z(o[6819]) );
  AND U10607 ( .A(p_input[26819]), .B(p_input[16819]), .Z(n7072) );
  AND U10608 ( .A(p_input[6819]), .B(p_input[36819]), .Z(n7071) );
  AND U10609 ( .A(n7073), .B(n7074), .Z(o[6818]) );
  AND U10610 ( .A(p_input[26818]), .B(p_input[16818]), .Z(n7074) );
  AND U10611 ( .A(p_input[6818]), .B(p_input[36818]), .Z(n7073) );
  AND U10612 ( .A(n7075), .B(n7076), .Z(o[6817]) );
  AND U10613 ( .A(p_input[26817]), .B(p_input[16817]), .Z(n7076) );
  AND U10614 ( .A(p_input[6817]), .B(p_input[36817]), .Z(n7075) );
  AND U10615 ( .A(n7077), .B(n7078), .Z(o[6816]) );
  AND U10616 ( .A(p_input[26816]), .B(p_input[16816]), .Z(n7078) );
  AND U10617 ( .A(p_input[6816]), .B(p_input[36816]), .Z(n7077) );
  AND U10618 ( .A(n7079), .B(n7080), .Z(o[6815]) );
  AND U10619 ( .A(p_input[26815]), .B(p_input[16815]), .Z(n7080) );
  AND U10620 ( .A(p_input[6815]), .B(p_input[36815]), .Z(n7079) );
  AND U10621 ( .A(n7081), .B(n7082), .Z(o[6814]) );
  AND U10622 ( .A(p_input[26814]), .B(p_input[16814]), .Z(n7082) );
  AND U10623 ( .A(p_input[6814]), .B(p_input[36814]), .Z(n7081) );
  AND U10624 ( .A(n7083), .B(n7084), .Z(o[6813]) );
  AND U10625 ( .A(p_input[26813]), .B(p_input[16813]), .Z(n7084) );
  AND U10626 ( .A(p_input[6813]), .B(p_input[36813]), .Z(n7083) );
  AND U10627 ( .A(n7085), .B(n7086), .Z(o[6812]) );
  AND U10628 ( .A(p_input[26812]), .B(p_input[16812]), .Z(n7086) );
  AND U10629 ( .A(p_input[6812]), .B(p_input[36812]), .Z(n7085) );
  AND U10630 ( .A(n7087), .B(n7088), .Z(o[6811]) );
  AND U10631 ( .A(p_input[26811]), .B(p_input[16811]), .Z(n7088) );
  AND U10632 ( .A(p_input[6811]), .B(p_input[36811]), .Z(n7087) );
  AND U10633 ( .A(n7089), .B(n7090), .Z(o[6810]) );
  AND U10634 ( .A(p_input[26810]), .B(p_input[16810]), .Z(n7090) );
  AND U10635 ( .A(p_input[6810]), .B(p_input[36810]), .Z(n7089) );
  AND U10636 ( .A(n7091), .B(n7092), .Z(o[680]) );
  AND U10637 ( .A(p_input[20680]), .B(p_input[10680]), .Z(n7092) );
  AND U10638 ( .A(p_input[680]), .B(p_input[30680]), .Z(n7091) );
  AND U10639 ( .A(n7093), .B(n7094), .Z(o[6809]) );
  AND U10640 ( .A(p_input[26809]), .B(p_input[16809]), .Z(n7094) );
  AND U10641 ( .A(p_input[6809]), .B(p_input[36809]), .Z(n7093) );
  AND U10642 ( .A(n7095), .B(n7096), .Z(o[6808]) );
  AND U10643 ( .A(p_input[26808]), .B(p_input[16808]), .Z(n7096) );
  AND U10644 ( .A(p_input[6808]), .B(p_input[36808]), .Z(n7095) );
  AND U10645 ( .A(n7097), .B(n7098), .Z(o[6807]) );
  AND U10646 ( .A(p_input[26807]), .B(p_input[16807]), .Z(n7098) );
  AND U10647 ( .A(p_input[6807]), .B(p_input[36807]), .Z(n7097) );
  AND U10648 ( .A(n7099), .B(n7100), .Z(o[6806]) );
  AND U10649 ( .A(p_input[26806]), .B(p_input[16806]), .Z(n7100) );
  AND U10650 ( .A(p_input[6806]), .B(p_input[36806]), .Z(n7099) );
  AND U10651 ( .A(n7101), .B(n7102), .Z(o[6805]) );
  AND U10652 ( .A(p_input[26805]), .B(p_input[16805]), .Z(n7102) );
  AND U10653 ( .A(p_input[6805]), .B(p_input[36805]), .Z(n7101) );
  AND U10654 ( .A(n7103), .B(n7104), .Z(o[6804]) );
  AND U10655 ( .A(p_input[26804]), .B(p_input[16804]), .Z(n7104) );
  AND U10656 ( .A(p_input[6804]), .B(p_input[36804]), .Z(n7103) );
  AND U10657 ( .A(n7105), .B(n7106), .Z(o[6803]) );
  AND U10658 ( .A(p_input[26803]), .B(p_input[16803]), .Z(n7106) );
  AND U10659 ( .A(p_input[6803]), .B(p_input[36803]), .Z(n7105) );
  AND U10660 ( .A(n7107), .B(n7108), .Z(o[6802]) );
  AND U10661 ( .A(p_input[26802]), .B(p_input[16802]), .Z(n7108) );
  AND U10662 ( .A(p_input[6802]), .B(p_input[36802]), .Z(n7107) );
  AND U10663 ( .A(n7109), .B(n7110), .Z(o[6801]) );
  AND U10664 ( .A(p_input[26801]), .B(p_input[16801]), .Z(n7110) );
  AND U10665 ( .A(p_input[6801]), .B(p_input[36801]), .Z(n7109) );
  AND U10666 ( .A(n7111), .B(n7112), .Z(o[6800]) );
  AND U10667 ( .A(p_input[26800]), .B(p_input[16800]), .Z(n7112) );
  AND U10668 ( .A(p_input[6800]), .B(p_input[36800]), .Z(n7111) );
  AND U10669 ( .A(n7113), .B(n7114), .Z(o[67]) );
  AND U10670 ( .A(p_input[20067]), .B(p_input[10067]), .Z(n7114) );
  AND U10671 ( .A(p_input[67]), .B(p_input[30067]), .Z(n7113) );
  AND U10672 ( .A(n7115), .B(n7116), .Z(o[679]) );
  AND U10673 ( .A(p_input[20679]), .B(p_input[10679]), .Z(n7116) );
  AND U10674 ( .A(p_input[679]), .B(p_input[30679]), .Z(n7115) );
  AND U10675 ( .A(n7117), .B(n7118), .Z(o[6799]) );
  AND U10676 ( .A(p_input[26799]), .B(p_input[16799]), .Z(n7118) );
  AND U10677 ( .A(p_input[6799]), .B(p_input[36799]), .Z(n7117) );
  AND U10678 ( .A(n7119), .B(n7120), .Z(o[6798]) );
  AND U10679 ( .A(p_input[26798]), .B(p_input[16798]), .Z(n7120) );
  AND U10680 ( .A(p_input[6798]), .B(p_input[36798]), .Z(n7119) );
  AND U10681 ( .A(n7121), .B(n7122), .Z(o[6797]) );
  AND U10682 ( .A(p_input[26797]), .B(p_input[16797]), .Z(n7122) );
  AND U10683 ( .A(p_input[6797]), .B(p_input[36797]), .Z(n7121) );
  AND U10684 ( .A(n7123), .B(n7124), .Z(o[6796]) );
  AND U10685 ( .A(p_input[26796]), .B(p_input[16796]), .Z(n7124) );
  AND U10686 ( .A(p_input[6796]), .B(p_input[36796]), .Z(n7123) );
  AND U10687 ( .A(n7125), .B(n7126), .Z(o[6795]) );
  AND U10688 ( .A(p_input[26795]), .B(p_input[16795]), .Z(n7126) );
  AND U10689 ( .A(p_input[6795]), .B(p_input[36795]), .Z(n7125) );
  AND U10690 ( .A(n7127), .B(n7128), .Z(o[6794]) );
  AND U10691 ( .A(p_input[26794]), .B(p_input[16794]), .Z(n7128) );
  AND U10692 ( .A(p_input[6794]), .B(p_input[36794]), .Z(n7127) );
  AND U10693 ( .A(n7129), .B(n7130), .Z(o[6793]) );
  AND U10694 ( .A(p_input[26793]), .B(p_input[16793]), .Z(n7130) );
  AND U10695 ( .A(p_input[6793]), .B(p_input[36793]), .Z(n7129) );
  AND U10696 ( .A(n7131), .B(n7132), .Z(o[6792]) );
  AND U10697 ( .A(p_input[26792]), .B(p_input[16792]), .Z(n7132) );
  AND U10698 ( .A(p_input[6792]), .B(p_input[36792]), .Z(n7131) );
  AND U10699 ( .A(n7133), .B(n7134), .Z(o[6791]) );
  AND U10700 ( .A(p_input[26791]), .B(p_input[16791]), .Z(n7134) );
  AND U10701 ( .A(p_input[6791]), .B(p_input[36791]), .Z(n7133) );
  AND U10702 ( .A(n7135), .B(n7136), .Z(o[6790]) );
  AND U10703 ( .A(p_input[26790]), .B(p_input[16790]), .Z(n7136) );
  AND U10704 ( .A(p_input[6790]), .B(p_input[36790]), .Z(n7135) );
  AND U10705 ( .A(n7137), .B(n7138), .Z(o[678]) );
  AND U10706 ( .A(p_input[20678]), .B(p_input[10678]), .Z(n7138) );
  AND U10707 ( .A(p_input[678]), .B(p_input[30678]), .Z(n7137) );
  AND U10708 ( .A(n7139), .B(n7140), .Z(o[6789]) );
  AND U10709 ( .A(p_input[26789]), .B(p_input[16789]), .Z(n7140) );
  AND U10710 ( .A(p_input[6789]), .B(p_input[36789]), .Z(n7139) );
  AND U10711 ( .A(n7141), .B(n7142), .Z(o[6788]) );
  AND U10712 ( .A(p_input[26788]), .B(p_input[16788]), .Z(n7142) );
  AND U10713 ( .A(p_input[6788]), .B(p_input[36788]), .Z(n7141) );
  AND U10714 ( .A(n7143), .B(n7144), .Z(o[6787]) );
  AND U10715 ( .A(p_input[26787]), .B(p_input[16787]), .Z(n7144) );
  AND U10716 ( .A(p_input[6787]), .B(p_input[36787]), .Z(n7143) );
  AND U10717 ( .A(n7145), .B(n7146), .Z(o[6786]) );
  AND U10718 ( .A(p_input[26786]), .B(p_input[16786]), .Z(n7146) );
  AND U10719 ( .A(p_input[6786]), .B(p_input[36786]), .Z(n7145) );
  AND U10720 ( .A(n7147), .B(n7148), .Z(o[6785]) );
  AND U10721 ( .A(p_input[26785]), .B(p_input[16785]), .Z(n7148) );
  AND U10722 ( .A(p_input[6785]), .B(p_input[36785]), .Z(n7147) );
  AND U10723 ( .A(n7149), .B(n7150), .Z(o[6784]) );
  AND U10724 ( .A(p_input[26784]), .B(p_input[16784]), .Z(n7150) );
  AND U10725 ( .A(p_input[6784]), .B(p_input[36784]), .Z(n7149) );
  AND U10726 ( .A(n7151), .B(n7152), .Z(o[6783]) );
  AND U10727 ( .A(p_input[26783]), .B(p_input[16783]), .Z(n7152) );
  AND U10728 ( .A(p_input[6783]), .B(p_input[36783]), .Z(n7151) );
  AND U10729 ( .A(n7153), .B(n7154), .Z(o[6782]) );
  AND U10730 ( .A(p_input[26782]), .B(p_input[16782]), .Z(n7154) );
  AND U10731 ( .A(p_input[6782]), .B(p_input[36782]), .Z(n7153) );
  AND U10732 ( .A(n7155), .B(n7156), .Z(o[6781]) );
  AND U10733 ( .A(p_input[26781]), .B(p_input[16781]), .Z(n7156) );
  AND U10734 ( .A(p_input[6781]), .B(p_input[36781]), .Z(n7155) );
  AND U10735 ( .A(n7157), .B(n7158), .Z(o[6780]) );
  AND U10736 ( .A(p_input[26780]), .B(p_input[16780]), .Z(n7158) );
  AND U10737 ( .A(p_input[6780]), .B(p_input[36780]), .Z(n7157) );
  AND U10738 ( .A(n7159), .B(n7160), .Z(o[677]) );
  AND U10739 ( .A(p_input[20677]), .B(p_input[10677]), .Z(n7160) );
  AND U10740 ( .A(p_input[677]), .B(p_input[30677]), .Z(n7159) );
  AND U10741 ( .A(n7161), .B(n7162), .Z(o[6779]) );
  AND U10742 ( .A(p_input[26779]), .B(p_input[16779]), .Z(n7162) );
  AND U10743 ( .A(p_input[6779]), .B(p_input[36779]), .Z(n7161) );
  AND U10744 ( .A(n7163), .B(n7164), .Z(o[6778]) );
  AND U10745 ( .A(p_input[26778]), .B(p_input[16778]), .Z(n7164) );
  AND U10746 ( .A(p_input[6778]), .B(p_input[36778]), .Z(n7163) );
  AND U10747 ( .A(n7165), .B(n7166), .Z(o[6777]) );
  AND U10748 ( .A(p_input[26777]), .B(p_input[16777]), .Z(n7166) );
  AND U10749 ( .A(p_input[6777]), .B(p_input[36777]), .Z(n7165) );
  AND U10750 ( .A(n7167), .B(n7168), .Z(o[6776]) );
  AND U10751 ( .A(p_input[26776]), .B(p_input[16776]), .Z(n7168) );
  AND U10752 ( .A(p_input[6776]), .B(p_input[36776]), .Z(n7167) );
  AND U10753 ( .A(n7169), .B(n7170), .Z(o[6775]) );
  AND U10754 ( .A(p_input[26775]), .B(p_input[16775]), .Z(n7170) );
  AND U10755 ( .A(p_input[6775]), .B(p_input[36775]), .Z(n7169) );
  AND U10756 ( .A(n7171), .B(n7172), .Z(o[6774]) );
  AND U10757 ( .A(p_input[26774]), .B(p_input[16774]), .Z(n7172) );
  AND U10758 ( .A(p_input[6774]), .B(p_input[36774]), .Z(n7171) );
  AND U10759 ( .A(n7173), .B(n7174), .Z(o[6773]) );
  AND U10760 ( .A(p_input[26773]), .B(p_input[16773]), .Z(n7174) );
  AND U10761 ( .A(p_input[6773]), .B(p_input[36773]), .Z(n7173) );
  AND U10762 ( .A(n7175), .B(n7176), .Z(o[6772]) );
  AND U10763 ( .A(p_input[26772]), .B(p_input[16772]), .Z(n7176) );
  AND U10764 ( .A(p_input[6772]), .B(p_input[36772]), .Z(n7175) );
  AND U10765 ( .A(n7177), .B(n7178), .Z(o[6771]) );
  AND U10766 ( .A(p_input[26771]), .B(p_input[16771]), .Z(n7178) );
  AND U10767 ( .A(p_input[6771]), .B(p_input[36771]), .Z(n7177) );
  AND U10768 ( .A(n7179), .B(n7180), .Z(o[6770]) );
  AND U10769 ( .A(p_input[26770]), .B(p_input[16770]), .Z(n7180) );
  AND U10770 ( .A(p_input[6770]), .B(p_input[36770]), .Z(n7179) );
  AND U10771 ( .A(n7181), .B(n7182), .Z(o[676]) );
  AND U10772 ( .A(p_input[20676]), .B(p_input[10676]), .Z(n7182) );
  AND U10773 ( .A(p_input[676]), .B(p_input[30676]), .Z(n7181) );
  AND U10774 ( .A(n7183), .B(n7184), .Z(o[6769]) );
  AND U10775 ( .A(p_input[26769]), .B(p_input[16769]), .Z(n7184) );
  AND U10776 ( .A(p_input[6769]), .B(p_input[36769]), .Z(n7183) );
  AND U10777 ( .A(n7185), .B(n7186), .Z(o[6768]) );
  AND U10778 ( .A(p_input[26768]), .B(p_input[16768]), .Z(n7186) );
  AND U10779 ( .A(p_input[6768]), .B(p_input[36768]), .Z(n7185) );
  AND U10780 ( .A(n7187), .B(n7188), .Z(o[6767]) );
  AND U10781 ( .A(p_input[26767]), .B(p_input[16767]), .Z(n7188) );
  AND U10782 ( .A(p_input[6767]), .B(p_input[36767]), .Z(n7187) );
  AND U10783 ( .A(n7189), .B(n7190), .Z(o[6766]) );
  AND U10784 ( .A(p_input[26766]), .B(p_input[16766]), .Z(n7190) );
  AND U10785 ( .A(p_input[6766]), .B(p_input[36766]), .Z(n7189) );
  AND U10786 ( .A(n7191), .B(n7192), .Z(o[6765]) );
  AND U10787 ( .A(p_input[26765]), .B(p_input[16765]), .Z(n7192) );
  AND U10788 ( .A(p_input[6765]), .B(p_input[36765]), .Z(n7191) );
  AND U10789 ( .A(n7193), .B(n7194), .Z(o[6764]) );
  AND U10790 ( .A(p_input[26764]), .B(p_input[16764]), .Z(n7194) );
  AND U10791 ( .A(p_input[6764]), .B(p_input[36764]), .Z(n7193) );
  AND U10792 ( .A(n7195), .B(n7196), .Z(o[6763]) );
  AND U10793 ( .A(p_input[26763]), .B(p_input[16763]), .Z(n7196) );
  AND U10794 ( .A(p_input[6763]), .B(p_input[36763]), .Z(n7195) );
  AND U10795 ( .A(n7197), .B(n7198), .Z(o[6762]) );
  AND U10796 ( .A(p_input[26762]), .B(p_input[16762]), .Z(n7198) );
  AND U10797 ( .A(p_input[6762]), .B(p_input[36762]), .Z(n7197) );
  AND U10798 ( .A(n7199), .B(n7200), .Z(o[6761]) );
  AND U10799 ( .A(p_input[26761]), .B(p_input[16761]), .Z(n7200) );
  AND U10800 ( .A(p_input[6761]), .B(p_input[36761]), .Z(n7199) );
  AND U10801 ( .A(n7201), .B(n7202), .Z(o[6760]) );
  AND U10802 ( .A(p_input[26760]), .B(p_input[16760]), .Z(n7202) );
  AND U10803 ( .A(p_input[6760]), .B(p_input[36760]), .Z(n7201) );
  AND U10804 ( .A(n7203), .B(n7204), .Z(o[675]) );
  AND U10805 ( .A(p_input[20675]), .B(p_input[10675]), .Z(n7204) );
  AND U10806 ( .A(p_input[675]), .B(p_input[30675]), .Z(n7203) );
  AND U10807 ( .A(n7205), .B(n7206), .Z(o[6759]) );
  AND U10808 ( .A(p_input[26759]), .B(p_input[16759]), .Z(n7206) );
  AND U10809 ( .A(p_input[6759]), .B(p_input[36759]), .Z(n7205) );
  AND U10810 ( .A(n7207), .B(n7208), .Z(o[6758]) );
  AND U10811 ( .A(p_input[26758]), .B(p_input[16758]), .Z(n7208) );
  AND U10812 ( .A(p_input[6758]), .B(p_input[36758]), .Z(n7207) );
  AND U10813 ( .A(n7209), .B(n7210), .Z(o[6757]) );
  AND U10814 ( .A(p_input[26757]), .B(p_input[16757]), .Z(n7210) );
  AND U10815 ( .A(p_input[6757]), .B(p_input[36757]), .Z(n7209) );
  AND U10816 ( .A(n7211), .B(n7212), .Z(o[6756]) );
  AND U10817 ( .A(p_input[26756]), .B(p_input[16756]), .Z(n7212) );
  AND U10818 ( .A(p_input[6756]), .B(p_input[36756]), .Z(n7211) );
  AND U10819 ( .A(n7213), .B(n7214), .Z(o[6755]) );
  AND U10820 ( .A(p_input[26755]), .B(p_input[16755]), .Z(n7214) );
  AND U10821 ( .A(p_input[6755]), .B(p_input[36755]), .Z(n7213) );
  AND U10822 ( .A(n7215), .B(n7216), .Z(o[6754]) );
  AND U10823 ( .A(p_input[26754]), .B(p_input[16754]), .Z(n7216) );
  AND U10824 ( .A(p_input[6754]), .B(p_input[36754]), .Z(n7215) );
  AND U10825 ( .A(n7217), .B(n7218), .Z(o[6753]) );
  AND U10826 ( .A(p_input[26753]), .B(p_input[16753]), .Z(n7218) );
  AND U10827 ( .A(p_input[6753]), .B(p_input[36753]), .Z(n7217) );
  AND U10828 ( .A(n7219), .B(n7220), .Z(o[6752]) );
  AND U10829 ( .A(p_input[26752]), .B(p_input[16752]), .Z(n7220) );
  AND U10830 ( .A(p_input[6752]), .B(p_input[36752]), .Z(n7219) );
  AND U10831 ( .A(n7221), .B(n7222), .Z(o[6751]) );
  AND U10832 ( .A(p_input[26751]), .B(p_input[16751]), .Z(n7222) );
  AND U10833 ( .A(p_input[6751]), .B(p_input[36751]), .Z(n7221) );
  AND U10834 ( .A(n7223), .B(n7224), .Z(o[6750]) );
  AND U10835 ( .A(p_input[26750]), .B(p_input[16750]), .Z(n7224) );
  AND U10836 ( .A(p_input[6750]), .B(p_input[36750]), .Z(n7223) );
  AND U10837 ( .A(n7225), .B(n7226), .Z(o[674]) );
  AND U10838 ( .A(p_input[20674]), .B(p_input[10674]), .Z(n7226) );
  AND U10839 ( .A(p_input[674]), .B(p_input[30674]), .Z(n7225) );
  AND U10840 ( .A(n7227), .B(n7228), .Z(o[6749]) );
  AND U10841 ( .A(p_input[26749]), .B(p_input[16749]), .Z(n7228) );
  AND U10842 ( .A(p_input[6749]), .B(p_input[36749]), .Z(n7227) );
  AND U10843 ( .A(n7229), .B(n7230), .Z(o[6748]) );
  AND U10844 ( .A(p_input[26748]), .B(p_input[16748]), .Z(n7230) );
  AND U10845 ( .A(p_input[6748]), .B(p_input[36748]), .Z(n7229) );
  AND U10846 ( .A(n7231), .B(n7232), .Z(o[6747]) );
  AND U10847 ( .A(p_input[26747]), .B(p_input[16747]), .Z(n7232) );
  AND U10848 ( .A(p_input[6747]), .B(p_input[36747]), .Z(n7231) );
  AND U10849 ( .A(n7233), .B(n7234), .Z(o[6746]) );
  AND U10850 ( .A(p_input[26746]), .B(p_input[16746]), .Z(n7234) );
  AND U10851 ( .A(p_input[6746]), .B(p_input[36746]), .Z(n7233) );
  AND U10852 ( .A(n7235), .B(n7236), .Z(o[6745]) );
  AND U10853 ( .A(p_input[26745]), .B(p_input[16745]), .Z(n7236) );
  AND U10854 ( .A(p_input[6745]), .B(p_input[36745]), .Z(n7235) );
  AND U10855 ( .A(n7237), .B(n7238), .Z(o[6744]) );
  AND U10856 ( .A(p_input[26744]), .B(p_input[16744]), .Z(n7238) );
  AND U10857 ( .A(p_input[6744]), .B(p_input[36744]), .Z(n7237) );
  AND U10858 ( .A(n7239), .B(n7240), .Z(o[6743]) );
  AND U10859 ( .A(p_input[26743]), .B(p_input[16743]), .Z(n7240) );
  AND U10860 ( .A(p_input[6743]), .B(p_input[36743]), .Z(n7239) );
  AND U10861 ( .A(n7241), .B(n7242), .Z(o[6742]) );
  AND U10862 ( .A(p_input[26742]), .B(p_input[16742]), .Z(n7242) );
  AND U10863 ( .A(p_input[6742]), .B(p_input[36742]), .Z(n7241) );
  AND U10864 ( .A(n7243), .B(n7244), .Z(o[6741]) );
  AND U10865 ( .A(p_input[26741]), .B(p_input[16741]), .Z(n7244) );
  AND U10866 ( .A(p_input[6741]), .B(p_input[36741]), .Z(n7243) );
  AND U10867 ( .A(n7245), .B(n7246), .Z(o[6740]) );
  AND U10868 ( .A(p_input[26740]), .B(p_input[16740]), .Z(n7246) );
  AND U10869 ( .A(p_input[6740]), .B(p_input[36740]), .Z(n7245) );
  AND U10870 ( .A(n7247), .B(n7248), .Z(o[673]) );
  AND U10871 ( .A(p_input[20673]), .B(p_input[10673]), .Z(n7248) );
  AND U10872 ( .A(p_input[673]), .B(p_input[30673]), .Z(n7247) );
  AND U10873 ( .A(n7249), .B(n7250), .Z(o[6739]) );
  AND U10874 ( .A(p_input[26739]), .B(p_input[16739]), .Z(n7250) );
  AND U10875 ( .A(p_input[6739]), .B(p_input[36739]), .Z(n7249) );
  AND U10876 ( .A(n7251), .B(n7252), .Z(o[6738]) );
  AND U10877 ( .A(p_input[26738]), .B(p_input[16738]), .Z(n7252) );
  AND U10878 ( .A(p_input[6738]), .B(p_input[36738]), .Z(n7251) );
  AND U10879 ( .A(n7253), .B(n7254), .Z(o[6737]) );
  AND U10880 ( .A(p_input[26737]), .B(p_input[16737]), .Z(n7254) );
  AND U10881 ( .A(p_input[6737]), .B(p_input[36737]), .Z(n7253) );
  AND U10882 ( .A(n7255), .B(n7256), .Z(o[6736]) );
  AND U10883 ( .A(p_input[26736]), .B(p_input[16736]), .Z(n7256) );
  AND U10884 ( .A(p_input[6736]), .B(p_input[36736]), .Z(n7255) );
  AND U10885 ( .A(n7257), .B(n7258), .Z(o[6735]) );
  AND U10886 ( .A(p_input[26735]), .B(p_input[16735]), .Z(n7258) );
  AND U10887 ( .A(p_input[6735]), .B(p_input[36735]), .Z(n7257) );
  AND U10888 ( .A(n7259), .B(n7260), .Z(o[6734]) );
  AND U10889 ( .A(p_input[26734]), .B(p_input[16734]), .Z(n7260) );
  AND U10890 ( .A(p_input[6734]), .B(p_input[36734]), .Z(n7259) );
  AND U10891 ( .A(n7261), .B(n7262), .Z(o[6733]) );
  AND U10892 ( .A(p_input[26733]), .B(p_input[16733]), .Z(n7262) );
  AND U10893 ( .A(p_input[6733]), .B(p_input[36733]), .Z(n7261) );
  AND U10894 ( .A(n7263), .B(n7264), .Z(o[6732]) );
  AND U10895 ( .A(p_input[26732]), .B(p_input[16732]), .Z(n7264) );
  AND U10896 ( .A(p_input[6732]), .B(p_input[36732]), .Z(n7263) );
  AND U10897 ( .A(n7265), .B(n7266), .Z(o[6731]) );
  AND U10898 ( .A(p_input[26731]), .B(p_input[16731]), .Z(n7266) );
  AND U10899 ( .A(p_input[6731]), .B(p_input[36731]), .Z(n7265) );
  AND U10900 ( .A(n7267), .B(n7268), .Z(o[6730]) );
  AND U10901 ( .A(p_input[26730]), .B(p_input[16730]), .Z(n7268) );
  AND U10902 ( .A(p_input[6730]), .B(p_input[36730]), .Z(n7267) );
  AND U10903 ( .A(n7269), .B(n7270), .Z(o[672]) );
  AND U10904 ( .A(p_input[20672]), .B(p_input[10672]), .Z(n7270) );
  AND U10905 ( .A(p_input[672]), .B(p_input[30672]), .Z(n7269) );
  AND U10906 ( .A(n7271), .B(n7272), .Z(o[6729]) );
  AND U10907 ( .A(p_input[26729]), .B(p_input[16729]), .Z(n7272) );
  AND U10908 ( .A(p_input[6729]), .B(p_input[36729]), .Z(n7271) );
  AND U10909 ( .A(n7273), .B(n7274), .Z(o[6728]) );
  AND U10910 ( .A(p_input[26728]), .B(p_input[16728]), .Z(n7274) );
  AND U10911 ( .A(p_input[6728]), .B(p_input[36728]), .Z(n7273) );
  AND U10912 ( .A(n7275), .B(n7276), .Z(o[6727]) );
  AND U10913 ( .A(p_input[26727]), .B(p_input[16727]), .Z(n7276) );
  AND U10914 ( .A(p_input[6727]), .B(p_input[36727]), .Z(n7275) );
  AND U10915 ( .A(n7277), .B(n7278), .Z(o[6726]) );
  AND U10916 ( .A(p_input[26726]), .B(p_input[16726]), .Z(n7278) );
  AND U10917 ( .A(p_input[6726]), .B(p_input[36726]), .Z(n7277) );
  AND U10918 ( .A(n7279), .B(n7280), .Z(o[6725]) );
  AND U10919 ( .A(p_input[26725]), .B(p_input[16725]), .Z(n7280) );
  AND U10920 ( .A(p_input[6725]), .B(p_input[36725]), .Z(n7279) );
  AND U10921 ( .A(n7281), .B(n7282), .Z(o[6724]) );
  AND U10922 ( .A(p_input[26724]), .B(p_input[16724]), .Z(n7282) );
  AND U10923 ( .A(p_input[6724]), .B(p_input[36724]), .Z(n7281) );
  AND U10924 ( .A(n7283), .B(n7284), .Z(o[6723]) );
  AND U10925 ( .A(p_input[26723]), .B(p_input[16723]), .Z(n7284) );
  AND U10926 ( .A(p_input[6723]), .B(p_input[36723]), .Z(n7283) );
  AND U10927 ( .A(n7285), .B(n7286), .Z(o[6722]) );
  AND U10928 ( .A(p_input[26722]), .B(p_input[16722]), .Z(n7286) );
  AND U10929 ( .A(p_input[6722]), .B(p_input[36722]), .Z(n7285) );
  AND U10930 ( .A(n7287), .B(n7288), .Z(o[6721]) );
  AND U10931 ( .A(p_input[26721]), .B(p_input[16721]), .Z(n7288) );
  AND U10932 ( .A(p_input[6721]), .B(p_input[36721]), .Z(n7287) );
  AND U10933 ( .A(n7289), .B(n7290), .Z(o[6720]) );
  AND U10934 ( .A(p_input[26720]), .B(p_input[16720]), .Z(n7290) );
  AND U10935 ( .A(p_input[6720]), .B(p_input[36720]), .Z(n7289) );
  AND U10936 ( .A(n7291), .B(n7292), .Z(o[671]) );
  AND U10937 ( .A(p_input[20671]), .B(p_input[10671]), .Z(n7292) );
  AND U10938 ( .A(p_input[671]), .B(p_input[30671]), .Z(n7291) );
  AND U10939 ( .A(n7293), .B(n7294), .Z(o[6719]) );
  AND U10940 ( .A(p_input[26719]), .B(p_input[16719]), .Z(n7294) );
  AND U10941 ( .A(p_input[6719]), .B(p_input[36719]), .Z(n7293) );
  AND U10942 ( .A(n7295), .B(n7296), .Z(o[6718]) );
  AND U10943 ( .A(p_input[26718]), .B(p_input[16718]), .Z(n7296) );
  AND U10944 ( .A(p_input[6718]), .B(p_input[36718]), .Z(n7295) );
  AND U10945 ( .A(n7297), .B(n7298), .Z(o[6717]) );
  AND U10946 ( .A(p_input[26717]), .B(p_input[16717]), .Z(n7298) );
  AND U10947 ( .A(p_input[6717]), .B(p_input[36717]), .Z(n7297) );
  AND U10948 ( .A(n7299), .B(n7300), .Z(o[6716]) );
  AND U10949 ( .A(p_input[26716]), .B(p_input[16716]), .Z(n7300) );
  AND U10950 ( .A(p_input[6716]), .B(p_input[36716]), .Z(n7299) );
  AND U10951 ( .A(n7301), .B(n7302), .Z(o[6715]) );
  AND U10952 ( .A(p_input[26715]), .B(p_input[16715]), .Z(n7302) );
  AND U10953 ( .A(p_input[6715]), .B(p_input[36715]), .Z(n7301) );
  AND U10954 ( .A(n7303), .B(n7304), .Z(o[6714]) );
  AND U10955 ( .A(p_input[26714]), .B(p_input[16714]), .Z(n7304) );
  AND U10956 ( .A(p_input[6714]), .B(p_input[36714]), .Z(n7303) );
  AND U10957 ( .A(n7305), .B(n7306), .Z(o[6713]) );
  AND U10958 ( .A(p_input[26713]), .B(p_input[16713]), .Z(n7306) );
  AND U10959 ( .A(p_input[6713]), .B(p_input[36713]), .Z(n7305) );
  AND U10960 ( .A(n7307), .B(n7308), .Z(o[6712]) );
  AND U10961 ( .A(p_input[26712]), .B(p_input[16712]), .Z(n7308) );
  AND U10962 ( .A(p_input[6712]), .B(p_input[36712]), .Z(n7307) );
  AND U10963 ( .A(n7309), .B(n7310), .Z(o[6711]) );
  AND U10964 ( .A(p_input[26711]), .B(p_input[16711]), .Z(n7310) );
  AND U10965 ( .A(p_input[6711]), .B(p_input[36711]), .Z(n7309) );
  AND U10966 ( .A(n7311), .B(n7312), .Z(o[6710]) );
  AND U10967 ( .A(p_input[26710]), .B(p_input[16710]), .Z(n7312) );
  AND U10968 ( .A(p_input[6710]), .B(p_input[36710]), .Z(n7311) );
  AND U10969 ( .A(n7313), .B(n7314), .Z(o[670]) );
  AND U10970 ( .A(p_input[20670]), .B(p_input[10670]), .Z(n7314) );
  AND U10971 ( .A(p_input[670]), .B(p_input[30670]), .Z(n7313) );
  AND U10972 ( .A(n7315), .B(n7316), .Z(o[6709]) );
  AND U10973 ( .A(p_input[26709]), .B(p_input[16709]), .Z(n7316) );
  AND U10974 ( .A(p_input[6709]), .B(p_input[36709]), .Z(n7315) );
  AND U10975 ( .A(n7317), .B(n7318), .Z(o[6708]) );
  AND U10976 ( .A(p_input[26708]), .B(p_input[16708]), .Z(n7318) );
  AND U10977 ( .A(p_input[6708]), .B(p_input[36708]), .Z(n7317) );
  AND U10978 ( .A(n7319), .B(n7320), .Z(o[6707]) );
  AND U10979 ( .A(p_input[26707]), .B(p_input[16707]), .Z(n7320) );
  AND U10980 ( .A(p_input[6707]), .B(p_input[36707]), .Z(n7319) );
  AND U10981 ( .A(n7321), .B(n7322), .Z(o[6706]) );
  AND U10982 ( .A(p_input[26706]), .B(p_input[16706]), .Z(n7322) );
  AND U10983 ( .A(p_input[6706]), .B(p_input[36706]), .Z(n7321) );
  AND U10984 ( .A(n7323), .B(n7324), .Z(o[6705]) );
  AND U10985 ( .A(p_input[26705]), .B(p_input[16705]), .Z(n7324) );
  AND U10986 ( .A(p_input[6705]), .B(p_input[36705]), .Z(n7323) );
  AND U10987 ( .A(n7325), .B(n7326), .Z(o[6704]) );
  AND U10988 ( .A(p_input[26704]), .B(p_input[16704]), .Z(n7326) );
  AND U10989 ( .A(p_input[6704]), .B(p_input[36704]), .Z(n7325) );
  AND U10990 ( .A(n7327), .B(n7328), .Z(o[6703]) );
  AND U10991 ( .A(p_input[26703]), .B(p_input[16703]), .Z(n7328) );
  AND U10992 ( .A(p_input[6703]), .B(p_input[36703]), .Z(n7327) );
  AND U10993 ( .A(n7329), .B(n7330), .Z(o[6702]) );
  AND U10994 ( .A(p_input[26702]), .B(p_input[16702]), .Z(n7330) );
  AND U10995 ( .A(p_input[6702]), .B(p_input[36702]), .Z(n7329) );
  AND U10996 ( .A(n7331), .B(n7332), .Z(o[6701]) );
  AND U10997 ( .A(p_input[26701]), .B(p_input[16701]), .Z(n7332) );
  AND U10998 ( .A(p_input[6701]), .B(p_input[36701]), .Z(n7331) );
  AND U10999 ( .A(n7333), .B(n7334), .Z(o[6700]) );
  AND U11000 ( .A(p_input[26700]), .B(p_input[16700]), .Z(n7334) );
  AND U11001 ( .A(p_input[6700]), .B(p_input[36700]), .Z(n7333) );
  AND U11002 ( .A(n7335), .B(n7336), .Z(o[66]) );
  AND U11003 ( .A(p_input[20066]), .B(p_input[10066]), .Z(n7336) );
  AND U11004 ( .A(p_input[66]), .B(p_input[30066]), .Z(n7335) );
  AND U11005 ( .A(n7337), .B(n7338), .Z(o[669]) );
  AND U11006 ( .A(p_input[20669]), .B(p_input[10669]), .Z(n7338) );
  AND U11007 ( .A(p_input[669]), .B(p_input[30669]), .Z(n7337) );
  AND U11008 ( .A(n7339), .B(n7340), .Z(o[6699]) );
  AND U11009 ( .A(p_input[26699]), .B(p_input[16699]), .Z(n7340) );
  AND U11010 ( .A(p_input[6699]), .B(p_input[36699]), .Z(n7339) );
  AND U11011 ( .A(n7341), .B(n7342), .Z(o[6698]) );
  AND U11012 ( .A(p_input[26698]), .B(p_input[16698]), .Z(n7342) );
  AND U11013 ( .A(p_input[6698]), .B(p_input[36698]), .Z(n7341) );
  AND U11014 ( .A(n7343), .B(n7344), .Z(o[6697]) );
  AND U11015 ( .A(p_input[26697]), .B(p_input[16697]), .Z(n7344) );
  AND U11016 ( .A(p_input[6697]), .B(p_input[36697]), .Z(n7343) );
  AND U11017 ( .A(n7345), .B(n7346), .Z(o[6696]) );
  AND U11018 ( .A(p_input[26696]), .B(p_input[16696]), .Z(n7346) );
  AND U11019 ( .A(p_input[6696]), .B(p_input[36696]), .Z(n7345) );
  AND U11020 ( .A(n7347), .B(n7348), .Z(o[6695]) );
  AND U11021 ( .A(p_input[26695]), .B(p_input[16695]), .Z(n7348) );
  AND U11022 ( .A(p_input[6695]), .B(p_input[36695]), .Z(n7347) );
  AND U11023 ( .A(n7349), .B(n7350), .Z(o[6694]) );
  AND U11024 ( .A(p_input[26694]), .B(p_input[16694]), .Z(n7350) );
  AND U11025 ( .A(p_input[6694]), .B(p_input[36694]), .Z(n7349) );
  AND U11026 ( .A(n7351), .B(n7352), .Z(o[6693]) );
  AND U11027 ( .A(p_input[26693]), .B(p_input[16693]), .Z(n7352) );
  AND U11028 ( .A(p_input[6693]), .B(p_input[36693]), .Z(n7351) );
  AND U11029 ( .A(n7353), .B(n7354), .Z(o[6692]) );
  AND U11030 ( .A(p_input[26692]), .B(p_input[16692]), .Z(n7354) );
  AND U11031 ( .A(p_input[6692]), .B(p_input[36692]), .Z(n7353) );
  AND U11032 ( .A(n7355), .B(n7356), .Z(o[6691]) );
  AND U11033 ( .A(p_input[26691]), .B(p_input[16691]), .Z(n7356) );
  AND U11034 ( .A(p_input[6691]), .B(p_input[36691]), .Z(n7355) );
  AND U11035 ( .A(n7357), .B(n7358), .Z(o[6690]) );
  AND U11036 ( .A(p_input[26690]), .B(p_input[16690]), .Z(n7358) );
  AND U11037 ( .A(p_input[6690]), .B(p_input[36690]), .Z(n7357) );
  AND U11038 ( .A(n7359), .B(n7360), .Z(o[668]) );
  AND U11039 ( .A(p_input[20668]), .B(p_input[10668]), .Z(n7360) );
  AND U11040 ( .A(p_input[668]), .B(p_input[30668]), .Z(n7359) );
  AND U11041 ( .A(n7361), .B(n7362), .Z(o[6689]) );
  AND U11042 ( .A(p_input[26689]), .B(p_input[16689]), .Z(n7362) );
  AND U11043 ( .A(p_input[6689]), .B(p_input[36689]), .Z(n7361) );
  AND U11044 ( .A(n7363), .B(n7364), .Z(o[6688]) );
  AND U11045 ( .A(p_input[26688]), .B(p_input[16688]), .Z(n7364) );
  AND U11046 ( .A(p_input[6688]), .B(p_input[36688]), .Z(n7363) );
  AND U11047 ( .A(n7365), .B(n7366), .Z(o[6687]) );
  AND U11048 ( .A(p_input[26687]), .B(p_input[16687]), .Z(n7366) );
  AND U11049 ( .A(p_input[6687]), .B(p_input[36687]), .Z(n7365) );
  AND U11050 ( .A(n7367), .B(n7368), .Z(o[6686]) );
  AND U11051 ( .A(p_input[26686]), .B(p_input[16686]), .Z(n7368) );
  AND U11052 ( .A(p_input[6686]), .B(p_input[36686]), .Z(n7367) );
  AND U11053 ( .A(n7369), .B(n7370), .Z(o[6685]) );
  AND U11054 ( .A(p_input[26685]), .B(p_input[16685]), .Z(n7370) );
  AND U11055 ( .A(p_input[6685]), .B(p_input[36685]), .Z(n7369) );
  AND U11056 ( .A(n7371), .B(n7372), .Z(o[6684]) );
  AND U11057 ( .A(p_input[26684]), .B(p_input[16684]), .Z(n7372) );
  AND U11058 ( .A(p_input[6684]), .B(p_input[36684]), .Z(n7371) );
  AND U11059 ( .A(n7373), .B(n7374), .Z(o[6683]) );
  AND U11060 ( .A(p_input[26683]), .B(p_input[16683]), .Z(n7374) );
  AND U11061 ( .A(p_input[6683]), .B(p_input[36683]), .Z(n7373) );
  AND U11062 ( .A(n7375), .B(n7376), .Z(o[6682]) );
  AND U11063 ( .A(p_input[26682]), .B(p_input[16682]), .Z(n7376) );
  AND U11064 ( .A(p_input[6682]), .B(p_input[36682]), .Z(n7375) );
  AND U11065 ( .A(n7377), .B(n7378), .Z(o[6681]) );
  AND U11066 ( .A(p_input[26681]), .B(p_input[16681]), .Z(n7378) );
  AND U11067 ( .A(p_input[6681]), .B(p_input[36681]), .Z(n7377) );
  AND U11068 ( .A(n7379), .B(n7380), .Z(o[6680]) );
  AND U11069 ( .A(p_input[26680]), .B(p_input[16680]), .Z(n7380) );
  AND U11070 ( .A(p_input[6680]), .B(p_input[36680]), .Z(n7379) );
  AND U11071 ( .A(n7381), .B(n7382), .Z(o[667]) );
  AND U11072 ( .A(p_input[20667]), .B(p_input[10667]), .Z(n7382) );
  AND U11073 ( .A(p_input[667]), .B(p_input[30667]), .Z(n7381) );
  AND U11074 ( .A(n7383), .B(n7384), .Z(o[6679]) );
  AND U11075 ( .A(p_input[26679]), .B(p_input[16679]), .Z(n7384) );
  AND U11076 ( .A(p_input[6679]), .B(p_input[36679]), .Z(n7383) );
  AND U11077 ( .A(n7385), .B(n7386), .Z(o[6678]) );
  AND U11078 ( .A(p_input[26678]), .B(p_input[16678]), .Z(n7386) );
  AND U11079 ( .A(p_input[6678]), .B(p_input[36678]), .Z(n7385) );
  AND U11080 ( .A(n7387), .B(n7388), .Z(o[6677]) );
  AND U11081 ( .A(p_input[26677]), .B(p_input[16677]), .Z(n7388) );
  AND U11082 ( .A(p_input[6677]), .B(p_input[36677]), .Z(n7387) );
  AND U11083 ( .A(n7389), .B(n7390), .Z(o[6676]) );
  AND U11084 ( .A(p_input[26676]), .B(p_input[16676]), .Z(n7390) );
  AND U11085 ( .A(p_input[6676]), .B(p_input[36676]), .Z(n7389) );
  AND U11086 ( .A(n7391), .B(n7392), .Z(o[6675]) );
  AND U11087 ( .A(p_input[26675]), .B(p_input[16675]), .Z(n7392) );
  AND U11088 ( .A(p_input[6675]), .B(p_input[36675]), .Z(n7391) );
  AND U11089 ( .A(n7393), .B(n7394), .Z(o[6674]) );
  AND U11090 ( .A(p_input[26674]), .B(p_input[16674]), .Z(n7394) );
  AND U11091 ( .A(p_input[6674]), .B(p_input[36674]), .Z(n7393) );
  AND U11092 ( .A(n7395), .B(n7396), .Z(o[6673]) );
  AND U11093 ( .A(p_input[26673]), .B(p_input[16673]), .Z(n7396) );
  AND U11094 ( .A(p_input[6673]), .B(p_input[36673]), .Z(n7395) );
  AND U11095 ( .A(n7397), .B(n7398), .Z(o[6672]) );
  AND U11096 ( .A(p_input[26672]), .B(p_input[16672]), .Z(n7398) );
  AND U11097 ( .A(p_input[6672]), .B(p_input[36672]), .Z(n7397) );
  AND U11098 ( .A(n7399), .B(n7400), .Z(o[6671]) );
  AND U11099 ( .A(p_input[26671]), .B(p_input[16671]), .Z(n7400) );
  AND U11100 ( .A(p_input[6671]), .B(p_input[36671]), .Z(n7399) );
  AND U11101 ( .A(n7401), .B(n7402), .Z(o[6670]) );
  AND U11102 ( .A(p_input[26670]), .B(p_input[16670]), .Z(n7402) );
  AND U11103 ( .A(p_input[6670]), .B(p_input[36670]), .Z(n7401) );
  AND U11104 ( .A(n7403), .B(n7404), .Z(o[666]) );
  AND U11105 ( .A(p_input[20666]), .B(p_input[10666]), .Z(n7404) );
  AND U11106 ( .A(p_input[666]), .B(p_input[30666]), .Z(n7403) );
  AND U11107 ( .A(n7405), .B(n7406), .Z(o[6669]) );
  AND U11108 ( .A(p_input[26669]), .B(p_input[16669]), .Z(n7406) );
  AND U11109 ( .A(p_input[6669]), .B(p_input[36669]), .Z(n7405) );
  AND U11110 ( .A(n7407), .B(n7408), .Z(o[6668]) );
  AND U11111 ( .A(p_input[26668]), .B(p_input[16668]), .Z(n7408) );
  AND U11112 ( .A(p_input[6668]), .B(p_input[36668]), .Z(n7407) );
  AND U11113 ( .A(n7409), .B(n7410), .Z(o[6667]) );
  AND U11114 ( .A(p_input[26667]), .B(p_input[16667]), .Z(n7410) );
  AND U11115 ( .A(p_input[6667]), .B(p_input[36667]), .Z(n7409) );
  AND U11116 ( .A(n7411), .B(n7412), .Z(o[6666]) );
  AND U11117 ( .A(p_input[26666]), .B(p_input[16666]), .Z(n7412) );
  AND U11118 ( .A(p_input[6666]), .B(p_input[36666]), .Z(n7411) );
  AND U11119 ( .A(n7413), .B(n7414), .Z(o[6665]) );
  AND U11120 ( .A(p_input[26665]), .B(p_input[16665]), .Z(n7414) );
  AND U11121 ( .A(p_input[6665]), .B(p_input[36665]), .Z(n7413) );
  AND U11122 ( .A(n7415), .B(n7416), .Z(o[6664]) );
  AND U11123 ( .A(p_input[26664]), .B(p_input[16664]), .Z(n7416) );
  AND U11124 ( .A(p_input[6664]), .B(p_input[36664]), .Z(n7415) );
  AND U11125 ( .A(n7417), .B(n7418), .Z(o[6663]) );
  AND U11126 ( .A(p_input[26663]), .B(p_input[16663]), .Z(n7418) );
  AND U11127 ( .A(p_input[6663]), .B(p_input[36663]), .Z(n7417) );
  AND U11128 ( .A(n7419), .B(n7420), .Z(o[6662]) );
  AND U11129 ( .A(p_input[26662]), .B(p_input[16662]), .Z(n7420) );
  AND U11130 ( .A(p_input[6662]), .B(p_input[36662]), .Z(n7419) );
  AND U11131 ( .A(n7421), .B(n7422), .Z(o[6661]) );
  AND U11132 ( .A(p_input[26661]), .B(p_input[16661]), .Z(n7422) );
  AND U11133 ( .A(p_input[6661]), .B(p_input[36661]), .Z(n7421) );
  AND U11134 ( .A(n7423), .B(n7424), .Z(o[6660]) );
  AND U11135 ( .A(p_input[26660]), .B(p_input[16660]), .Z(n7424) );
  AND U11136 ( .A(p_input[6660]), .B(p_input[36660]), .Z(n7423) );
  AND U11137 ( .A(n7425), .B(n7426), .Z(o[665]) );
  AND U11138 ( .A(p_input[20665]), .B(p_input[10665]), .Z(n7426) );
  AND U11139 ( .A(p_input[665]), .B(p_input[30665]), .Z(n7425) );
  AND U11140 ( .A(n7427), .B(n7428), .Z(o[6659]) );
  AND U11141 ( .A(p_input[26659]), .B(p_input[16659]), .Z(n7428) );
  AND U11142 ( .A(p_input[6659]), .B(p_input[36659]), .Z(n7427) );
  AND U11143 ( .A(n7429), .B(n7430), .Z(o[6658]) );
  AND U11144 ( .A(p_input[26658]), .B(p_input[16658]), .Z(n7430) );
  AND U11145 ( .A(p_input[6658]), .B(p_input[36658]), .Z(n7429) );
  AND U11146 ( .A(n7431), .B(n7432), .Z(o[6657]) );
  AND U11147 ( .A(p_input[26657]), .B(p_input[16657]), .Z(n7432) );
  AND U11148 ( .A(p_input[6657]), .B(p_input[36657]), .Z(n7431) );
  AND U11149 ( .A(n7433), .B(n7434), .Z(o[6656]) );
  AND U11150 ( .A(p_input[26656]), .B(p_input[16656]), .Z(n7434) );
  AND U11151 ( .A(p_input[6656]), .B(p_input[36656]), .Z(n7433) );
  AND U11152 ( .A(n7435), .B(n7436), .Z(o[6655]) );
  AND U11153 ( .A(p_input[26655]), .B(p_input[16655]), .Z(n7436) );
  AND U11154 ( .A(p_input[6655]), .B(p_input[36655]), .Z(n7435) );
  AND U11155 ( .A(n7437), .B(n7438), .Z(o[6654]) );
  AND U11156 ( .A(p_input[26654]), .B(p_input[16654]), .Z(n7438) );
  AND U11157 ( .A(p_input[6654]), .B(p_input[36654]), .Z(n7437) );
  AND U11158 ( .A(n7439), .B(n7440), .Z(o[6653]) );
  AND U11159 ( .A(p_input[26653]), .B(p_input[16653]), .Z(n7440) );
  AND U11160 ( .A(p_input[6653]), .B(p_input[36653]), .Z(n7439) );
  AND U11161 ( .A(n7441), .B(n7442), .Z(o[6652]) );
  AND U11162 ( .A(p_input[26652]), .B(p_input[16652]), .Z(n7442) );
  AND U11163 ( .A(p_input[6652]), .B(p_input[36652]), .Z(n7441) );
  AND U11164 ( .A(n7443), .B(n7444), .Z(o[6651]) );
  AND U11165 ( .A(p_input[26651]), .B(p_input[16651]), .Z(n7444) );
  AND U11166 ( .A(p_input[6651]), .B(p_input[36651]), .Z(n7443) );
  AND U11167 ( .A(n7445), .B(n7446), .Z(o[6650]) );
  AND U11168 ( .A(p_input[26650]), .B(p_input[16650]), .Z(n7446) );
  AND U11169 ( .A(p_input[6650]), .B(p_input[36650]), .Z(n7445) );
  AND U11170 ( .A(n7447), .B(n7448), .Z(o[664]) );
  AND U11171 ( .A(p_input[20664]), .B(p_input[10664]), .Z(n7448) );
  AND U11172 ( .A(p_input[664]), .B(p_input[30664]), .Z(n7447) );
  AND U11173 ( .A(n7449), .B(n7450), .Z(o[6649]) );
  AND U11174 ( .A(p_input[26649]), .B(p_input[16649]), .Z(n7450) );
  AND U11175 ( .A(p_input[6649]), .B(p_input[36649]), .Z(n7449) );
  AND U11176 ( .A(n7451), .B(n7452), .Z(o[6648]) );
  AND U11177 ( .A(p_input[26648]), .B(p_input[16648]), .Z(n7452) );
  AND U11178 ( .A(p_input[6648]), .B(p_input[36648]), .Z(n7451) );
  AND U11179 ( .A(n7453), .B(n7454), .Z(o[6647]) );
  AND U11180 ( .A(p_input[26647]), .B(p_input[16647]), .Z(n7454) );
  AND U11181 ( .A(p_input[6647]), .B(p_input[36647]), .Z(n7453) );
  AND U11182 ( .A(n7455), .B(n7456), .Z(o[6646]) );
  AND U11183 ( .A(p_input[26646]), .B(p_input[16646]), .Z(n7456) );
  AND U11184 ( .A(p_input[6646]), .B(p_input[36646]), .Z(n7455) );
  AND U11185 ( .A(n7457), .B(n7458), .Z(o[6645]) );
  AND U11186 ( .A(p_input[26645]), .B(p_input[16645]), .Z(n7458) );
  AND U11187 ( .A(p_input[6645]), .B(p_input[36645]), .Z(n7457) );
  AND U11188 ( .A(n7459), .B(n7460), .Z(o[6644]) );
  AND U11189 ( .A(p_input[26644]), .B(p_input[16644]), .Z(n7460) );
  AND U11190 ( .A(p_input[6644]), .B(p_input[36644]), .Z(n7459) );
  AND U11191 ( .A(n7461), .B(n7462), .Z(o[6643]) );
  AND U11192 ( .A(p_input[26643]), .B(p_input[16643]), .Z(n7462) );
  AND U11193 ( .A(p_input[6643]), .B(p_input[36643]), .Z(n7461) );
  AND U11194 ( .A(n7463), .B(n7464), .Z(o[6642]) );
  AND U11195 ( .A(p_input[26642]), .B(p_input[16642]), .Z(n7464) );
  AND U11196 ( .A(p_input[6642]), .B(p_input[36642]), .Z(n7463) );
  AND U11197 ( .A(n7465), .B(n7466), .Z(o[6641]) );
  AND U11198 ( .A(p_input[26641]), .B(p_input[16641]), .Z(n7466) );
  AND U11199 ( .A(p_input[6641]), .B(p_input[36641]), .Z(n7465) );
  AND U11200 ( .A(n7467), .B(n7468), .Z(o[6640]) );
  AND U11201 ( .A(p_input[26640]), .B(p_input[16640]), .Z(n7468) );
  AND U11202 ( .A(p_input[6640]), .B(p_input[36640]), .Z(n7467) );
  AND U11203 ( .A(n7469), .B(n7470), .Z(o[663]) );
  AND U11204 ( .A(p_input[20663]), .B(p_input[10663]), .Z(n7470) );
  AND U11205 ( .A(p_input[663]), .B(p_input[30663]), .Z(n7469) );
  AND U11206 ( .A(n7471), .B(n7472), .Z(o[6639]) );
  AND U11207 ( .A(p_input[26639]), .B(p_input[16639]), .Z(n7472) );
  AND U11208 ( .A(p_input[6639]), .B(p_input[36639]), .Z(n7471) );
  AND U11209 ( .A(n7473), .B(n7474), .Z(o[6638]) );
  AND U11210 ( .A(p_input[26638]), .B(p_input[16638]), .Z(n7474) );
  AND U11211 ( .A(p_input[6638]), .B(p_input[36638]), .Z(n7473) );
  AND U11212 ( .A(n7475), .B(n7476), .Z(o[6637]) );
  AND U11213 ( .A(p_input[26637]), .B(p_input[16637]), .Z(n7476) );
  AND U11214 ( .A(p_input[6637]), .B(p_input[36637]), .Z(n7475) );
  AND U11215 ( .A(n7477), .B(n7478), .Z(o[6636]) );
  AND U11216 ( .A(p_input[26636]), .B(p_input[16636]), .Z(n7478) );
  AND U11217 ( .A(p_input[6636]), .B(p_input[36636]), .Z(n7477) );
  AND U11218 ( .A(n7479), .B(n7480), .Z(o[6635]) );
  AND U11219 ( .A(p_input[26635]), .B(p_input[16635]), .Z(n7480) );
  AND U11220 ( .A(p_input[6635]), .B(p_input[36635]), .Z(n7479) );
  AND U11221 ( .A(n7481), .B(n7482), .Z(o[6634]) );
  AND U11222 ( .A(p_input[26634]), .B(p_input[16634]), .Z(n7482) );
  AND U11223 ( .A(p_input[6634]), .B(p_input[36634]), .Z(n7481) );
  AND U11224 ( .A(n7483), .B(n7484), .Z(o[6633]) );
  AND U11225 ( .A(p_input[26633]), .B(p_input[16633]), .Z(n7484) );
  AND U11226 ( .A(p_input[6633]), .B(p_input[36633]), .Z(n7483) );
  AND U11227 ( .A(n7485), .B(n7486), .Z(o[6632]) );
  AND U11228 ( .A(p_input[26632]), .B(p_input[16632]), .Z(n7486) );
  AND U11229 ( .A(p_input[6632]), .B(p_input[36632]), .Z(n7485) );
  AND U11230 ( .A(n7487), .B(n7488), .Z(o[6631]) );
  AND U11231 ( .A(p_input[26631]), .B(p_input[16631]), .Z(n7488) );
  AND U11232 ( .A(p_input[6631]), .B(p_input[36631]), .Z(n7487) );
  AND U11233 ( .A(n7489), .B(n7490), .Z(o[6630]) );
  AND U11234 ( .A(p_input[26630]), .B(p_input[16630]), .Z(n7490) );
  AND U11235 ( .A(p_input[6630]), .B(p_input[36630]), .Z(n7489) );
  AND U11236 ( .A(n7491), .B(n7492), .Z(o[662]) );
  AND U11237 ( .A(p_input[20662]), .B(p_input[10662]), .Z(n7492) );
  AND U11238 ( .A(p_input[662]), .B(p_input[30662]), .Z(n7491) );
  AND U11239 ( .A(n7493), .B(n7494), .Z(o[6629]) );
  AND U11240 ( .A(p_input[26629]), .B(p_input[16629]), .Z(n7494) );
  AND U11241 ( .A(p_input[6629]), .B(p_input[36629]), .Z(n7493) );
  AND U11242 ( .A(n7495), .B(n7496), .Z(o[6628]) );
  AND U11243 ( .A(p_input[26628]), .B(p_input[16628]), .Z(n7496) );
  AND U11244 ( .A(p_input[6628]), .B(p_input[36628]), .Z(n7495) );
  AND U11245 ( .A(n7497), .B(n7498), .Z(o[6627]) );
  AND U11246 ( .A(p_input[26627]), .B(p_input[16627]), .Z(n7498) );
  AND U11247 ( .A(p_input[6627]), .B(p_input[36627]), .Z(n7497) );
  AND U11248 ( .A(n7499), .B(n7500), .Z(o[6626]) );
  AND U11249 ( .A(p_input[26626]), .B(p_input[16626]), .Z(n7500) );
  AND U11250 ( .A(p_input[6626]), .B(p_input[36626]), .Z(n7499) );
  AND U11251 ( .A(n7501), .B(n7502), .Z(o[6625]) );
  AND U11252 ( .A(p_input[26625]), .B(p_input[16625]), .Z(n7502) );
  AND U11253 ( .A(p_input[6625]), .B(p_input[36625]), .Z(n7501) );
  AND U11254 ( .A(n7503), .B(n7504), .Z(o[6624]) );
  AND U11255 ( .A(p_input[26624]), .B(p_input[16624]), .Z(n7504) );
  AND U11256 ( .A(p_input[6624]), .B(p_input[36624]), .Z(n7503) );
  AND U11257 ( .A(n7505), .B(n7506), .Z(o[6623]) );
  AND U11258 ( .A(p_input[26623]), .B(p_input[16623]), .Z(n7506) );
  AND U11259 ( .A(p_input[6623]), .B(p_input[36623]), .Z(n7505) );
  AND U11260 ( .A(n7507), .B(n7508), .Z(o[6622]) );
  AND U11261 ( .A(p_input[26622]), .B(p_input[16622]), .Z(n7508) );
  AND U11262 ( .A(p_input[6622]), .B(p_input[36622]), .Z(n7507) );
  AND U11263 ( .A(n7509), .B(n7510), .Z(o[6621]) );
  AND U11264 ( .A(p_input[26621]), .B(p_input[16621]), .Z(n7510) );
  AND U11265 ( .A(p_input[6621]), .B(p_input[36621]), .Z(n7509) );
  AND U11266 ( .A(n7511), .B(n7512), .Z(o[6620]) );
  AND U11267 ( .A(p_input[26620]), .B(p_input[16620]), .Z(n7512) );
  AND U11268 ( .A(p_input[6620]), .B(p_input[36620]), .Z(n7511) );
  AND U11269 ( .A(n7513), .B(n7514), .Z(o[661]) );
  AND U11270 ( .A(p_input[20661]), .B(p_input[10661]), .Z(n7514) );
  AND U11271 ( .A(p_input[661]), .B(p_input[30661]), .Z(n7513) );
  AND U11272 ( .A(n7515), .B(n7516), .Z(o[6619]) );
  AND U11273 ( .A(p_input[26619]), .B(p_input[16619]), .Z(n7516) );
  AND U11274 ( .A(p_input[6619]), .B(p_input[36619]), .Z(n7515) );
  AND U11275 ( .A(n7517), .B(n7518), .Z(o[6618]) );
  AND U11276 ( .A(p_input[26618]), .B(p_input[16618]), .Z(n7518) );
  AND U11277 ( .A(p_input[6618]), .B(p_input[36618]), .Z(n7517) );
  AND U11278 ( .A(n7519), .B(n7520), .Z(o[6617]) );
  AND U11279 ( .A(p_input[26617]), .B(p_input[16617]), .Z(n7520) );
  AND U11280 ( .A(p_input[6617]), .B(p_input[36617]), .Z(n7519) );
  AND U11281 ( .A(n7521), .B(n7522), .Z(o[6616]) );
  AND U11282 ( .A(p_input[26616]), .B(p_input[16616]), .Z(n7522) );
  AND U11283 ( .A(p_input[6616]), .B(p_input[36616]), .Z(n7521) );
  AND U11284 ( .A(n7523), .B(n7524), .Z(o[6615]) );
  AND U11285 ( .A(p_input[26615]), .B(p_input[16615]), .Z(n7524) );
  AND U11286 ( .A(p_input[6615]), .B(p_input[36615]), .Z(n7523) );
  AND U11287 ( .A(n7525), .B(n7526), .Z(o[6614]) );
  AND U11288 ( .A(p_input[26614]), .B(p_input[16614]), .Z(n7526) );
  AND U11289 ( .A(p_input[6614]), .B(p_input[36614]), .Z(n7525) );
  AND U11290 ( .A(n7527), .B(n7528), .Z(o[6613]) );
  AND U11291 ( .A(p_input[26613]), .B(p_input[16613]), .Z(n7528) );
  AND U11292 ( .A(p_input[6613]), .B(p_input[36613]), .Z(n7527) );
  AND U11293 ( .A(n7529), .B(n7530), .Z(o[6612]) );
  AND U11294 ( .A(p_input[26612]), .B(p_input[16612]), .Z(n7530) );
  AND U11295 ( .A(p_input[6612]), .B(p_input[36612]), .Z(n7529) );
  AND U11296 ( .A(n7531), .B(n7532), .Z(o[6611]) );
  AND U11297 ( .A(p_input[26611]), .B(p_input[16611]), .Z(n7532) );
  AND U11298 ( .A(p_input[6611]), .B(p_input[36611]), .Z(n7531) );
  AND U11299 ( .A(n7533), .B(n7534), .Z(o[6610]) );
  AND U11300 ( .A(p_input[26610]), .B(p_input[16610]), .Z(n7534) );
  AND U11301 ( .A(p_input[6610]), .B(p_input[36610]), .Z(n7533) );
  AND U11302 ( .A(n7535), .B(n7536), .Z(o[660]) );
  AND U11303 ( .A(p_input[20660]), .B(p_input[10660]), .Z(n7536) );
  AND U11304 ( .A(p_input[660]), .B(p_input[30660]), .Z(n7535) );
  AND U11305 ( .A(n7537), .B(n7538), .Z(o[6609]) );
  AND U11306 ( .A(p_input[26609]), .B(p_input[16609]), .Z(n7538) );
  AND U11307 ( .A(p_input[6609]), .B(p_input[36609]), .Z(n7537) );
  AND U11308 ( .A(n7539), .B(n7540), .Z(o[6608]) );
  AND U11309 ( .A(p_input[26608]), .B(p_input[16608]), .Z(n7540) );
  AND U11310 ( .A(p_input[6608]), .B(p_input[36608]), .Z(n7539) );
  AND U11311 ( .A(n7541), .B(n7542), .Z(o[6607]) );
  AND U11312 ( .A(p_input[26607]), .B(p_input[16607]), .Z(n7542) );
  AND U11313 ( .A(p_input[6607]), .B(p_input[36607]), .Z(n7541) );
  AND U11314 ( .A(n7543), .B(n7544), .Z(o[6606]) );
  AND U11315 ( .A(p_input[26606]), .B(p_input[16606]), .Z(n7544) );
  AND U11316 ( .A(p_input[6606]), .B(p_input[36606]), .Z(n7543) );
  AND U11317 ( .A(n7545), .B(n7546), .Z(o[6605]) );
  AND U11318 ( .A(p_input[26605]), .B(p_input[16605]), .Z(n7546) );
  AND U11319 ( .A(p_input[6605]), .B(p_input[36605]), .Z(n7545) );
  AND U11320 ( .A(n7547), .B(n7548), .Z(o[6604]) );
  AND U11321 ( .A(p_input[26604]), .B(p_input[16604]), .Z(n7548) );
  AND U11322 ( .A(p_input[6604]), .B(p_input[36604]), .Z(n7547) );
  AND U11323 ( .A(n7549), .B(n7550), .Z(o[6603]) );
  AND U11324 ( .A(p_input[26603]), .B(p_input[16603]), .Z(n7550) );
  AND U11325 ( .A(p_input[6603]), .B(p_input[36603]), .Z(n7549) );
  AND U11326 ( .A(n7551), .B(n7552), .Z(o[6602]) );
  AND U11327 ( .A(p_input[26602]), .B(p_input[16602]), .Z(n7552) );
  AND U11328 ( .A(p_input[6602]), .B(p_input[36602]), .Z(n7551) );
  AND U11329 ( .A(n7553), .B(n7554), .Z(o[6601]) );
  AND U11330 ( .A(p_input[26601]), .B(p_input[16601]), .Z(n7554) );
  AND U11331 ( .A(p_input[6601]), .B(p_input[36601]), .Z(n7553) );
  AND U11332 ( .A(n7555), .B(n7556), .Z(o[6600]) );
  AND U11333 ( .A(p_input[26600]), .B(p_input[16600]), .Z(n7556) );
  AND U11334 ( .A(p_input[6600]), .B(p_input[36600]), .Z(n7555) );
  AND U11335 ( .A(n7557), .B(n7558), .Z(o[65]) );
  AND U11336 ( .A(p_input[20065]), .B(p_input[10065]), .Z(n7558) );
  AND U11337 ( .A(p_input[65]), .B(p_input[30065]), .Z(n7557) );
  AND U11338 ( .A(n7559), .B(n7560), .Z(o[659]) );
  AND U11339 ( .A(p_input[20659]), .B(p_input[10659]), .Z(n7560) );
  AND U11340 ( .A(p_input[659]), .B(p_input[30659]), .Z(n7559) );
  AND U11341 ( .A(n7561), .B(n7562), .Z(o[6599]) );
  AND U11342 ( .A(p_input[26599]), .B(p_input[16599]), .Z(n7562) );
  AND U11343 ( .A(p_input[6599]), .B(p_input[36599]), .Z(n7561) );
  AND U11344 ( .A(n7563), .B(n7564), .Z(o[6598]) );
  AND U11345 ( .A(p_input[26598]), .B(p_input[16598]), .Z(n7564) );
  AND U11346 ( .A(p_input[6598]), .B(p_input[36598]), .Z(n7563) );
  AND U11347 ( .A(n7565), .B(n7566), .Z(o[6597]) );
  AND U11348 ( .A(p_input[26597]), .B(p_input[16597]), .Z(n7566) );
  AND U11349 ( .A(p_input[6597]), .B(p_input[36597]), .Z(n7565) );
  AND U11350 ( .A(n7567), .B(n7568), .Z(o[6596]) );
  AND U11351 ( .A(p_input[26596]), .B(p_input[16596]), .Z(n7568) );
  AND U11352 ( .A(p_input[6596]), .B(p_input[36596]), .Z(n7567) );
  AND U11353 ( .A(n7569), .B(n7570), .Z(o[6595]) );
  AND U11354 ( .A(p_input[26595]), .B(p_input[16595]), .Z(n7570) );
  AND U11355 ( .A(p_input[6595]), .B(p_input[36595]), .Z(n7569) );
  AND U11356 ( .A(n7571), .B(n7572), .Z(o[6594]) );
  AND U11357 ( .A(p_input[26594]), .B(p_input[16594]), .Z(n7572) );
  AND U11358 ( .A(p_input[6594]), .B(p_input[36594]), .Z(n7571) );
  AND U11359 ( .A(n7573), .B(n7574), .Z(o[6593]) );
  AND U11360 ( .A(p_input[26593]), .B(p_input[16593]), .Z(n7574) );
  AND U11361 ( .A(p_input[6593]), .B(p_input[36593]), .Z(n7573) );
  AND U11362 ( .A(n7575), .B(n7576), .Z(o[6592]) );
  AND U11363 ( .A(p_input[26592]), .B(p_input[16592]), .Z(n7576) );
  AND U11364 ( .A(p_input[6592]), .B(p_input[36592]), .Z(n7575) );
  AND U11365 ( .A(n7577), .B(n7578), .Z(o[6591]) );
  AND U11366 ( .A(p_input[26591]), .B(p_input[16591]), .Z(n7578) );
  AND U11367 ( .A(p_input[6591]), .B(p_input[36591]), .Z(n7577) );
  AND U11368 ( .A(n7579), .B(n7580), .Z(o[6590]) );
  AND U11369 ( .A(p_input[26590]), .B(p_input[16590]), .Z(n7580) );
  AND U11370 ( .A(p_input[6590]), .B(p_input[36590]), .Z(n7579) );
  AND U11371 ( .A(n7581), .B(n7582), .Z(o[658]) );
  AND U11372 ( .A(p_input[20658]), .B(p_input[10658]), .Z(n7582) );
  AND U11373 ( .A(p_input[658]), .B(p_input[30658]), .Z(n7581) );
  AND U11374 ( .A(n7583), .B(n7584), .Z(o[6589]) );
  AND U11375 ( .A(p_input[26589]), .B(p_input[16589]), .Z(n7584) );
  AND U11376 ( .A(p_input[6589]), .B(p_input[36589]), .Z(n7583) );
  AND U11377 ( .A(n7585), .B(n7586), .Z(o[6588]) );
  AND U11378 ( .A(p_input[26588]), .B(p_input[16588]), .Z(n7586) );
  AND U11379 ( .A(p_input[6588]), .B(p_input[36588]), .Z(n7585) );
  AND U11380 ( .A(n7587), .B(n7588), .Z(o[6587]) );
  AND U11381 ( .A(p_input[26587]), .B(p_input[16587]), .Z(n7588) );
  AND U11382 ( .A(p_input[6587]), .B(p_input[36587]), .Z(n7587) );
  AND U11383 ( .A(n7589), .B(n7590), .Z(o[6586]) );
  AND U11384 ( .A(p_input[26586]), .B(p_input[16586]), .Z(n7590) );
  AND U11385 ( .A(p_input[6586]), .B(p_input[36586]), .Z(n7589) );
  AND U11386 ( .A(n7591), .B(n7592), .Z(o[6585]) );
  AND U11387 ( .A(p_input[26585]), .B(p_input[16585]), .Z(n7592) );
  AND U11388 ( .A(p_input[6585]), .B(p_input[36585]), .Z(n7591) );
  AND U11389 ( .A(n7593), .B(n7594), .Z(o[6584]) );
  AND U11390 ( .A(p_input[26584]), .B(p_input[16584]), .Z(n7594) );
  AND U11391 ( .A(p_input[6584]), .B(p_input[36584]), .Z(n7593) );
  AND U11392 ( .A(n7595), .B(n7596), .Z(o[6583]) );
  AND U11393 ( .A(p_input[26583]), .B(p_input[16583]), .Z(n7596) );
  AND U11394 ( .A(p_input[6583]), .B(p_input[36583]), .Z(n7595) );
  AND U11395 ( .A(n7597), .B(n7598), .Z(o[6582]) );
  AND U11396 ( .A(p_input[26582]), .B(p_input[16582]), .Z(n7598) );
  AND U11397 ( .A(p_input[6582]), .B(p_input[36582]), .Z(n7597) );
  AND U11398 ( .A(n7599), .B(n7600), .Z(o[6581]) );
  AND U11399 ( .A(p_input[26581]), .B(p_input[16581]), .Z(n7600) );
  AND U11400 ( .A(p_input[6581]), .B(p_input[36581]), .Z(n7599) );
  AND U11401 ( .A(n7601), .B(n7602), .Z(o[6580]) );
  AND U11402 ( .A(p_input[26580]), .B(p_input[16580]), .Z(n7602) );
  AND U11403 ( .A(p_input[6580]), .B(p_input[36580]), .Z(n7601) );
  AND U11404 ( .A(n7603), .B(n7604), .Z(o[657]) );
  AND U11405 ( .A(p_input[20657]), .B(p_input[10657]), .Z(n7604) );
  AND U11406 ( .A(p_input[657]), .B(p_input[30657]), .Z(n7603) );
  AND U11407 ( .A(n7605), .B(n7606), .Z(o[6579]) );
  AND U11408 ( .A(p_input[26579]), .B(p_input[16579]), .Z(n7606) );
  AND U11409 ( .A(p_input[6579]), .B(p_input[36579]), .Z(n7605) );
  AND U11410 ( .A(n7607), .B(n7608), .Z(o[6578]) );
  AND U11411 ( .A(p_input[26578]), .B(p_input[16578]), .Z(n7608) );
  AND U11412 ( .A(p_input[6578]), .B(p_input[36578]), .Z(n7607) );
  AND U11413 ( .A(n7609), .B(n7610), .Z(o[6577]) );
  AND U11414 ( .A(p_input[26577]), .B(p_input[16577]), .Z(n7610) );
  AND U11415 ( .A(p_input[6577]), .B(p_input[36577]), .Z(n7609) );
  AND U11416 ( .A(n7611), .B(n7612), .Z(o[6576]) );
  AND U11417 ( .A(p_input[26576]), .B(p_input[16576]), .Z(n7612) );
  AND U11418 ( .A(p_input[6576]), .B(p_input[36576]), .Z(n7611) );
  AND U11419 ( .A(n7613), .B(n7614), .Z(o[6575]) );
  AND U11420 ( .A(p_input[26575]), .B(p_input[16575]), .Z(n7614) );
  AND U11421 ( .A(p_input[6575]), .B(p_input[36575]), .Z(n7613) );
  AND U11422 ( .A(n7615), .B(n7616), .Z(o[6574]) );
  AND U11423 ( .A(p_input[26574]), .B(p_input[16574]), .Z(n7616) );
  AND U11424 ( .A(p_input[6574]), .B(p_input[36574]), .Z(n7615) );
  AND U11425 ( .A(n7617), .B(n7618), .Z(o[6573]) );
  AND U11426 ( .A(p_input[26573]), .B(p_input[16573]), .Z(n7618) );
  AND U11427 ( .A(p_input[6573]), .B(p_input[36573]), .Z(n7617) );
  AND U11428 ( .A(n7619), .B(n7620), .Z(o[6572]) );
  AND U11429 ( .A(p_input[26572]), .B(p_input[16572]), .Z(n7620) );
  AND U11430 ( .A(p_input[6572]), .B(p_input[36572]), .Z(n7619) );
  AND U11431 ( .A(n7621), .B(n7622), .Z(o[6571]) );
  AND U11432 ( .A(p_input[26571]), .B(p_input[16571]), .Z(n7622) );
  AND U11433 ( .A(p_input[6571]), .B(p_input[36571]), .Z(n7621) );
  AND U11434 ( .A(n7623), .B(n7624), .Z(o[6570]) );
  AND U11435 ( .A(p_input[26570]), .B(p_input[16570]), .Z(n7624) );
  AND U11436 ( .A(p_input[6570]), .B(p_input[36570]), .Z(n7623) );
  AND U11437 ( .A(n7625), .B(n7626), .Z(o[656]) );
  AND U11438 ( .A(p_input[20656]), .B(p_input[10656]), .Z(n7626) );
  AND U11439 ( .A(p_input[656]), .B(p_input[30656]), .Z(n7625) );
  AND U11440 ( .A(n7627), .B(n7628), .Z(o[6569]) );
  AND U11441 ( .A(p_input[26569]), .B(p_input[16569]), .Z(n7628) );
  AND U11442 ( .A(p_input[6569]), .B(p_input[36569]), .Z(n7627) );
  AND U11443 ( .A(n7629), .B(n7630), .Z(o[6568]) );
  AND U11444 ( .A(p_input[26568]), .B(p_input[16568]), .Z(n7630) );
  AND U11445 ( .A(p_input[6568]), .B(p_input[36568]), .Z(n7629) );
  AND U11446 ( .A(n7631), .B(n7632), .Z(o[6567]) );
  AND U11447 ( .A(p_input[26567]), .B(p_input[16567]), .Z(n7632) );
  AND U11448 ( .A(p_input[6567]), .B(p_input[36567]), .Z(n7631) );
  AND U11449 ( .A(n7633), .B(n7634), .Z(o[6566]) );
  AND U11450 ( .A(p_input[26566]), .B(p_input[16566]), .Z(n7634) );
  AND U11451 ( .A(p_input[6566]), .B(p_input[36566]), .Z(n7633) );
  AND U11452 ( .A(n7635), .B(n7636), .Z(o[6565]) );
  AND U11453 ( .A(p_input[26565]), .B(p_input[16565]), .Z(n7636) );
  AND U11454 ( .A(p_input[6565]), .B(p_input[36565]), .Z(n7635) );
  AND U11455 ( .A(n7637), .B(n7638), .Z(o[6564]) );
  AND U11456 ( .A(p_input[26564]), .B(p_input[16564]), .Z(n7638) );
  AND U11457 ( .A(p_input[6564]), .B(p_input[36564]), .Z(n7637) );
  AND U11458 ( .A(n7639), .B(n7640), .Z(o[6563]) );
  AND U11459 ( .A(p_input[26563]), .B(p_input[16563]), .Z(n7640) );
  AND U11460 ( .A(p_input[6563]), .B(p_input[36563]), .Z(n7639) );
  AND U11461 ( .A(n7641), .B(n7642), .Z(o[6562]) );
  AND U11462 ( .A(p_input[26562]), .B(p_input[16562]), .Z(n7642) );
  AND U11463 ( .A(p_input[6562]), .B(p_input[36562]), .Z(n7641) );
  AND U11464 ( .A(n7643), .B(n7644), .Z(o[6561]) );
  AND U11465 ( .A(p_input[26561]), .B(p_input[16561]), .Z(n7644) );
  AND U11466 ( .A(p_input[6561]), .B(p_input[36561]), .Z(n7643) );
  AND U11467 ( .A(n7645), .B(n7646), .Z(o[6560]) );
  AND U11468 ( .A(p_input[26560]), .B(p_input[16560]), .Z(n7646) );
  AND U11469 ( .A(p_input[6560]), .B(p_input[36560]), .Z(n7645) );
  AND U11470 ( .A(n7647), .B(n7648), .Z(o[655]) );
  AND U11471 ( .A(p_input[20655]), .B(p_input[10655]), .Z(n7648) );
  AND U11472 ( .A(p_input[655]), .B(p_input[30655]), .Z(n7647) );
  AND U11473 ( .A(n7649), .B(n7650), .Z(o[6559]) );
  AND U11474 ( .A(p_input[26559]), .B(p_input[16559]), .Z(n7650) );
  AND U11475 ( .A(p_input[6559]), .B(p_input[36559]), .Z(n7649) );
  AND U11476 ( .A(n7651), .B(n7652), .Z(o[6558]) );
  AND U11477 ( .A(p_input[26558]), .B(p_input[16558]), .Z(n7652) );
  AND U11478 ( .A(p_input[6558]), .B(p_input[36558]), .Z(n7651) );
  AND U11479 ( .A(n7653), .B(n7654), .Z(o[6557]) );
  AND U11480 ( .A(p_input[26557]), .B(p_input[16557]), .Z(n7654) );
  AND U11481 ( .A(p_input[6557]), .B(p_input[36557]), .Z(n7653) );
  AND U11482 ( .A(n7655), .B(n7656), .Z(o[6556]) );
  AND U11483 ( .A(p_input[26556]), .B(p_input[16556]), .Z(n7656) );
  AND U11484 ( .A(p_input[6556]), .B(p_input[36556]), .Z(n7655) );
  AND U11485 ( .A(n7657), .B(n7658), .Z(o[6555]) );
  AND U11486 ( .A(p_input[26555]), .B(p_input[16555]), .Z(n7658) );
  AND U11487 ( .A(p_input[6555]), .B(p_input[36555]), .Z(n7657) );
  AND U11488 ( .A(n7659), .B(n7660), .Z(o[6554]) );
  AND U11489 ( .A(p_input[26554]), .B(p_input[16554]), .Z(n7660) );
  AND U11490 ( .A(p_input[6554]), .B(p_input[36554]), .Z(n7659) );
  AND U11491 ( .A(n7661), .B(n7662), .Z(o[6553]) );
  AND U11492 ( .A(p_input[26553]), .B(p_input[16553]), .Z(n7662) );
  AND U11493 ( .A(p_input[6553]), .B(p_input[36553]), .Z(n7661) );
  AND U11494 ( .A(n7663), .B(n7664), .Z(o[6552]) );
  AND U11495 ( .A(p_input[26552]), .B(p_input[16552]), .Z(n7664) );
  AND U11496 ( .A(p_input[6552]), .B(p_input[36552]), .Z(n7663) );
  AND U11497 ( .A(n7665), .B(n7666), .Z(o[6551]) );
  AND U11498 ( .A(p_input[26551]), .B(p_input[16551]), .Z(n7666) );
  AND U11499 ( .A(p_input[6551]), .B(p_input[36551]), .Z(n7665) );
  AND U11500 ( .A(n7667), .B(n7668), .Z(o[6550]) );
  AND U11501 ( .A(p_input[26550]), .B(p_input[16550]), .Z(n7668) );
  AND U11502 ( .A(p_input[6550]), .B(p_input[36550]), .Z(n7667) );
  AND U11503 ( .A(n7669), .B(n7670), .Z(o[654]) );
  AND U11504 ( .A(p_input[20654]), .B(p_input[10654]), .Z(n7670) );
  AND U11505 ( .A(p_input[654]), .B(p_input[30654]), .Z(n7669) );
  AND U11506 ( .A(n7671), .B(n7672), .Z(o[6549]) );
  AND U11507 ( .A(p_input[26549]), .B(p_input[16549]), .Z(n7672) );
  AND U11508 ( .A(p_input[6549]), .B(p_input[36549]), .Z(n7671) );
  AND U11509 ( .A(n7673), .B(n7674), .Z(o[6548]) );
  AND U11510 ( .A(p_input[26548]), .B(p_input[16548]), .Z(n7674) );
  AND U11511 ( .A(p_input[6548]), .B(p_input[36548]), .Z(n7673) );
  AND U11512 ( .A(n7675), .B(n7676), .Z(o[6547]) );
  AND U11513 ( .A(p_input[26547]), .B(p_input[16547]), .Z(n7676) );
  AND U11514 ( .A(p_input[6547]), .B(p_input[36547]), .Z(n7675) );
  AND U11515 ( .A(n7677), .B(n7678), .Z(o[6546]) );
  AND U11516 ( .A(p_input[26546]), .B(p_input[16546]), .Z(n7678) );
  AND U11517 ( .A(p_input[6546]), .B(p_input[36546]), .Z(n7677) );
  AND U11518 ( .A(n7679), .B(n7680), .Z(o[6545]) );
  AND U11519 ( .A(p_input[26545]), .B(p_input[16545]), .Z(n7680) );
  AND U11520 ( .A(p_input[6545]), .B(p_input[36545]), .Z(n7679) );
  AND U11521 ( .A(n7681), .B(n7682), .Z(o[6544]) );
  AND U11522 ( .A(p_input[26544]), .B(p_input[16544]), .Z(n7682) );
  AND U11523 ( .A(p_input[6544]), .B(p_input[36544]), .Z(n7681) );
  AND U11524 ( .A(n7683), .B(n7684), .Z(o[6543]) );
  AND U11525 ( .A(p_input[26543]), .B(p_input[16543]), .Z(n7684) );
  AND U11526 ( .A(p_input[6543]), .B(p_input[36543]), .Z(n7683) );
  AND U11527 ( .A(n7685), .B(n7686), .Z(o[6542]) );
  AND U11528 ( .A(p_input[26542]), .B(p_input[16542]), .Z(n7686) );
  AND U11529 ( .A(p_input[6542]), .B(p_input[36542]), .Z(n7685) );
  AND U11530 ( .A(n7687), .B(n7688), .Z(o[6541]) );
  AND U11531 ( .A(p_input[26541]), .B(p_input[16541]), .Z(n7688) );
  AND U11532 ( .A(p_input[6541]), .B(p_input[36541]), .Z(n7687) );
  AND U11533 ( .A(n7689), .B(n7690), .Z(o[6540]) );
  AND U11534 ( .A(p_input[26540]), .B(p_input[16540]), .Z(n7690) );
  AND U11535 ( .A(p_input[6540]), .B(p_input[36540]), .Z(n7689) );
  AND U11536 ( .A(n7691), .B(n7692), .Z(o[653]) );
  AND U11537 ( .A(p_input[20653]), .B(p_input[10653]), .Z(n7692) );
  AND U11538 ( .A(p_input[653]), .B(p_input[30653]), .Z(n7691) );
  AND U11539 ( .A(n7693), .B(n7694), .Z(o[6539]) );
  AND U11540 ( .A(p_input[26539]), .B(p_input[16539]), .Z(n7694) );
  AND U11541 ( .A(p_input[6539]), .B(p_input[36539]), .Z(n7693) );
  AND U11542 ( .A(n7695), .B(n7696), .Z(o[6538]) );
  AND U11543 ( .A(p_input[26538]), .B(p_input[16538]), .Z(n7696) );
  AND U11544 ( .A(p_input[6538]), .B(p_input[36538]), .Z(n7695) );
  AND U11545 ( .A(n7697), .B(n7698), .Z(o[6537]) );
  AND U11546 ( .A(p_input[26537]), .B(p_input[16537]), .Z(n7698) );
  AND U11547 ( .A(p_input[6537]), .B(p_input[36537]), .Z(n7697) );
  AND U11548 ( .A(n7699), .B(n7700), .Z(o[6536]) );
  AND U11549 ( .A(p_input[26536]), .B(p_input[16536]), .Z(n7700) );
  AND U11550 ( .A(p_input[6536]), .B(p_input[36536]), .Z(n7699) );
  AND U11551 ( .A(n7701), .B(n7702), .Z(o[6535]) );
  AND U11552 ( .A(p_input[26535]), .B(p_input[16535]), .Z(n7702) );
  AND U11553 ( .A(p_input[6535]), .B(p_input[36535]), .Z(n7701) );
  AND U11554 ( .A(n7703), .B(n7704), .Z(o[6534]) );
  AND U11555 ( .A(p_input[26534]), .B(p_input[16534]), .Z(n7704) );
  AND U11556 ( .A(p_input[6534]), .B(p_input[36534]), .Z(n7703) );
  AND U11557 ( .A(n7705), .B(n7706), .Z(o[6533]) );
  AND U11558 ( .A(p_input[26533]), .B(p_input[16533]), .Z(n7706) );
  AND U11559 ( .A(p_input[6533]), .B(p_input[36533]), .Z(n7705) );
  AND U11560 ( .A(n7707), .B(n7708), .Z(o[6532]) );
  AND U11561 ( .A(p_input[26532]), .B(p_input[16532]), .Z(n7708) );
  AND U11562 ( .A(p_input[6532]), .B(p_input[36532]), .Z(n7707) );
  AND U11563 ( .A(n7709), .B(n7710), .Z(o[6531]) );
  AND U11564 ( .A(p_input[26531]), .B(p_input[16531]), .Z(n7710) );
  AND U11565 ( .A(p_input[6531]), .B(p_input[36531]), .Z(n7709) );
  AND U11566 ( .A(n7711), .B(n7712), .Z(o[6530]) );
  AND U11567 ( .A(p_input[26530]), .B(p_input[16530]), .Z(n7712) );
  AND U11568 ( .A(p_input[6530]), .B(p_input[36530]), .Z(n7711) );
  AND U11569 ( .A(n7713), .B(n7714), .Z(o[652]) );
  AND U11570 ( .A(p_input[20652]), .B(p_input[10652]), .Z(n7714) );
  AND U11571 ( .A(p_input[652]), .B(p_input[30652]), .Z(n7713) );
  AND U11572 ( .A(n7715), .B(n7716), .Z(o[6529]) );
  AND U11573 ( .A(p_input[26529]), .B(p_input[16529]), .Z(n7716) );
  AND U11574 ( .A(p_input[6529]), .B(p_input[36529]), .Z(n7715) );
  AND U11575 ( .A(n7717), .B(n7718), .Z(o[6528]) );
  AND U11576 ( .A(p_input[26528]), .B(p_input[16528]), .Z(n7718) );
  AND U11577 ( .A(p_input[6528]), .B(p_input[36528]), .Z(n7717) );
  AND U11578 ( .A(n7719), .B(n7720), .Z(o[6527]) );
  AND U11579 ( .A(p_input[26527]), .B(p_input[16527]), .Z(n7720) );
  AND U11580 ( .A(p_input[6527]), .B(p_input[36527]), .Z(n7719) );
  AND U11581 ( .A(n7721), .B(n7722), .Z(o[6526]) );
  AND U11582 ( .A(p_input[26526]), .B(p_input[16526]), .Z(n7722) );
  AND U11583 ( .A(p_input[6526]), .B(p_input[36526]), .Z(n7721) );
  AND U11584 ( .A(n7723), .B(n7724), .Z(o[6525]) );
  AND U11585 ( .A(p_input[26525]), .B(p_input[16525]), .Z(n7724) );
  AND U11586 ( .A(p_input[6525]), .B(p_input[36525]), .Z(n7723) );
  AND U11587 ( .A(n7725), .B(n7726), .Z(o[6524]) );
  AND U11588 ( .A(p_input[26524]), .B(p_input[16524]), .Z(n7726) );
  AND U11589 ( .A(p_input[6524]), .B(p_input[36524]), .Z(n7725) );
  AND U11590 ( .A(n7727), .B(n7728), .Z(o[6523]) );
  AND U11591 ( .A(p_input[26523]), .B(p_input[16523]), .Z(n7728) );
  AND U11592 ( .A(p_input[6523]), .B(p_input[36523]), .Z(n7727) );
  AND U11593 ( .A(n7729), .B(n7730), .Z(o[6522]) );
  AND U11594 ( .A(p_input[26522]), .B(p_input[16522]), .Z(n7730) );
  AND U11595 ( .A(p_input[6522]), .B(p_input[36522]), .Z(n7729) );
  AND U11596 ( .A(n7731), .B(n7732), .Z(o[6521]) );
  AND U11597 ( .A(p_input[26521]), .B(p_input[16521]), .Z(n7732) );
  AND U11598 ( .A(p_input[6521]), .B(p_input[36521]), .Z(n7731) );
  AND U11599 ( .A(n7733), .B(n7734), .Z(o[6520]) );
  AND U11600 ( .A(p_input[26520]), .B(p_input[16520]), .Z(n7734) );
  AND U11601 ( .A(p_input[6520]), .B(p_input[36520]), .Z(n7733) );
  AND U11602 ( .A(n7735), .B(n7736), .Z(o[651]) );
  AND U11603 ( .A(p_input[20651]), .B(p_input[10651]), .Z(n7736) );
  AND U11604 ( .A(p_input[651]), .B(p_input[30651]), .Z(n7735) );
  AND U11605 ( .A(n7737), .B(n7738), .Z(o[6519]) );
  AND U11606 ( .A(p_input[26519]), .B(p_input[16519]), .Z(n7738) );
  AND U11607 ( .A(p_input[6519]), .B(p_input[36519]), .Z(n7737) );
  AND U11608 ( .A(n7739), .B(n7740), .Z(o[6518]) );
  AND U11609 ( .A(p_input[26518]), .B(p_input[16518]), .Z(n7740) );
  AND U11610 ( .A(p_input[6518]), .B(p_input[36518]), .Z(n7739) );
  AND U11611 ( .A(n7741), .B(n7742), .Z(o[6517]) );
  AND U11612 ( .A(p_input[26517]), .B(p_input[16517]), .Z(n7742) );
  AND U11613 ( .A(p_input[6517]), .B(p_input[36517]), .Z(n7741) );
  AND U11614 ( .A(n7743), .B(n7744), .Z(o[6516]) );
  AND U11615 ( .A(p_input[26516]), .B(p_input[16516]), .Z(n7744) );
  AND U11616 ( .A(p_input[6516]), .B(p_input[36516]), .Z(n7743) );
  AND U11617 ( .A(n7745), .B(n7746), .Z(o[6515]) );
  AND U11618 ( .A(p_input[26515]), .B(p_input[16515]), .Z(n7746) );
  AND U11619 ( .A(p_input[6515]), .B(p_input[36515]), .Z(n7745) );
  AND U11620 ( .A(n7747), .B(n7748), .Z(o[6514]) );
  AND U11621 ( .A(p_input[26514]), .B(p_input[16514]), .Z(n7748) );
  AND U11622 ( .A(p_input[6514]), .B(p_input[36514]), .Z(n7747) );
  AND U11623 ( .A(n7749), .B(n7750), .Z(o[6513]) );
  AND U11624 ( .A(p_input[26513]), .B(p_input[16513]), .Z(n7750) );
  AND U11625 ( .A(p_input[6513]), .B(p_input[36513]), .Z(n7749) );
  AND U11626 ( .A(n7751), .B(n7752), .Z(o[6512]) );
  AND U11627 ( .A(p_input[26512]), .B(p_input[16512]), .Z(n7752) );
  AND U11628 ( .A(p_input[6512]), .B(p_input[36512]), .Z(n7751) );
  AND U11629 ( .A(n7753), .B(n7754), .Z(o[6511]) );
  AND U11630 ( .A(p_input[26511]), .B(p_input[16511]), .Z(n7754) );
  AND U11631 ( .A(p_input[6511]), .B(p_input[36511]), .Z(n7753) );
  AND U11632 ( .A(n7755), .B(n7756), .Z(o[6510]) );
  AND U11633 ( .A(p_input[26510]), .B(p_input[16510]), .Z(n7756) );
  AND U11634 ( .A(p_input[6510]), .B(p_input[36510]), .Z(n7755) );
  AND U11635 ( .A(n7757), .B(n7758), .Z(o[650]) );
  AND U11636 ( .A(p_input[20650]), .B(p_input[10650]), .Z(n7758) );
  AND U11637 ( .A(p_input[650]), .B(p_input[30650]), .Z(n7757) );
  AND U11638 ( .A(n7759), .B(n7760), .Z(o[6509]) );
  AND U11639 ( .A(p_input[26509]), .B(p_input[16509]), .Z(n7760) );
  AND U11640 ( .A(p_input[6509]), .B(p_input[36509]), .Z(n7759) );
  AND U11641 ( .A(n7761), .B(n7762), .Z(o[6508]) );
  AND U11642 ( .A(p_input[26508]), .B(p_input[16508]), .Z(n7762) );
  AND U11643 ( .A(p_input[6508]), .B(p_input[36508]), .Z(n7761) );
  AND U11644 ( .A(n7763), .B(n7764), .Z(o[6507]) );
  AND U11645 ( .A(p_input[26507]), .B(p_input[16507]), .Z(n7764) );
  AND U11646 ( .A(p_input[6507]), .B(p_input[36507]), .Z(n7763) );
  AND U11647 ( .A(n7765), .B(n7766), .Z(o[6506]) );
  AND U11648 ( .A(p_input[26506]), .B(p_input[16506]), .Z(n7766) );
  AND U11649 ( .A(p_input[6506]), .B(p_input[36506]), .Z(n7765) );
  AND U11650 ( .A(n7767), .B(n7768), .Z(o[6505]) );
  AND U11651 ( .A(p_input[26505]), .B(p_input[16505]), .Z(n7768) );
  AND U11652 ( .A(p_input[6505]), .B(p_input[36505]), .Z(n7767) );
  AND U11653 ( .A(n7769), .B(n7770), .Z(o[6504]) );
  AND U11654 ( .A(p_input[26504]), .B(p_input[16504]), .Z(n7770) );
  AND U11655 ( .A(p_input[6504]), .B(p_input[36504]), .Z(n7769) );
  AND U11656 ( .A(n7771), .B(n7772), .Z(o[6503]) );
  AND U11657 ( .A(p_input[26503]), .B(p_input[16503]), .Z(n7772) );
  AND U11658 ( .A(p_input[6503]), .B(p_input[36503]), .Z(n7771) );
  AND U11659 ( .A(n7773), .B(n7774), .Z(o[6502]) );
  AND U11660 ( .A(p_input[26502]), .B(p_input[16502]), .Z(n7774) );
  AND U11661 ( .A(p_input[6502]), .B(p_input[36502]), .Z(n7773) );
  AND U11662 ( .A(n7775), .B(n7776), .Z(o[6501]) );
  AND U11663 ( .A(p_input[26501]), .B(p_input[16501]), .Z(n7776) );
  AND U11664 ( .A(p_input[6501]), .B(p_input[36501]), .Z(n7775) );
  AND U11665 ( .A(n7777), .B(n7778), .Z(o[6500]) );
  AND U11666 ( .A(p_input[26500]), .B(p_input[16500]), .Z(n7778) );
  AND U11667 ( .A(p_input[6500]), .B(p_input[36500]), .Z(n7777) );
  AND U11668 ( .A(n7779), .B(n7780), .Z(o[64]) );
  AND U11669 ( .A(p_input[20064]), .B(p_input[10064]), .Z(n7780) );
  AND U11670 ( .A(p_input[64]), .B(p_input[30064]), .Z(n7779) );
  AND U11671 ( .A(n7781), .B(n7782), .Z(o[649]) );
  AND U11672 ( .A(p_input[20649]), .B(p_input[10649]), .Z(n7782) );
  AND U11673 ( .A(p_input[649]), .B(p_input[30649]), .Z(n7781) );
  AND U11674 ( .A(n7783), .B(n7784), .Z(o[6499]) );
  AND U11675 ( .A(p_input[26499]), .B(p_input[16499]), .Z(n7784) );
  AND U11676 ( .A(p_input[6499]), .B(p_input[36499]), .Z(n7783) );
  AND U11677 ( .A(n7785), .B(n7786), .Z(o[6498]) );
  AND U11678 ( .A(p_input[26498]), .B(p_input[16498]), .Z(n7786) );
  AND U11679 ( .A(p_input[6498]), .B(p_input[36498]), .Z(n7785) );
  AND U11680 ( .A(n7787), .B(n7788), .Z(o[6497]) );
  AND U11681 ( .A(p_input[26497]), .B(p_input[16497]), .Z(n7788) );
  AND U11682 ( .A(p_input[6497]), .B(p_input[36497]), .Z(n7787) );
  AND U11683 ( .A(n7789), .B(n7790), .Z(o[6496]) );
  AND U11684 ( .A(p_input[26496]), .B(p_input[16496]), .Z(n7790) );
  AND U11685 ( .A(p_input[6496]), .B(p_input[36496]), .Z(n7789) );
  AND U11686 ( .A(n7791), .B(n7792), .Z(o[6495]) );
  AND U11687 ( .A(p_input[26495]), .B(p_input[16495]), .Z(n7792) );
  AND U11688 ( .A(p_input[6495]), .B(p_input[36495]), .Z(n7791) );
  AND U11689 ( .A(n7793), .B(n7794), .Z(o[6494]) );
  AND U11690 ( .A(p_input[26494]), .B(p_input[16494]), .Z(n7794) );
  AND U11691 ( .A(p_input[6494]), .B(p_input[36494]), .Z(n7793) );
  AND U11692 ( .A(n7795), .B(n7796), .Z(o[6493]) );
  AND U11693 ( .A(p_input[26493]), .B(p_input[16493]), .Z(n7796) );
  AND U11694 ( .A(p_input[6493]), .B(p_input[36493]), .Z(n7795) );
  AND U11695 ( .A(n7797), .B(n7798), .Z(o[6492]) );
  AND U11696 ( .A(p_input[26492]), .B(p_input[16492]), .Z(n7798) );
  AND U11697 ( .A(p_input[6492]), .B(p_input[36492]), .Z(n7797) );
  AND U11698 ( .A(n7799), .B(n7800), .Z(o[6491]) );
  AND U11699 ( .A(p_input[26491]), .B(p_input[16491]), .Z(n7800) );
  AND U11700 ( .A(p_input[6491]), .B(p_input[36491]), .Z(n7799) );
  AND U11701 ( .A(n7801), .B(n7802), .Z(o[6490]) );
  AND U11702 ( .A(p_input[26490]), .B(p_input[16490]), .Z(n7802) );
  AND U11703 ( .A(p_input[6490]), .B(p_input[36490]), .Z(n7801) );
  AND U11704 ( .A(n7803), .B(n7804), .Z(o[648]) );
  AND U11705 ( .A(p_input[20648]), .B(p_input[10648]), .Z(n7804) );
  AND U11706 ( .A(p_input[648]), .B(p_input[30648]), .Z(n7803) );
  AND U11707 ( .A(n7805), .B(n7806), .Z(o[6489]) );
  AND U11708 ( .A(p_input[26489]), .B(p_input[16489]), .Z(n7806) );
  AND U11709 ( .A(p_input[6489]), .B(p_input[36489]), .Z(n7805) );
  AND U11710 ( .A(n7807), .B(n7808), .Z(o[6488]) );
  AND U11711 ( .A(p_input[26488]), .B(p_input[16488]), .Z(n7808) );
  AND U11712 ( .A(p_input[6488]), .B(p_input[36488]), .Z(n7807) );
  AND U11713 ( .A(n7809), .B(n7810), .Z(o[6487]) );
  AND U11714 ( .A(p_input[26487]), .B(p_input[16487]), .Z(n7810) );
  AND U11715 ( .A(p_input[6487]), .B(p_input[36487]), .Z(n7809) );
  AND U11716 ( .A(n7811), .B(n7812), .Z(o[6486]) );
  AND U11717 ( .A(p_input[26486]), .B(p_input[16486]), .Z(n7812) );
  AND U11718 ( .A(p_input[6486]), .B(p_input[36486]), .Z(n7811) );
  AND U11719 ( .A(n7813), .B(n7814), .Z(o[6485]) );
  AND U11720 ( .A(p_input[26485]), .B(p_input[16485]), .Z(n7814) );
  AND U11721 ( .A(p_input[6485]), .B(p_input[36485]), .Z(n7813) );
  AND U11722 ( .A(n7815), .B(n7816), .Z(o[6484]) );
  AND U11723 ( .A(p_input[26484]), .B(p_input[16484]), .Z(n7816) );
  AND U11724 ( .A(p_input[6484]), .B(p_input[36484]), .Z(n7815) );
  AND U11725 ( .A(n7817), .B(n7818), .Z(o[6483]) );
  AND U11726 ( .A(p_input[26483]), .B(p_input[16483]), .Z(n7818) );
  AND U11727 ( .A(p_input[6483]), .B(p_input[36483]), .Z(n7817) );
  AND U11728 ( .A(n7819), .B(n7820), .Z(o[6482]) );
  AND U11729 ( .A(p_input[26482]), .B(p_input[16482]), .Z(n7820) );
  AND U11730 ( .A(p_input[6482]), .B(p_input[36482]), .Z(n7819) );
  AND U11731 ( .A(n7821), .B(n7822), .Z(o[6481]) );
  AND U11732 ( .A(p_input[26481]), .B(p_input[16481]), .Z(n7822) );
  AND U11733 ( .A(p_input[6481]), .B(p_input[36481]), .Z(n7821) );
  AND U11734 ( .A(n7823), .B(n7824), .Z(o[6480]) );
  AND U11735 ( .A(p_input[26480]), .B(p_input[16480]), .Z(n7824) );
  AND U11736 ( .A(p_input[6480]), .B(p_input[36480]), .Z(n7823) );
  AND U11737 ( .A(n7825), .B(n7826), .Z(o[647]) );
  AND U11738 ( .A(p_input[20647]), .B(p_input[10647]), .Z(n7826) );
  AND U11739 ( .A(p_input[647]), .B(p_input[30647]), .Z(n7825) );
  AND U11740 ( .A(n7827), .B(n7828), .Z(o[6479]) );
  AND U11741 ( .A(p_input[26479]), .B(p_input[16479]), .Z(n7828) );
  AND U11742 ( .A(p_input[6479]), .B(p_input[36479]), .Z(n7827) );
  AND U11743 ( .A(n7829), .B(n7830), .Z(o[6478]) );
  AND U11744 ( .A(p_input[26478]), .B(p_input[16478]), .Z(n7830) );
  AND U11745 ( .A(p_input[6478]), .B(p_input[36478]), .Z(n7829) );
  AND U11746 ( .A(n7831), .B(n7832), .Z(o[6477]) );
  AND U11747 ( .A(p_input[26477]), .B(p_input[16477]), .Z(n7832) );
  AND U11748 ( .A(p_input[6477]), .B(p_input[36477]), .Z(n7831) );
  AND U11749 ( .A(n7833), .B(n7834), .Z(o[6476]) );
  AND U11750 ( .A(p_input[26476]), .B(p_input[16476]), .Z(n7834) );
  AND U11751 ( .A(p_input[6476]), .B(p_input[36476]), .Z(n7833) );
  AND U11752 ( .A(n7835), .B(n7836), .Z(o[6475]) );
  AND U11753 ( .A(p_input[26475]), .B(p_input[16475]), .Z(n7836) );
  AND U11754 ( .A(p_input[6475]), .B(p_input[36475]), .Z(n7835) );
  AND U11755 ( .A(n7837), .B(n7838), .Z(o[6474]) );
  AND U11756 ( .A(p_input[26474]), .B(p_input[16474]), .Z(n7838) );
  AND U11757 ( .A(p_input[6474]), .B(p_input[36474]), .Z(n7837) );
  AND U11758 ( .A(n7839), .B(n7840), .Z(o[6473]) );
  AND U11759 ( .A(p_input[26473]), .B(p_input[16473]), .Z(n7840) );
  AND U11760 ( .A(p_input[6473]), .B(p_input[36473]), .Z(n7839) );
  AND U11761 ( .A(n7841), .B(n7842), .Z(o[6472]) );
  AND U11762 ( .A(p_input[26472]), .B(p_input[16472]), .Z(n7842) );
  AND U11763 ( .A(p_input[6472]), .B(p_input[36472]), .Z(n7841) );
  AND U11764 ( .A(n7843), .B(n7844), .Z(o[6471]) );
  AND U11765 ( .A(p_input[26471]), .B(p_input[16471]), .Z(n7844) );
  AND U11766 ( .A(p_input[6471]), .B(p_input[36471]), .Z(n7843) );
  AND U11767 ( .A(n7845), .B(n7846), .Z(o[6470]) );
  AND U11768 ( .A(p_input[26470]), .B(p_input[16470]), .Z(n7846) );
  AND U11769 ( .A(p_input[6470]), .B(p_input[36470]), .Z(n7845) );
  AND U11770 ( .A(n7847), .B(n7848), .Z(o[646]) );
  AND U11771 ( .A(p_input[20646]), .B(p_input[10646]), .Z(n7848) );
  AND U11772 ( .A(p_input[646]), .B(p_input[30646]), .Z(n7847) );
  AND U11773 ( .A(n7849), .B(n7850), .Z(o[6469]) );
  AND U11774 ( .A(p_input[26469]), .B(p_input[16469]), .Z(n7850) );
  AND U11775 ( .A(p_input[6469]), .B(p_input[36469]), .Z(n7849) );
  AND U11776 ( .A(n7851), .B(n7852), .Z(o[6468]) );
  AND U11777 ( .A(p_input[26468]), .B(p_input[16468]), .Z(n7852) );
  AND U11778 ( .A(p_input[6468]), .B(p_input[36468]), .Z(n7851) );
  AND U11779 ( .A(n7853), .B(n7854), .Z(o[6467]) );
  AND U11780 ( .A(p_input[26467]), .B(p_input[16467]), .Z(n7854) );
  AND U11781 ( .A(p_input[6467]), .B(p_input[36467]), .Z(n7853) );
  AND U11782 ( .A(n7855), .B(n7856), .Z(o[6466]) );
  AND U11783 ( .A(p_input[26466]), .B(p_input[16466]), .Z(n7856) );
  AND U11784 ( .A(p_input[6466]), .B(p_input[36466]), .Z(n7855) );
  AND U11785 ( .A(n7857), .B(n7858), .Z(o[6465]) );
  AND U11786 ( .A(p_input[26465]), .B(p_input[16465]), .Z(n7858) );
  AND U11787 ( .A(p_input[6465]), .B(p_input[36465]), .Z(n7857) );
  AND U11788 ( .A(n7859), .B(n7860), .Z(o[6464]) );
  AND U11789 ( .A(p_input[26464]), .B(p_input[16464]), .Z(n7860) );
  AND U11790 ( .A(p_input[6464]), .B(p_input[36464]), .Z(n7859) );
  AND U11791 ( .A(n7861), .B(n7862), .Z(o[6463]) );
  AND U11792 ( .A(p_input[26463]), .B(p_input[16463]), .Z(n7862) );
  AND U11793 ( .A(p_input[6463]), .B(p_input[36463]), .Z(n7861) );
  AND U11794 ( .A(n7863), .B(n7864), .Z(o[6462]) );
  AND U11795 ( .A(p_input[26462]), .B(p_input[16462]), .Z(n7864) );
  AND U11796 ( .A(p_input[6462]), .B(p_input[36462]), .Z(n7863) );
  AND U11797 ( .A(n7865), .B(n7866), .Z(o[6461]) );
  AND U11798 ( .A(p_input[26461]), .B(p_input[16461]), .Z(n7866) );
  AND U11799 ( .A(p_input[6461]), .B(p_input[36461]), .Z(n7865) );
  AND U11800 ( .A(n7867), .B(n7868), .Z(o[6460]) );
  AND U11801 ( .A(p_input[26460]), .B(p_input[16460]), .Z(n7868) );
  AND U11802 ( .A(p_input[6460]), .B(p_input[36460]), .Z(n7867) );
  AND U11803 ( .A(n7869), .B(n7870), .Z(o[645]) );
  AND U11804 ( .A(p_input[20645]), .B(p_input[10645]), .Z(n7870) );
  AND U11805 ( .A(p_input[645]), .B(p_input[30645]), .Z(n7869) );
  AND U11806 ( .A(n7871), .B(n7872), .Z(o[6459]) );
  AND U11807 ( .A(p_input[26459]), .B(p_input[16459]), .Z(n7872) );
  AND U11808 ( .A(p_input[6459]), .B(p_input[36459]), .Z(n7871) );
  AND U11809 ( .A(n7873), .B(n7874), .Z(o[6458]) );
  AND U11810 ( .A(p_input[26458]), .B(p_input[16458]), .Z(n7874) );
  AND U11811 ( .A(p_input[6458]), .B(p_input[36458]), .Z(n7873) );
  AND U11812 ( .A(n7875), .B(n7876), .Z(o[6457]) );
  AND U11813 ( .A(p_input[26457]), .B(p_input[16457]), .Z(n7876) );
  AND U11814 ( .A(p_input[6457]), .B(p_input[36457]), .Z(n7875) );
  AND U11815 ( .A(n7877), .B(n7878), .Z(o[6456]) );
  AND U11816 ( .A(p_input[26456]), .B(p_input[16456]), .Z(n7878) );
  AND U11817 ( .A(p_input[6456]), .B(p_input[36456]), .Z(n7877) );
  AND U11818 ( .A(n7879), .B(n7880), .Z(o[6455]) );
  AND U11819 ( .A(p_input[26455]), .B(p_input[16455]), .Z(n7880) );
  AND U11820 ( .A(p_input[6455]), .B(p_input[36455]), .Z(n7879) );
  AND U11821 ( .A(n7881), .B(n7882), .Z(o[6454]) );
  AND U11822 ( .A(p_input[26454]), .B(p_input[16454]), .Z(n7882) );
  AND U11823 ( .A(p_input[6454]), .B(p_input[36454]), .Z(n7881) );
  AND U11824 ( .A(n7883), .B(n7884), .Z(o[6453]) );
  AND U11825 ( .A(p_input[26453]), .B(p_input[16453]), .Z(n7884) );
  AND U11826 ( .A(p_input[6453]), .B(p_input[36453]), .Z(n7883) );
  AND U11827 ( .A(n7885), .B(n7886), .Z(o[6452]) );
  AND U11828 ( .A(p_input[26452]), .B(p_input[16452]), .Z(n7886) );
  AND U11829 ( .A(p_input[6452]), .B(p_input[36452]), .Z(n7885) );
  AND U11830 ( .A(n7887), .B(n7888), .Z(o[6451]) );
  AND U11831 ( .A(p_input[26451]), .B(p_input[16451]), .Z(n7888) );
  AND U11832 ( .A(p_input[6451]), .B(p_input[36451]), .Z(n7887) );
  AND U11833 ( .A(n7889), .B(n7890), .Z(o[6450]) );
  AND U11834 ( .A(p_input[26450]), .B(p_input[16450]), .Z(n7890) );
  AND U11835 ( .A(p_input[6450]), .B(p_input[36450]), .Z(n7889) );
  AND U11836 ( .A(n7891), .B(n7892), .Z(o[644]) );
  AND U11837 ( .A(p_input[20644]), .B(p_input[10644]), .Z(n7892) );
  AND U11838 ( .A(p_input[644]), .B(p_input[30644]), .Z(n7891) );
  AND U11839 ( .A(n7893), .B(n7894), .Z(o[6449]) );
  AND U11840 ( .A(p_input[26449]), .B(p_input[16449]), .Z(n7894) );
  AND U11841 ( .A(p_input[6449]), .B(p_input[36449]), .Z(n7893) );
  AND U11842 ( .A(n7895), .B(n7896), .Z(o[6448]) );
  AND U11843 ( .A(p_input[26448]), .B(p_input[16448]), .Z(n7896) );
  AND U11844 ( .A(p_input[6448]), .B(p_input[36448]), .Z(n7895) );
  AND U11845 ( .A(n7897), .B(n7898), .Z(o[6447]) );
  AND U11846 ( .A(p_input[26447]), .B(p_input[16447]), .Z(n7898) );
  AND U11847 ( .A(p_input[6447]), .B(p_input[36447]), .Z(n7897) );
  AND U11848 ( .A(n7899), .B(n7900), .Z(o[6446]) );
  AND U11849 ( .A(p_input[26446]), .B(p_input[16446]), .Z(n7900) );
  AND U11850 ( .A(p_input[6446]), .B(p_input[36446]), .Z(n7899) );
  AND U11851 ( .A(n7901), .B(n7902), .Z(o[6445]) );
  AND U11852 ( .A(p_input[26445]), .B(p_input[16445]), .Z(n7902) );
  AND U11853 ( .A(p_input[6445]), .B(p_input[36445]), .Z(n7901) );
  AND U11854 ( .A(n7903), .B(n7904), .Z(o[6444]) );
  AND U11855 ( .A(p_input[26444]), .B(p_input[16444]), .Z(n7904) );
  AND U11856 ( .A(p_input[6444]), .B(p_input[36444]), .Z(n7903) );
  AND U11857 ( .A(n7905), .B(n7906), .Z(o[6443]) );
  AND U11858 ( .A(p_input[26443]), .B(p_input[16443]), .Z(n7906) );
  AND U11859 ( .A(p_input[6443]), .B(p_input[36443]), .Z(n7905) );
  AND U11860 ( .A(n7907), .B(n7908), .Z(o[6442]) );
  AND U11861 ( .A(p_input[26442]), .B(p_input[16442]), .Z(n7908) );
  AND U11862 ( .A(p_input[6442]), .B(p_input[36442]), .Z(n7907) );
  AND U11863 ( .A(n7909), .B(n7910), .Z(o[6441]) );
  AND U11864 ( .A(p_input[26441]), .B(p_input[16441]), .Z(n7910) );
  AND U11865 ( .A(p_input[6441]), .B(p_input[36441]), .Z(n7909) );
  AND U11866 ( .A(n7911), .B(n7912), .Z(o[6440]) );
  AND U11867 ( .A(p_input[26440]), .B(p_input[16440]), .Z(n7912) );
  AND U11868 ( .A(p_input[6440]), .B(p_input[36440]), .Z(n7911) );
  AND U11869 ( .A(n7913), .B(n7914), .Z(o[643]) );
  AND U11870 ( .A(p_input[20643]), .B(p_input[10643]), .Z(n7914) );
  AND U11871 ( .A(p_input[643]), .B(p_input[30643]), .Z(n7913) );
  AND U11872 ( .A(n7915), .B(n7916), .Z(o[6439]) );
  AND U11873 ( .A(p_input[26439]), .B(p_input[16439]), .Z(n7916) );
  AND U11874 ( .A(p_input[6439]), .B(p_input[36439]), .Z(n7915) );
  AND U11875 ( .A(n7917), .B(n7918), .Z(o[6438]) );
  AND U11876 ( .A(p_input[26438]), .B(p_input[16438]), .Z(n7918) );
  AND U11877 ( .A(p_input[6438]), .B(p_input[36438]), .Z(n7917) );
  AND U11878 ( .A(n7919), .B(n7920), .Z(o[6437]) );
  AND U11879 ( .A(p_input[26437]), .B(p_input[16437]), .Z(n7920) );
  AND U11880 ( .A(p_input[6437]), .B(p_input[36437]), .Z(n7919) );
  AND U11881 ( .A(n7921), .B(n7922), .Z(o[6436]) );
  AND U11882 ( .A(p_input[26436]), .B(p_input[16436]), .Z(n7922) );
  AND U11883 ( .A(p_input[6436]), .B(p_input[36436]), .Z(n7921) );
  AND U11884 ( .A(n7923), .B(n7924), .Z(o[6435]) );
  AND U11885 ( .A(p_input[26435]), .B(p_input[16435]), .Z(n7924) );
  AND U11886 ( .A(p_input[6435]), .B(p_input[36435]), .Z(n7923) );
  AND U11887 ( .A(n7925), .B(n7926), .Z(o[6434]) );
  AND U11888 ( .A(p_input[26434]), .B(p_input[16434]), .Z(n7926) );
  AND U11889 ( .A(p_input[6434]), .B(p_input[36434]), .Z(n7925) );
  AND U11890 ( .A(n7927), .B(n7928), .Z(o[6433]) );
  AND U11891 ( .A(p_input[26433]), .B(p_input[16433]), .Z(n7928) );
  AND U11892 ( .A(p_input[6433]), .B(p_input[36433]), .Z(n7927) );
  AND U11893 ( .A(n7929), .B(n7930), .Z(o[6432]) );
  AND U11894 ( .A(p_input[26432]), .B(p_input[16432]), .Z(n7930) );
  AND U11895 ( .A(p_input[6432]), .B(p_input[36432]), .Z(n7929) );
  AND U11896 ( .A(n7931), .B(n7932), .Z(o[6431]) );
  AND U11897 ( .A(p_input[26431]), .B(p_input[16431]), .Z(n7932) );
  AND U11898 ( .A(p_input[6431]), .B(p_input[36431]), .Z(n7931) );
  AND U11899 ( .A(n7933), .B(n7934), .Z(o[6430]) );
  AND U11900 ( .A(p_input[26430]), .B(p_input[16430]), .Z(n7934) );
  AND U11901 ( .A(p_input[6430]), .B(p_input[36430]), .Z(n7933) );
  AND U11902 ( .A(n7935), .B(n7936), .Z(o[642]) );
  AND U11903 ( .A(p_input[20642]), .B(p_input[10642]), .Z(n7936) );
  AND U11904 ( .A(p_input[642]), .B(p_input[30642]), .Z(n7935) );
  AND U11905 ( .A(n7937), .B(n7938), .Z(o[6429]) );
  AND U11906 ( .A(p_input[26429]), .B(p_input[16429]), .Z(n7938) );
  AND U11907 ( .A(p_input[6429]), .B(p_input[36429]), .Z(n7937) );
  AND U11908 ( .A(n7939), .B(n7940), .Z(o[6428]) );
  AND U11909 ( .A(p_input[26428]), .B(p_input[16428]), .Z(n7940) );
  AND U11910 ( .A(p_input[6428]), .B(p_input[36428]), .Z(n7939) );
  AND U11911 ( .A(n7941), .B(n7942), .Z(o[6427]) );
  AND U11912 ( .A(p_input[26427]), .B(p_input[16427]), .Z(n7942) );
  AND U11913 ( .A(p_input[6427]), .B(p_input[36427]), .Z(n7941) );
  AND U11914 ( .A(n7943), .B(n7944), .Z(o[6426]) );
  AND U11915 ( .A(p_input[26426]), .B(p_input[16426]), .Z(n7944) );
  AND U11916 ( .A(p_input[6426]), .B(p_input[36426]), .Z(n7943) );
  AND U11917 ( .A(n7945), .B(n7946), .Z(o[6425]) );
  AND U11918 ( .A(p_input[26425]), .B(p_input[16425]), .Z(n7946) );
  AND U11919 ( .A(p_input[6425]), .B(p_input[36425]), .Z(n7945) );
  AND U11920 ( .A(n7947), .B(n7948), .Z(o[6424]) );
  AND U11921 ( .A(p_input[26424]), .B(p_input[16424]), .Z(n7948) );
  AND U11922 ( .A(p_input[6424]), .B(p_input[36424]), .Z(n7947) );
  AND U11923 ( .A(n7949), .B(n7950), .Z(o[6423]) );
  AND U11924 ( .A(p_input[26423]), .B(p_input[16423]), .Z(n7950) );
  AND U11925 ( .A(p_input[6423]), .B(p_input[36423]), .Z(n7949) );
  AND U11926 ( .A(n7951), .B(n7952), .Z(o[6422]) );
  AND U11927 ( .A(p_input[26422]), .B(p_input[16422]), .Z(n7952) );
  AND U11928 ( .A(p_input[6422]), .B(p_input[36422]), .Z(n7951) );
  AND U11929 ( .A(n7953), .B(n7954), .Z(o[6421]) );
  AND U11930 ( .A(p_input[26421]), .B(p_input[16421]), .Z(n7954) );
  AND U11931 ( .A(p_input[6421]), .B(p_input[36421]), .Z(n7953) );
  AND U11932 ( .A(n7955), .B(n7956), .Z(o[6420]) );
  AND U11933 ( .A(p_input[26420]), .B(p_input[16420]), .Z(n7956) );
  AND U11934 ( .A(p_input[6420]), .B(p_input[36420]), .Z(n7955) );
  AND U11935 ( .A(n7957), .B(n7958), .Z(o[641]) );
  AND U11936 ( .A(p_input[20641]), .B(p_input[10641]), .Z(n7958) );
  AND U11937 ( .A(p_input[641]), .B(p_input[30641]), .Z(n7957) );
  AND U11938 ( .A(n7959), .B(n7960), .Z(o[6419]) );
  AND U11939 ( .A(p_input[26419]), .B(p_input[16419]), .Z(n7960) );
  AND U11940 ( .A(p_input[6419]), .B(p_input[36419]), .Z(n7959) );
  AND U11941 ( .A(n7961), .B(n7962), .Z(o[6418]) );
  AND U11942 ( .A(p_input[26418]), .B(p_input[16418]), .Z(n7962) );
  AND U11943 ( .A(p_input[6418]), .B(p_input[36418]), .Z(n7961) );
  AND U11944 ( .A(n7963), .B(n7964), .Z(o[6417]) );
  AND U11945 ( .A(p_input[26417]), .B(p_input[16417]), .Z(n7964) );
  AND U11946 ( .A(p_input[6417]), .B(p_input[36417]), .Z(n7963) );
  AND U11947 ( .A(n7965), .B(n7966), .Z(o[6416]) );
  AND U11948 ( .A(p_input[26416]), .B(p_input[16416]), .Z(n7966) );
  AND U11949 ( .A(p_input[6416]), .B(p_input[36416]), .Z(n7965) );
  AND U11950 ( .A(n7967), .B(n7968), .Z(o[6415]) );
  AND U11951 ( .A(p_input[26415]), .B(p_input[16415]), .Z(n7968) );
  AND U11952 ( .A(p_input[6415]), .B(p_input[36415]), .Z(n7967) );
  AND U11953 ( .A(n7969), .B(n7970), .Z(o[6414]) );
  AND U11954 ( .A(p_input[26414]), .B(p_input[16414]), .Z(n7970) );
  AND U11955 ( .A(p_input[6414]), .B(p_input[36414]), .Z(n7969) );
  AND U11956 ( .A(n7971), .B(n7972), .Z(o[6413]) );
  AND U11957 ( .A(p_input[26413]), .B(p_input[16413]), .Z(n7972) );
  AND U11958 ( .A(p_input[6413]), .B(p_input[36413]), .Z(n7971) );
  AND U11959 ( .A(n7973), .B(n7974), .Z(o[6412]) );
  AND U11960 ( .A(p_input[26412]), .B(p_input[16412]), .Z(n7974) );
  AND U11961 ( .A(p_input[6412]), .B(p_input[36412]), .Z(n7973) );
  AND U11962 ( .A(n7975), .B(n7976), .Z(o[6411]) );
  AND U11963 ( .A(p_input[26411]), .B(p_input[16411]), .Z(n7976) );
  AND U11964 ( .A(p_input[6411]), .B(p_input[36411]), .Z(n7975) );
  AND U11965 ( .A(n7977), .B(n7978), .Z(o[6410]) );
  AND U11966 ( .A(p_input[26410]), .B(p_input[16410]), .Z(n7978) );
  AND U11967 ( .A(p_input[6410]), .B(p_input[36410]), .Z(n7977) );
  AND U11968 ( .A(n7979), .B(n7980), .Z(o[640]) );
  AND U11969 ( .A(p_input[20640]), .B(p_input[10640]), .Z(n7980) );
  AND U11970 ( .A(p_input[640]), .B(p_input[30640]), .Z(n7979) );
  AND U11971 ( .A(n7981), .B(n7982), .Z(o[6409]) );
  AND U11972 ( .A(p_input[26409]), .B(p_input[16409]), .Z(n7982) );
  AND U11973 ( .A(p_input[6409]), .B(p_input[36409]), .Z(n7981) );
  AND U11974 ( .A(n7983), .B(n7984), .Z(o[6408]) );
  AND U11975 ( .A(p_input[26408]), .B(p_input[16408]), .Z(n7984) );
  AND U11976 ( .A(p_input[6408]), .B(p_input[36408]), .Z(n7983) );
  AND U11977 ( .A(n7985), .B(n7986), .Z(o[6407]) );
  AND U11978 ( .A(p_input[26407]), .B(p_input[16407]), .Z(n7986) );
  AND U11979 ( .A(p_input[6407]), .B(p_input[36407]), .Z(n7985) );
  AND U11980 ( .A(n7987), .B(n7988), .Z(o[6406]) );
  AND U11981 ( .A(p_input[26406]), .B(p_input[16406]), .Z(n7988) );
  AND U11982 ( .A(p_input[6406]), .B(p_input[36406]), .Z(n7987) );
  AND U11983 ( .A(n7989), .B(n7990), .Z(o[6405]) );
  AND U11984 ( .A(p_input[26405]), .B(p_input[16405]), .Z(n7990) );
  AND U11985 ( .A(p_input[6405]), .B(p_input[36405]), .Z(n7989) );
  AND U11986 ( .A(n7991), .B(n7992), .Z(o[6404]) );
  AND U11987 ( .A(p_input[26404]), .B(p_input[16404]), .Z(n7992) );
  AND U11988 ( .A(p_input[6404]), .B(p_input[36404]), .Z(n7991) );
  AND U11989 ( .A(n7993), .B(n7994), .Z(o[6403]) );
  AND U11990 ( .A(p_input[26403]), .B(p_input[16403]), .Z(n7994) );
  AND U11991 ( .A(p_input[6403]), .B(p_input[36403]), .Z(n7993) );
  AND U11992 ( .A(n7995), .B(n7996), .Z(o[6402]) );
  AND U11993 ( .A(p_input[26402]), .B(p_input[16402]), .Z(n7996) );
  AND U11994 ( .A(p_input[6402]), .B(p_input[36402]), .Z(n7995) );
  AND U11995 ( .A(n7997), .B(n7998), .Z(o[6401]) );
  AND U11996 ( .A(p_input[26401]), .B(p_input[16401]), .Z(n7998) );
  AND U11997 ( .A(p_input[6401]), .B(p_input[36401]), .Z(n7997) );
  AND U11998 ( .A(n7999), .B(n8000), .Z(o[6400]) );
  AND U11999 ( .A(p_input[26400]), .B(p_input[16400]), .Z(n8000) );
  AND U12000 ( .A(p_input[6400]), .B(p_input[36400]), .Z(n7999) );
  AND U12001 ( .A(n8001), .B(n8002), .Z(o[63]) );
  AND U12002 ( .A(p_input[20063]), .B(p_input[10063]), .Z(n8002) );
  AND U12003 ( .A(p_input[63]), .B(p_input[30063]), .Z(n8001) );
  AND U12004 ( .A(n8003), .B(n8004), .Z(o[639]) );
  AND U12005 ( .A(p_input[20639]), .B(p_input[10639]), .Z(n8004) );
  AND U12006 ( .A(p_input[639]), .B(p_input[30639]), .Z(n8003) );
  AND U12007 ( .A(n8005), .B(n8006), .Z(o[6399]) );
  AND U12008 ( .A(p_input[26399]), .B(p_input[16399]), .Z(n8006) );
  AND U12009 ( .A(p_input[6399]), .B(p_input[36399]), .Z(n8005) );
  AND U12010 ( .A(n8007), .B(n8008), .Z(o[6398]) );
  AND U12011 ( .A(p_input[26398]), .B(p_input[16398]), .Z(n8008) );
  AND U12012 ( .A(p_input[6398]), .B(p_input[36398]), .Z(n8007) );
  AND U12013 ( .A(n8009), .B(n8010), .Z(o[6397]) );
  AND U12014 ( .A(p_input[26397]), .B(p_input[16397]), .Z(n8010) );
  AND U12015 ( .A(p_input[6397]), .B(p_input[36397]), .Z(n8009) );
  AND U12016 ( .A(n8011), .B(n8012), .Z(o[6396]) );
  AND U12017 ( .A(p_input[26396]), .B(p_input[16396]), .Z(n8012) );
  AND U12018 ( .A(p_input[6396]), .B(p_input[36396]), .Z(n8011) );
  AND U12019 ( .A(n8013), .B(n8014), .Z(o[6395]) );
  AND U12020 ( .A(p_input[26395]), .B(p_input[16395]), .Z(n8014) );
  AND U12021 ( .A(p_input[6395]), .B(p_input[36395]), .Z(n8013) );
  AND U12022 ( .A(n8015), .B(n8016), .Z(o[6394]) );
  AND U12023 ( .A(p_input[26394]), .B(p_input[16394]), .Z(n8016) );
  AND U12024 ( .A(p_input[6394]), .B(p_input[36394]), .Z(n8015) );
  AND U12025 ( .A(n8017), .B(n8018), .Z(o[6393]) );
  AND U12026 ( .A(p_input[26393]), .B(p_input[16393]), .Z(n8018) );
  AND U12027 ( .A(p_input[6393]), .B(p_input[36393]), .Z(n8017) );
  AND U12028 ( .A(n8019), .B(n8020), .Z(o[6392]) );
  AND U12029 ( .A(p_input[26392]), .B(p_input[16392]), .Z(n8020) );
  AND U12030 ( .A(p_input[6392]), .B(p_input[36392]), .Z(n8019) );
  AND U12031 ( .A(n8021), .B(n8022), .Z(o[6391]) );
  AND U12032 ( .A(p_input[26391]), .B(p_input[16391]), .Z(n8022) );
  AND U12033 ( .A(p_input[6391]), .B(p_input[36391]), .Z(n8021) );
  AND U12034 ( .A(n8023), .B(n8024), .Z(o[6390]) );
  AND U12035 ( .A(p_input[26390]), .B(p_input[16390]), .Z(n8024) );
  AND U12036 ( .A(p_input[6390]), .B(p_input[36390]), .Z(n8023) );
  AND U12037 ( .A(n8025), .B(n8026), .Z(o[638]) );
  AND U12038 ( .A(p_input[20638]), .B(p_input[10638]), .Z(n8026) );
  AND U12039 ( .A(p_input[638]), .B(p_input[30638]), .Z(n8025) );
  AND U12040 ( .A(n8027), .B(n8028), .Z(o[6389]) );
  AND U12041 ( .A(p_input[26389]), .B(p_input[16389]), .Z(n8028) );
  AND U12042 ( .A(p_input[6389]), .B(p_input[36389]), .Z(n8027) );
  AND U12043 ( .A(n8029), .B(n8030), .Z(o[6388]) );
  AND U12044 ( .A(p_input[26388]), .B(p_input[16388]), .Z(n8030) );
  AND U12045 ( .A(p_input[6388]), .B(p_input[36388]), .Z(n8029) );
  AND U12046 ( .A(n8031), .B(n8032), .Z(o[6387]) );
  AND U12047 ( .A(p_input[26387]), .B(p_input[16387]), .Z(n8032) );
  AND U12048 ( .A(p_input[6387]), .B(p_input[36387]), .Z(n8031) );
  AND U12049 ( .A(n8033), .B(n8034), .Z(o[6386]) );
  AND U12050 ( .A(p_input[26386]), .B(p_input[16386]), .Z(n8034) );
  AND U12051 ( .A(p_input[6386]), .B(p_input[36386]), .Z(n8033) );
  AND U12052 ( .A(n8035), .B(n8036), .Z(o[6385]) );
  AND U12053 ( .A(p_input[26385]), .B(p_input[16385]), .Z(n8036) );
  AND U12054 ( .A(p_input[6385]), .B(p_input[36385]), .Z(n8035) );
  AND U12055 ( .A(n8037), .B(n8038), .Z(o[6384]) );
  AND U12056 ( .A(p_input[26384]), .B(p_input[16384]), .Z(n8038) );
  AND U12057 ( .A(p_input[6384]), .B(p_input[36384]), .Z(n8037) );
  AND U12058 ( .A(n8039), .B(n8040), .Z(o[6383]) );
  AND U12059 ( .A(p_input[26383]), .B(p_input[16383]), .Z(n8040) );
  AND U12060 ( .A(p_input[6383]), .B(p_input[36383]), .Z(n8039) );
  AND U12061 ( .A(n8041), .B(n8042), .Z(o[6382]) );
  AND U12062 ( .A(p_input[26382]), .B(p_input[16382]), .Z(n8042) );
  AND U12063 ( .A(p_input[6382]), .B(p_input[36382]), .Z(n8041) );
  AND U12064 ( .A(n8043), .B(n8044), .Z(o[6381]) );
  AND U12065 ( .A(p_input[26381]), .B(p_input[16381]), .Z(n8044) );
  AND U12066 ( .A(p_input[6381]), .B(p_input[36381]), .Z(n8043) );
  AND U12067 ( .A(n8045), .B(n8046), .Z(o[6380]) );
  AND U12068 ( .A(p_input[26380]), .B(p_input[16380]), .Z(n8046) );
  AND U12069 ( .A(p_input[6380]), .B(p_input[36380]), .Z(n8045) );
  AND U12070 ( .A(n8047), .B(n8048), .Z(o[637]) );
  AND U12071 ( .A(p_input[20637]), .B(p_input[10637]), .Z(n8048) );
  AND U12072 ( .A(p_input[637]), .B(p_input[30637]), .Z(n8047) );
  AND U12073 ( .A(n8049), .B(n8050), .Z(o[6379]) );
  AND U12074 ( .A(p_input[26379]), .B(p_input[16379]), .Z(n8050) );
  AND U12075 ( .A(p_input[6379]), .B(p_input[36379]), .Z(n8049) );
  AND U12076 ( .A(n8051), .B(n8052), .Z(o[6378]) );
  AND U12077 ( .A(p_input[26378]), .B(p_input[16378]), .Z(n8052) );
  AND U12078 ( .A(p_input[6378]), .B(p_input[36378]), .Z(n8051) );
  AND U12079 ( .A(n8053), .B(n8054), .Z(o[6377]) );
  AND U12080 ( .A(p_input[26377]), .B(p_input[16377]), .Z(n8054) );
  AND U12081 ( .A(p_input[6377]), .B(p_input[36377]), .Z(n8053) );
  AND U12082 ( .A(n8055), .B(n8056), .Z(o[6376]) );
  AND U12083 ( .A(p_input[26376]), .B(p_input[16376]), .Z(n8056) );
  AND U12084 ( .A(p_input[6376]), .B(p_input[36376]), .Z(n8055) );
  AND U12085 ( .A(n8057), .B(n8058), .Z(o[6375]) );
  AND U12086 ( .A(p_input[26375]), .B(p_input[16375]), .Z(n8058) );
  AND U12087 ( .A(p_input[6375]), .B(p_input[36375]), .Z(n8057) );
  AND U12088 ( .A(n8059), .B(n8060), .Z(o[6374]) );
  AND U12089 ( .A(p_input[26374]), .B(p_input[16374]), .Z(n8060) );
  AND U12090 ( .A(p_input[6374]), .B(p_input[36374]), .Z(n8059) );
  AND U12091 ( .A(n8061), .B(n8062), .Z(o[6373]) );
  AND U12092 ( .A(p_input[26373]), .B(p_input[16373]), .Z(n8062) );
  AND U12093 ( .A(p_input[6373]), .B(p_input[36373]), .Z(n8061) );
  AND U12094 ( .A(n8063), .B(n8064), .Z(o[6372]) );
  AND U12095 ( .A(p_input[26372]), .B(p_input[16372]), .Z(n8064) );
  AND U12096 ( .A(p_input[6372]), .B(p_input[36372]), .Z(n8063) );
  AND U12097 ( .A(n8065), .B(n8066), .Z(o[6371]) );
  AND U12098 ( .A(p_input[26371]), .B(p_input[16371]), .Z(n8066) );
  AND U12099 ( .A(p_input[6371]), .B(p_input[36371]), .Z(n8065) );
  AND U12100 ( .A(n8067), .B(n8068), .Z(o[6370]) );
  AND U12101 ( .A(p_input[26370]), .B(p_input[16370]), .Z(n8068) );
  AND U12102 ( .A(p_input[6370]), .B(p_input[36370]), .Z(n8067) );
  AND U12103 ( .A(n8069), .B(n8070), .Z(o[636]) );
  AND U12104 ( .A(p_input[20636]), .B(p_input[10636]), .Z(n8070) );
  AND U12105 ( .A(p_input[636]), .B(p_input[30636]), .Z(n8069) );
  AND U12106 ( .A(n8071), .B(n8072), .Z(o[6369]) );
  AND U12107 ( .A(p_input[26369]), .B(p_input[16369]), .Z(n8072) );
  AND U12108 ( .A(p_input[6369]), .B(p_input[36369]), .Z(n8071) );
  AND U12109 ( .A(n8073), .B(n8074), .Z(o[6368]) );
  AND U12110 ( .A(p_input[26368]), .B(p_input[16368]), .Z(n8074) );
  AND U12111 ( .A(p_input[6368]), .B(p_input[36368]), .Z(n8073) );
  AND U12112 ( .A(n8075), .B(n8076), .Z(o[6367]) );
  AND U12113 ( .A(p_input[26367]), .B(p_input[16367]), .Z(n8076) );
  AND U12114 ( .A(p_input[6367]), .B(p_input[36367]), .Z(n8075) );
  AND U12115 ( .A(n8077), .B(n8078), .Z(o[6366]) );
  AND U12116 ( .A(p_input[26366]), .B(p_input[16366]), .Z(n8078) );
  AND U12117 ( .A(p_input[6366]), .B(p_input[36366]), .Z(n8077) );
  AND U12118 ( .A(n8079), .B(n8080), .Z(o[6365]) );
  AND U12119 ( .A(p_input[26365]), .B(p_input[16365]), .Z(n8080) );
  AND U12120 ( .A(p_input[6365]), .B(p_input[36365]), .Z(n8079) );
  AND U12121 ( .A(n8081), .B(n8082), .Z(o[6364]) );
  AND U12122 ( .A(p_input[26364]), .B(p_input[16364]), .Z(n8082) );
  AND U12123 ( .A(p_input[6364]), .B(p_input[36364]), .Z(n8081) );
  AND U12124 ( .A(n8083), .B(n8084), .Z(o[6363]) );
  AND U12125 ( .A(p_input[26363]), .B(p_input[16363]), .Z(n8084) );
  AND U12126 ( .A(p_input[6363]), .B(p_input[36363]), .Z(n8083) );
  AND U12127 ( .A(n8085), .B(n8086), .Z(o[6362]) );
  AND U12128 ( .A(p_input[26362]), .B(p_input[16362]), .Z(n8086) );
  AND U12129 ( .A(p_input[6362]), .B(p_input[36362]), .Z(n8085) );
  AND U12130 ( .A(n8087), .B(n8088), .Z(o[6361]) );
  AND U12131 ( .A(p_input[26361]), .B(p_input[16361]), .Z(n8088) );
  AND U12132 ( .A(p_input[6361]), .B(p_input[36361]), .Z(n8087) );
  AND U12133 ( .A(n8089), .B(n8090), .Z(o[6360]) );
  AND U12134 ( .A(p_input[26360]), .B(p_input[16360]), .Z(n8090) );
  AND U12135 ( .A(p_input[6360]), .B(p_input[36360]), .Z(n8089) );
  AND U12136 ( .A(n8091), .B(n8092), .Z(o[635]) );
  AND U12137 ( .A(p_input[20635]), .B(p_input[10635]), .Z(n8092) );
  AND U12138 ( .A(p_input[635]), .B(p_input[30635]), .Z(n8091) );
  AND U12139 ( .A(n8093), .B(n8094), .Z(o[6359]) );
  AND U12140 ( .A(p_input[26359]), .B(p_input[16359]), .Z(n8094) );
  AND U12141 ( .A(p_input[6359]), .B(p_input[36359]), .Z(n8093) );
  AND U12142 ( .A(n8095), .B(n8096), .Z(o[6358]) );
  AND U12143 ( .A(p_input[26358]), .B(p_input[16358]), .Z(n8096) );
  AND U12144 ( .A(p_input[6358]), .B(p_input[36358]), .Z(n8095) );
  AND U12145 ( .A(n8097), .B(n8098), .Z(o[6357]) );
  AND U12146 ( .A(p_input[26357]), .B(p_input[16357]), .Z(n8098) );
  AND U12147 ( .A(p_input[6357]), .B(p_input[36357]), .Z(n8097) );
  AND U12148 ( .A(n8099), .B(n8100), .Z(o[6356]) );
  AND U12149 ( .A(p_input[26356]), .B(p_input[16356]), .Z(n8100) );
  AND U12150 ( .A(p_input[6356]), .B(p_input[36356]), .Z(n8099) );
  AND U12151 ( .A(n8101), .B(n8102), .Z(o[6355]) );
  AND U12152 ( .A(p_input[26355]), .B(p_input[16355]), .Z(n8102) );
  AND U12153 ( .A(p_input[6355]), .B(p_input[36355]), .Z(n8101) );
  AND U12154 ( .A(n8103), .B(n8104), .Z(o[6354]) );
  AND U12155 ( .A(p_input[26354]), .B(p_input[16354]), .Z(n8104) );
  AND U12156 ( .A(p_input[6354]), .B(p_input[36354]), .Z(n8103) );
  AND U12157 ( .A(n8105), .B(n8106), .Z(o[6353]) );
  AND U12158 ( .A(p_input[26353]), .B(p_input[16353]), .Z(n8106) );
  AND U12159 ( .A(p_input[6353]), .B(p_input[36353]), .Z(n8105) );
  AND U12160 ( .A(n8107), .B(n8108), .Z(o[6352]) );
  AND U12161 ( .A(p_input[26352]), .B(p_input[16352]), .Z(n8108) );
  AND U12162 ( .A(p_input[6352]), .B(p_input[36352]), .Z(n8107) );
  AND U12163 ( .A(n8109), .B(n8110), .Z(o[6351]) );
  AND U12164 ( .A(p_input[26351]), .B(p_input[16351]), .Z(n8110) );
  AND U12165 ( .A(p_input[6351]), .B(p_input[36351]), .Z(n8109) );
  AND U12166 ( .A(n8111), .B(n8112), .Z(o[6350]) );
  AND U12167 ( .A(p_input[26350]), .B(p_input[16350]), .Z(n8112) );
  AND U12168 ( .A(p_input[6350]), .B(p_input[36350]), .Z(n8111) );
  AND U12169 ( .A(n8113), .B(n8114), .Z(o[634]) );
  AND U12170 ( .A(p_input[20634]), .B(p_input[10634]), .Z(n8114) );
  AND U12171 ( .A(p_input[634]), .B(p_input[30634]), .Z(n8113) );
  AND U12172 ( .A(n8115), .B(n8116), .Z(o[6349]) );
  AND U12173 ( .A(p_input[26349]), .B(p_input[16349]), .Z(n8116) );
  AND U12174 ( .A(p_input[6349]), .B(p_input[36349]), .Z(n8115) );
  AND U12175 ( .A(n8117), .B(n8118), .Z(o[6348]) );
  AND U12176 ( .A(p_input[26348]), .B(p_input[16348]), .Z(n8118) );
  AND U12177 ( .A(p_input[6348]), .B(p_input[36348]), .Z(n8117) );
  AND U12178 ( .A(n8119), .B(n8120), .Z(o[6347]) );
  AND U12179 ( .A(p_input[26347]), .B(p_input[16347]), .Z(n8120) );
  AND U12180 ( .A(p_input[6347]), .B(p_input[36347]), .Z(n8119) );
  AND U12181 ( .A(n8121), .B(n8122), .Z(o[6346]) );
  AND U12182 ( .A(p_input[26346]), .B(p_input[16346]), .Z(n8122) );
  AND U12183 ( .A(p_input[6346]), .B(p_input[36346]), .Z(n8121) );
  AND U12184 ( .A(n8123), .B(n8124), .Z(o[6345]) );
  AND U12185 ( .A(p_input[26345]), .B(p_input[16345]), .Z(n8124) );
  AND U12186 ( .A(p_input[6345]), .B(p_input[36345]), .Z(n8123) );
  AND U12187 ( .A(n8125), .B(n8126), .Z(o[6344]) );
  AND U12188 ( .A(p_input[26344]), .B(p_input[16344]), .Z(n8126) );
  AND U12189 ( .A(p_input[6344]), .B(p_input[36344]), .Z(n8125) );
  AND U12190 ( .A(n8127), .B(n8128), .Z(o[6343]) );
  AND U12191 ( .A(p_input[26343]), .B(p_input[16343]), .Z(n8128) );
  AND U12192 ( .A(p_input[6343]), .B(p_input[36343]), .Z(n8127) );
  AND U12193 ( .A(n8129), .B(n8130), .Z(o[6342]) );
  AND U12194 ( .A(p_input[26342]), .B(p_input[16342]), .Z(n8130) );
  AND U12195 ( .A(p_input[6342]), .B(p_input[36342]), .Z(n8129) );
  AND U12196 ( .A(n8131), .B(n8132), .Z(o[6341]) );
  AND U12197 ( .A(p_input[26341]), .B(p_input[16341]), .Z(n8132) );
  AND U12198 ( .A(p_input[6341]), .B(p_input[36341]), .Z(n8131) );
  AND U12199 ( .A(n8133), .B(n8134), .Z(o[6340]) );
  AND U12200 ( .A(p_input[26340]), .B(p_input[16340]), .Z(n8134) );
  AND U12201 ( .A(p_input[6340]), .B(p_input[36340]), .Z(n8133) );
  AND U12202 ( .A(n8135), .B(n8136), .Z(o[633]) );
  AND U12203 ( .A(p_input[20633]), .B(p_input[10633]), .Z(n8136) );
  AND U12204 ( .A(p_input[633]), .B(p_input[30633]), .Z(n8135) );
  AND U12205 ( .A(n8137), .B(n8138), .Z(o[6339]) );
  AND U12206 ( .A(p_input[26339]), .B(p_input[16339]), .Z(n8138) );
  AND U12207 ( .A(p_input[6339]), .B(p_input[36339]), .Z(n8137) );
  AND U12208 ( .A(n8139), .B(n8140), .Z(o[6338]) );
  AND U12209 ( .A(p_input[26338]), .B(p_input[16338]), .Z(n8140) );
  AND U12210 ( .A(p_input[6338]), .B(p_input[36338]), .Z(n8139) );
  AND U12211 ( .A(n8141), .B(n8142), .Z(o[6337]) );
  AND U12212 ( .A(p_input[26337]), .B(p_input[16337]), .Z(n8142) );
  AND U12213 ( .A(p_input[6337]), .B(p_input[36337]), .Z(n8141) );
  AND U12214 ( .A(n8143), .B(n8144), .Z(o[6336]) );
  AND U12215 ( .A(p_input[26336]), .B(p_input[16336]), .Z(n8144) );
  AND U12216 ( .A(p_input[6336]), .B(p_input[36336]), .Z(n8143) );
  AND U12217 ( .A(n8145), .B(n8146), .Z(o[6335]) );
  AND U12218 ( .A(p_input[26335]), .B(p_input[16335]), .Z(n8146) );
  AND U12219 ( .A(p_input[6335]), .B(p_input[36335]), .Z(n8145) );
  AND U12220 ( .A(n8147), .B(n8148), .Z(o[6334]) );
  AND U12221 ( .A(p_input[26334]), .B(p_input[16334]), .Z(n8148) );
  AND U12222 ( .A(p_input[6334]), .B(p_input[36334]), .Z(n8147) );
  AND U12223 ( .A(n8149), .B(n8150), .Z(o[6333]) );
  AND U12224 ( .A(p_input[26333]), .B(p_input[16333]), .Z(n8150) );
  AND U12225 ( .A(p_input[6333]), .B(p_input[36333]), .Z(n8149) );
  AND U12226 ( .A(n8151), .B(n8152), .Z(o[6332]) );
  AND U12227 ( .A(p_input[26332]), .B(p_input[16332]), .Z(n8152) );
  AND U12228 ( .A(p_input[6332]), .B(p_input[36332]), .Z(n8151) );
  AND U12229 ( .A(n8153), .B(n8154), .Z(o[6331]) );
  AND U12230 ( .A(p_input[26331]), .B(p_input[16331]), .Z(n8154) );
  AND U12231 ( .A(p_input[6331]), .B(p_input[36331]), .Z(n8153) );
  AND U12232 ( .A(n8155), .B(n8156), .Z(o[6330]) );
  AND U12233 ( .A(p_input[26330]), .B(p_input[16330]), .Z(n8156) );
  AND U12234 ( .A(p_input[6330]), .B(p_input[36330]), .Z(n8155) );
  AND U12235 ( .A(n8157), .B(n8158), .Z(o[632]) );
  AND U12236 ( .A(p_input[20632]), .B(p_input[10632]), .Z(n8158) );
  AND U12237 ( .A(p_input[632]), .B(p_input[30632]), .Z(n8157) );
  AND U12238 ( .A(n8159), .B(n8160), .Z(o[6329]) );
  AND U12239 ( .A(p_input[26329]), .B(p_input[16329]), .Z(n8160) );
  AND U12240 ( .A(p_input[6329]), .B(p_input[36329]), .Z(n8159) );
  AND U12241 ( .A(n8161), .B(n8162), .Z(o[6328]) );
  AND U12242 ( .A(p_input[26328]), .B(p_input[16328]), .Z(n8162) );
  AND U12243 ( .A(p_input[6328]), .B(p_input[36328]), .Z(n8161) );
  AND U12244 ( .A(n8163), .B(n8164), .Z(o[6327]) );
  AND U12245 ( .A(p_input[26327]), .B(p_input[16327]), .Z(n8164) );
  AND U12246 ( .A(p_input[6327]), .B(p_input[36327]), .Z(n8163) );
  AND U12247 ( .A(n8165), .B(n8166), .Z(o[6326]) );
  AND U12248 ( .A(p_input[26326]), .B(p_input[16326]), .Z(n8166) );
  AND U12249 ( .A(p_input[6326]), .B(p_input[36326]), .Z(n8165) );
  AND U12250 ( .A(n8167), .B(n8168), .Z(o[6325]) );
  AND U12251 ( .A(p_input[26325]), .B(p_input[16325]), .Z(n8168) );
  AND U12252 ( .A(p_input[6325]), .B(p_input[36325]), .Z(n8167) );
  AND U12253 ( .A(n8169), .B(n8170), .Z(o[6324]) );
  AND U12254 ( .A(p_input[26324]), .B(p_input[16324]), .Z(n8170) );
  AND U12255 ( .A(p_input[6324]), .B(p_input[36324]), .Z(n8169) );
  AND U12256 ( .A(n8171), .B(n8172), .Z(o[6323]) );
  AND U12257 ( .A(p_input[26323]), .B(p_input[16323]), .Z(n8172) );
  AND U12258 ( .A(p_input[6323]), .B(p_input[36323]), .Z(n8171) );
  AND U12259 ( .A(n8173), .B(n8174), .Z(o[6322]) );
  AND U12260 ( .A(p_input[26322]), .B(p_input[16322]), .Z(n8174) );
  AND U12261 ( .A(p_input[6322]), .B(p_input[36322]), .Z(n8173) );
  AND U12262 ( .A(n8175), .B(n8176), .Z(o[6321]) );
  AND U12263 ( .A(p_input[26321]), .B(p_input[16321]), .Z(n8176) );
  AND U12264 ( .A(p_input[6321]), .B(p_input[36321]), .Z(n8175) );
  AND U12265 ( .A(n8177), .B(n8178), .Z(o[6320]) );
  AND U12266 ( .A(p_input[26320]), .B(p_input[16320]), .Z(n8178) );
  AND U12267 ( .A(p_input[6320]), .B(p_input[36320]), .Z(n8177) );
  AND U12268 ( .A(n8179), .B(n8180), .Z(o[631]) );
  AND U12269 ( .A(p_input[20631]), .B(p_input[10631]), .Z(n8180) );
  AND U12270 ( .A(p_input[631]), .B(p_input[30631]), .Z(n8179) );
  AND U12271 ( .A(n8181), .B(n8182), .Z(o[6319]) );
  AND U12272 ( .A(p_input[26319]), .B(p_input[16319]), .Z(n8182) );
  AND U12273 ( .A(p_input[6319]), .B(p_input[36319]), .Z(n8181) );
  AND U12274 ( .A(n8183), .B(n8184), .Z(o[6318]) );
  AND U12275 ( .A(p_input[26318]), .B(p_input[16318]), .Z(n8184) );
  AND U12276 ( .A(p_input[6318]), .B(p_input[36318]), .Z(n8183) );
  AND U12277 ( .A(n8185), .B(n8186), .Z(o[6317]) );
  AND U12278 ( .A(p_input[26317]), .B(p_input[16317]), .Z(n8186) );
  AND U12279 ( .A(p_input[6317]), .B(p_input[36317]), .Z(n8185) );
  AND U12280 ( .A(n8187), .B(n8188), .Z(o[6316]) );
  AND U12281 ( .A(p_input[26316]), .B(p_input[16316]), .Z(n8188) );
  AND U12282 ( .A(p_input[6316]), .B(p_input[36316]), .Z(n8187) );
  AND U12283 ( .A(n8189), .B(n8190), .Z(o[6315]) );
  AND U12284 ( .A(p_input[26315]), .B(p_input[16315]), .Z(n8190) );
  AND U12285 ( .A(p_input[6315]), .B(p_input[36315]), .Z(n8189) );
  AND U12286 ( .A(n8191), .B(n8192), .Z(o[6314]) );
  AND U12287 ( .A(p_input[26314]), .B(p_input[16314]), .Z(n8192) );
  AND U12288 ( .A(p_input[6314]), .B(p_input[36314]), .Z(n8191) );
  AND U12289 ( .A(n8193), .B(n8194), .Z(o[6313]) );
  AND U12290 ( .A(p_input[26313]), .B(p_input[16313]), .Z(n8194) );
  AND U12291 ( .A(p_input[6313]), .B(p_input[36313]), .Z(n8193) );
  AND U12292 ( .A(n8195), .B(n8196), .Z(o[6312]) );
  AND U12293 ( .A(p_input[26312]), .B(p_input[16312]), .Z(n8196) );
  AND U12294 ( .A(p_input[6312]), .B(p_input[36312]), .Z(n8195) );
  AND U12295 ( .A(n8197), .B(n8198), .Z(o[6311]) );
  AND U12296 ( .A(p_input[26311]), .B(p_input[16311]), .Z(n8198) );
  AND U12297 ( .A(p_input[6311]), .B(p_input[36311]), .Z(n8197) );
  AND U12298 ( .A(n8199), .B(n8200), .Z(o[6310]) );
  AND U12299 ( .A(p_input[26310]), .B(p_input[16310]), .Z(n8200) );
  AND U12300 ( .A(p_input[6310]), .B(p_input[36310]), .Z(n8199) );
  AND U12301 ( .A(n8201), .B(n8202), .Z(o[630]) );
  AND U12302 ( .A(p_input[20630]), .B(p_input[10630]), .Z(n8202) );
  AND U12303 ( .A(p_input[630]), .B(p_input[30630]), .Z(n8201) );
  AND U12304 ( .A(n8203), .B(n8204), .Z(o[6309]) );
  AND U12305 ( .A(p_input[26309]), .B(p_input[16309]), .Z(n8204) );
  AND U12306 ( .A(p_input[6309]), .B(p_input[36309]), .Z(n8203) );
  AND U12307 ( .A(n8205), .B(n8206), .Z(o[6308]) );
  AND U12308 ( .A(p_input[26308]), .B(p_input[16308]), .Z(n8206) );
  AND U12309 ( .A(p_input[6308]), .B(p_input[36308]), .Z(n8205) );
  AND U12310 ( .A(n8207), .B(n8208), .Z(o[6307]) );
  AND U12311 ( .A(p_input[26307]), .B(p_input[16307]), .Z(n8208) );
  AND U12312 ( .A(p_input[6307]), .B(p_input[36307]), .Z(n8207) );
  AND U12313 ( .A(n8209), .B(n8210), .Z(o[6306]) );
  AND U12314 ( .A(p_input[26306]), .B(p_input[16306]), .Z(n8210) );
  AND U12315 ( .A(p_input[6306]), .B(p_input[36306]), .Z(n8209) );
  AND U12316 ( .A(n8211), .B(n8212), .Z(o[6305]) );
  AND U12317 ( .A(p_input[26305]), .B(p_input[16305]), .Z(n8212) );
  AND U12318 ( .A(p_input[6305]), .B(p_input[36305]), .Z(n8211) );
  AND U12319 ( .A(n8213), .B(n8214), .Z(o[6304]) );
  AND U12320 ( .A(p_input[26304]), .B(p_input[16304]), .Z(n8214) );
  AND U12321 ( .A(p_input[6304]), .B(p_input[36304]), .Z(n8213) );
  AND U12322 ( .A(n8215), .B(n8216), .Z(o[6303]) );
  AND U12323 ( .A(p_input[26303]), .B(p_input[16303]), .Z(n8216) );
  AND U12324 ( .A(p_input[6303]), .B(p_input[36303]), .Z(n8215) );
  AND U12325 ( .A(n8217), .B(n8218), .Z(o[6302]) );
  AND U12326 ( .A(p_input[26302]), .B(p_input[16302]), .Z(n8218) );
  AND U12327 ( .A(p_input[6302]), .B(p_input[36302]), .Z(n8217) );
  AND U12328 ( .A(n8219), .B(n8220), .Z(o[6301]) );
  AND U12329 ( .A(p_input[26301]), .B(p_input[16301]), .Z(n8220) );
  AND U12330 ( .A(p_input[6301]), .B(p_input[36301]), .Z(n8219) );
  AND U12331 ( .A(n8221), .B(n8222), .Z(o[6300]) );
  AND U12332 ( .A(p_input[26300]), .B(p_input[16300]), .Z(n8222) );
  AND U12333 ( .A(p_input[6300]), .B(p_input[36300]), .Z(n8221) );
  AND U12334 ( .A(n8223), .B(n8224), .Z(o[62]) );
  AND U12335 ( .A(p_input[20062]), .B(p_input[10062]), .Z(n8224) );
  AND U12336 ( .A(p_input[62]), .B(p_input[30062]), .Z(n8223) );
  AND U12337 ( .A(n8225), .B(n8226), .Z(o[629]) );
  AND U12338 ( .A(p_input[20629]), .B(p_input[10629]), .Z(n8226) );
  AND U12339 ( .A(p_input[629]), .B(p_input[30629]), .Z(n8225) );
  AND U12340 ( .A(n8227), .B(n8228), .Z(o[6299]) );
  AND U12341 ( .A(p_input[26299]), .B(p_input[16299]), .Z(n8228) );
  AND U12342 ( .A(p_input[6299]), .B(p_input[36299]), .Z(n8227) );
  AND U12343 ( .A(n8229), .B(n8230), .Z(o[6298]) );
  AND U12344 ( .A(p_input[26298]), .B(p_input[16298]), .Z(n8230) );
  AND U12345 ( .A(p_input[6298]), .B(p_input[36298]), .Z(n8229) );
  AND U12346 ( .A(n8231), .B(n8232), .Z(o[6297]) );
  AND U12347 ( .A(p_input[26297]), .B(p_input[16297]), .Z(n8232) );
  AND U12348 ( .A(p_input[6297]), .B(p_input[36297]), .Z(n8231) );
  AND U12349 ( .A(n8233), .B(n8234), .Z(o[6296]) );
  AND U12350 ( .A(p_input[26296]), .B(p_input[16296]), .Z(n8234) );
  AND U12351 ( .A(p_input[6296]), .B(p_input[36296]), .Z(n8233) );
  AND U12352 ( .A(n8235), .B(n8236), .Z(o[6295]) );
  AND U12353 ( .A(p_input[26295]), .B(p_input[16295]), .Z(n8236) );
  AND U12354 ( .A(p_input[6295]), .B(p_input[36295]), .Z(n8235) );
  AND U12355 ( .A(n8237), .B(n8238), .Z(o[6294]) );
  AND U12356 ( .A(p_input[26294]), .B(p_input[16294]), .Z(n8238) );
  AND U12357 ( .A(p_input[6294]), .B(p_input[36294]), .Z(n8237) );
  AND U12358 ( .A(n8239), .B(n8240), .Z(o[6293]) );
  AND U12359 ( .A(p_input[26293]), .B(p_input[16293]), .Z(n8240) );
  AND U12360 ( .A(p_input[6293]), .B(p_input[36293]), .Z(n8239) );
  AND U12361 ( .A(n8241), .B(n8242), .Z(o[6292]) );
  AND U12362 ( .A(p_input[26292]), .B(p_input[16292]), .Z(n8242) );
  AND U12363 ( .A(p_input[6292]), .B(p_input[36292]), .Z(n8241) );
  AND U12364 ( .A(n8243), .B(n8244), .Z(o[6291]) );
  AND U12365 ( .A(p_input[26291]), .B(p_input[16291]), .Z(n8244) );
  AND U12366 ( .A(p_input[6291]), .B(p_input[36291]), .Z(n8243) );
  AND U12367 ( .A(n8245), .B(n8246), .Z(o[6290]) );
  AND U12368 ( .A(p_input[26290]), .B(p_input[16290]), .Z(n8246) );
  AND U12369 ( .A(p_input[6290]), .B(p_input[36290]), .Z(n8245) );
  AND U12370 ( .A(n8247), .B(n8248), .Z(o[628]) );
  AND U12371 ( .A(p_input[20628]), .B(p_input[10628]), .Z(n8248) );
  AND U12372 ( .A(p_input[628]), .B(p_input[30628]), .Z(n8247) );
  AND U12373 ( .A(n8249), .B(n8250), .Z(o[6289]) );
  AND U12374 ( .A(p_input[26289]), .B(p_input[16289]), .Z(n8250) );
  AND U12375 ( .A(p_input[6289]), .B(p_input[36289]), .Z(n8249) );
  AND U12376 ( .A(n8251), .B(n8252), .Z(o[6288]) );
  AND U12377 ( .A(p_input[26288]), .B(p_input[16288]), .Z(n8252) );
  AND U12378 ( .A(p_input[6288]), .B(p_input[36288]), .Z(n8251) );
  AND U12379 ( .A(n8253), .B(n8254), .Z(o[6287]) );
  AND U12380 ( .A(p_input[26287]), .B(p_input[16287]), .Z(n8254) );
  AND U12381 ( .A(p_input[6287]), .B(p_input[36287]), .Z(n8253) );
  AND U12382 ( .A(n8255), .B(n8256), .Z(o[6286]) );
  AND U12383 ( .A(p_input[26286]), .B(p_input[16286]), .Z(n8256) );
  AND U12384 ( .A(p_input[6286]), .B(p_input[36286]), .Z(n8255) );
  AND U12385 ( .A(n8257), .B(n8258), .Z(o[6285]) );
  AND U12386 ( .A(p_input[26285]), .B(p_input[16285]), .Z(n8258) );
  AND U12387 ( .A(p_input[6285]), .B(p_input[36285]), .Z(n8257) );
  AND U12388 ( .A(n8259), .B(n8260), .Z(o[6284]) );
  AND U12389 ( .A(p_input[26284]), .B(p_input[16284]), .Z(n8260) );
  AND U12390 ( .A(p_input[6284]), .B(p_input[36284]), .Z(n8259) );
  AND U12391 ( .A(n8261), .B(n8262), .Z(o[6283]) );
  AND U12392 ( .A(p_input[26283]), .B(p_input[16283]), .Z(n8262) );
  AND U12393 ( .A(p_input[6283]), .B(p_input[36283]), .Z(n8261) );
  AND U12394 ( .A(n8263), .B(n8264), .Z(o[6282]) );
  AND U12395 ( .A(p_input[26282]), .B(p_input[16282]), .Z(n8264) );
  AND U12396 ( .A(p_input[6282]), .B(p_input[36282]), .Z(n8263) );
  AND U12397 ( .A(n8265), .B(n8266), .Z(o[6281]) );
  AND U12398 ( .A(p_input[26281]), .B(p_input[16281]), .Z(n8266) );
  AND U12399 ( .A(p_input[6281]), .B(p_input[36281]), .Z(n8265) );
  AND U12400 ( .A(n8267), .B(n8268), .Z(o[6280]) );
  AND U12401 ( .A(p_input[26280]), .B(p_input[16280]), .Z(n8268) );
  AND U12402 ( .A(p_input[6280]), .B(p_input[36280]), .Z(n8267) );
  AND U12403 ( .A(n8269), .B(n8270), .Z(o[627]) );
  AND U12404 ( .A(p_input[20627]), .B(p_input[10627]), .Z(n8270) );
  AND U12405 ( .A(p_input[627]), .B(p_input[30627]), .Z(n8269) );
  AND U12406 ( .A(n8271), .B(n8272), .Z(o[6279]) );
  AND U12407 ( .A(p_input[26279]), .B(p_input[16279]), .Z(n8272) );
  AND U12408 ( .A(p_input[6279]), .B(p_input[36279]), .Z(n8271) );
  AND U12409 ( .A(n8273), .B(n8274), .Z(o[6278]) );
  AND U12410 ( .A(p_input[26278]), .B(p_input[16278]), .Z(n8274) );
  AND U12411 ( .A(p_input[6278]), .B(p_input[36278]), .Z(n8273) );
  AND U12412 ( .A(n8275), .B(n8276), .Z(o[6277]) );
  AND U12413 ( .A(p_input[26277]), .B(p_input[16277]), .Z(n8276) );
  AND U12414 ( .A(p_input[6277]), .B(p_input[36277]), .Z(n8275) );
  AND U12415 ( .A(n8277), .B(n8278), .Z(o[6276]) );
  AND U12416 ( .A(p_input[26276]), .B(p_input[16276]), .Z(n8278) );
  AND U12417 ( .A(p_input[6276]), .B(p_input[36276]), .Z(n8277) );
  AND U12418 ( .A(n8279), .B(n8280), .Z(o[6275]) );
  AND U12419 ( .A(p_input[26275]), .B(p_input[16275]), .Z(n8280) );
  AND U12420 ( .A(p_input[6275]), .B(p_input[36275]), .Z(n8279) );
  AND U12421 ( .A(n8281), .B(n8282), .Z(o[6274]) );
  AND U12422 ( .A(p_input[26274]), .B(p_input[16274]), .Z(n8282) );
  AND U12423 ( .A(p_input[6274]), .B(p_input[36274]), .Z(n8281) );
  AND U12424 ( .A(n8283), .B(n8284), .Z(o[6273]) );
  AND U12425 ( .A(p_input[26273]), .B(p_input[16273]), .Z(n8284) );
  AND U12426 ( .A(p_input[6273]), .B(p_input[36273]), .Z(n8283) );
  AND U12427 ( .A(n8285), .B(n8286), .Z(o[6272]) );
  AND U12428 ( .A(p_input[26272]), .B(p_input[16272]), .Z(n8286) );
  AND U12429 ( .A(p_input[6272]), .B(p_input[36272]), .Z(n8285) );
  AND U12430 ( .A(n8287), .B(n8288), .Z(o[6271]) );
  AND U12431 ( .A(p_input[26271]), .B(p_input[16271]), .Z(n8288) );
  AND U12432 ( .A(p_input[6271]), .B(p_input[36271]), .Z(n8287) );
  AND U12433 ( .A(n8289), .B(n8290), .Z(o[6270]) );
  AND U12434 ( .A(p_input[26270]), .B(p_input[16270]), .Z(n8290) );
  AND U12435 ( .A(p_input[6270]), .B(p_input[36270]), .Z(n8289) );
  AND U12436 ( .A(n8291), .B(n8292), .Z(o[626]) );
  AND U12437 ( .A(p_input[20626]), .B(p_input[10626]), .Z(n8292) );
  AND U12438 ( .A(p_input[626]), .B(p_input[30626]), .Z(n8291) );
  AND U12439 ( .A(n8293), .B(n8294), .Z(o[6269]) );
  AND U12440 ( .A(p_input[26269]), .B(p_input[16269]), .Z(n8294) );
  AND U12441 ( .A(p_input[6269]), .B(p_input[36269]), .Z(n8293) );
  AND U12442 ( .A(n8295), .B(n8296), .Z(o[6268]) );
  AND U12443 ( .A(p_input[26268]), .B(p_input[16268]), .Z(n8296) );
  AND U12444 ( .A(p_input[6268]), .B(p_input[36268]), .Z(n8295) );
  AND U12445 ( .A(n8297), .B(n8298), .Z(o[6267]) );
  AND U12446 ( .A(p_input[26267]), .B(p_input[16267]), .Z(n8298) );
  AND U12447 ( .A(p_input[6267]), .B(p_input[36267]), .Z(n8297) );
  AND U12448 ( .A(n8299), .B(n8300), .Z(o[6266]) );
  AND U12449 ( .A(p_input[26266]), .B(p_input[16266]), .Z(n8300) );
  AND U12450 ( .A(p_input[6266]), .B(p_input[36266]), .Z(n8299) );
  AND U12451 ( .A(n8301), .B(n8302), .Z(o[6265]) );
  AND U12452 ( .A(p_input[26265]), .B(p_input[16265]), .Z(n8302) );
  AND U12453 ( .A(p_input[6265]), .B(p_input[36265]), .Z(n8301) );
  AND U12454 ( .A(n8303), .B(n8304), .Z(o[6264]) );
  AND U12455 ( .A(p_input[26264]), .B(p_input[16264]), .Z(n8304) );
  AND U12456 ( .A(p_input[6264]), .B(p_input[36264]), .Z(n8303) );
  AND U12457 ( .A(n8305), .B(n8306), .Z(o[6263]) );
  AND U12458 ( .A(p_input[26263]), .B(p_input[16263]), .Z(n8306) );
  AND U12459 ( .A(p_input[6263]), .B(p_input[36263]), .Z(n8305) );
  AND U12460 ( .A(n8307), .B(n8308), .Z(o[6262]) );
  AND U12461 ( .A(p_input[26262]), .B(p_input[16262]), .Z(n8308) );
  AND U12462 ( .A(p_input[6262]), .B(p_input[36262]), .Z(n8307) );
  AND U12463 ( .A(n8309), .B(n8310), .Z(o[6261]) );
  AND U12464 ( .A(p_input[26261]), .B(p_input[16261]), .Z(n8310) );
  AND U12465 ( .A(p_input[6261]), .B(p_input[36261]), .Z(n8309) );
  AND U12466 ( .A(n8311), .B(n8312), .Z(o[6260]) );
  AND U12467 ( .A(p_input[26260]), .B(p_input[16260]), .Z(n8312) );
  AND U12468 ( .A(p_input[6260]), .B(p_input[36260]), .Z(n8311) );
  AND U12469 ( .A(n8313), .B(n8314), .Z(o[625]) );
  AND U12470 ( .A(p_input[20625]), .B(p_input[10625]), .Z(n8314) );
  AND U12471 ( .A(p_input[625]), .B(p_input[30625]), .Z(n8313) );
  AND U12472 ( .A(n8315), .B(n8316), .Z(o[6259]) );
  AND U12473 ( .A(p_input[26259]), .B(p_input[16259]), .Z(n8316) );
  AND U12474 ( .A(p_input[6259]), .B(p_input[36259]), .Z(n8315) );
  AND U12475 ( .A(n8317), .B(n8318), .Z(o[6258]) );
  AND U12476 ( .A(p_input[26258]), .B(p_input[16258]), .Z(n8318) );
  AND U12477 ( .A(p_input[6258]), .B(p_input[36258]), .Z(n8317) );
  AND U12478 ( .A(n8319), .B(n8320), .Z(o[6257]) );
  AND U12479 ( .A(p_input[26257]), .B(p_input[16257]), .Z(n8320) );
  AND U12480 ( .A(p_input[6257]), .B(p_input[36257]), .Z(n8319) );
  AND U12481 ( .A(n8321), .B(n8322), .Z(o[6256]) );
  AND U12482 ( .A(p_input[26256]), .B(p_input[16256]), .Z(n8322) );
  AND U12483 ( .A(p_input[6256]), .B(p_input[36256]), .Z(n8321) );
  AND U12484 ( .A(n8323), .B(n8324), .Z(o[6255]) );
  AND U12485 ( .A(p_input[26255]), .B(p_input[16255]), .Z(n8324) );
  AND U12486 ( .A(p_input[6255]), .B(p_input[36255]), .Z(n8323) );
  AND U12487 ( .A(n8325), .B(n8326), .Z(o[6254]) );
  AND U12488 ( .A(p_input[26254]), .B(p_input[16254]), .Z(n8326) );
  AND U12489 ( .A(p_input[6254]), .B(p_input[36254]), .Z(n8325) );
  AND U12490 ( .A(n8327), .B(n8328), .Z(o[6253]) );
  AND U12491 ( .A(p_input[26253]), .B(p_input[16253]), .Z(n8328) );
  AND U12492 ( .A(p_input[6253]), .B(p_input[36253]), .Z(n8327) );
  AND U12493 ( .A(n8329), .B(n8330), .Z(o[6252]) );
  AND U12494 ( .A(p_input[26252]), .B(p_input[16252]), .Z(n8330) );
  AND U12495 ( .A(p_input[6252]), .B(p_input[36252]), .Z(n8329) );
  AND U12496 ( .A(n8331), .B(n8332), .Z(o[6251]) );
  AND U12497 ( .A(p_input[26251]), .B(p_input[16251]), .Z(n8332) );
  AND U12498 ( .A(p_input[6251]), .B(p_input[36251]), .Z(n8331) );
  AND U12499 ( .A(n8333), .B(n8334), .Z(o[6250]) );
  AND U12500 ( .A(p_input[26250]), .B(p_input[16250]), .Z(n8334) );
  AND U12501 ( .A(p_input[6250]), .B(p_input[36250]), .Z(n8333) );
  AND U12502 ( .A(n8335), .B(n8336), .Z(o[624]) );
  AND U12503 ( .A(p_input[20624]), .B(p_input[10624]), .Z(n8336) );
  AND U12504 ( .A(p_input[624]), .B(p_input[30624]), .Z(n8335) );
  AND U12505 ( .A(n8337), .B(n8338), .Z(o[6249]) );
  AND U12506 ( .A(p_input[26249]), .B(p_input[16249]), .Z(n8338) );
  AND U12507 ( .A(p_input[6249]), .B(p_input[36249]), .Z(n8337) );
  AND U12508 ( .A(n8339), .B(n8340), .Z(o[6248]) );
  AND U12509 ( .A(p_input[26248]), .B(p_input[16248]), .Z(n8340) );
  AND U12510 ( .A(p_input[6248]), .B(p_input[36248]), .Z(n8339) );
  AND U12511 ( .A(n8341), .B(n8342), .Z(o[6247]) );
  AND U12512 ( .A(p_input[26247]), .B(p_input[16247]), .Z(n8342) );
  AND U12513 ( .A(p_input[6247]), .B(p_input[36247]), .Z(n8341) );
  AND U12514 ( .A(n8343), .B(n8344), .Z(o[6246]) );
  AND U12515 ( .A(p_input[26246]), .B(p_input[16246]), .Z(n8344) );
  AND U12516 ( .A(p_input[6246]), .B(p_input[36246]), .Z(n8343) );
  AND U12517 ( .A(n8345), .B(n8346), .Z(o[6245]) );
  AND U12518 ( .A(p_input[26245]), .B(p_input[16245]), .Z(n8346) );
  AND U12519 ( .A(p_input[6245]), .B(p_input[36245]), .Z(n8345) );
  AND U12520 ( .A(n8347), .B(n8348), .Z(o[6244]) );
  AND U12521 ( .A(p_input[26244]), .B(p_input[16244]), .Z(n8348) );
  AND U12522 ( .A(p_input[6244]), .B(p_input[36244]), .Z(n8347) );
  AND U12523 ( .A(n8349), .B(n8350), .Z(o[6243]) );
  AND U12524 ( .A(p_input[26243]), .B(p_input[16243]), .Z(n8350) );
  AND U12525 ( .A(p_input[6243]), .B(p_input[36243]), .Z(n8349) );
  AND U12526 ( .A(n8351), .B(n8352), .Z(o[6242]) );
  AND U12527 ( .A(p_input[26242]), .B(p_input[16242]), .Z(n8352) );
  AND U12528 ( .A(p_input[6242]), .B(p_input[36242]), .Z(n8351) );
  AND U12529 ( .A(n8353), .B(n8354), .Z(o[6241]) );
  AND U12530 ( .A(p_input[26241]), .B(p_input[16241]), .Z(n8354) );
  AND U12531 ( .A(p_input[6241]), .B(p_input[36241]), .Z(n8353) );
  AND U12532 ( .A(n8355), .B(n8356), .Z(o[6240]) );
  AND U12533 ( .A(p_input[26240]), .B(p_input[16240]), .Z(n8356) );
  AND U12534 ( .A(p_input[6240]), .B(p_input[36240]), .Z(n8355) );
  AND U12535 ( .A(n8357), .B(n8358), .Z(o[623]) );
  AND U12536 ( .A(p_input[20623]), .B(p_input[10623]), .Z(n8358) );
  AND U12537 ( .A(p_input[623]), .B(p_input[30623]), .Z(n8357) );
  AND U12538 ( .A(n8359), .B(n8360), .Z(o[6239]) );
  AND U12539 ( .A(p_input[26239]), .B(p_input[16239]), .Z(n8360) );
  AND U12540 ( .A(p_input[6239]), .B(p_input[36239]), .Z(n8359) );
  AND U12541 ( .A(n8361), .B(n8362), .Z(o[6238]) );
  AND U12542 ( .A(p_input[26238]), .B(p_input[16238]), .Z(n8362) );
  AND U12543 ( .A(p_input[6238]), .B(p_input[36238]), .Z(n8361) );
  AND U12544 ( .A(n8363), .B(n8364), .Z(o[6237]) );
  AND U12545 ( .A(p_input[26237]), .B(p_input[16237]), .Z(n8364) );
  AND U12546 ( .A(p_input[6237]), .B(p_input[36237]), .Z(n8363) );
  AND U12547 ( .A(n8365), .B(n8366), .Z(o[6236]) );
  AND U12548 ( .A(p_input[26236]), .B(p_input[16236]), .Z(n8366) );
  AND U12549 ( .A(p_input[6236]), .B(p_input[36236]), .Z(n8365) );
  AND U12550 ( .A(n8367), .B(n8368), .Z(o[6235]) );
  AND U12551 ( .A(p_input[26235]), .B(p_input[16235]), .Z(n8368) );
  AND U12552 ( .A(p_input[6235]), .B(p_input[36235]), .Z(n8367) );
  AND U12553 ( .A(n8369), .B(n8370), .Z(o[6234]) );
  AND U12554 ( .A(p_input[26234]), .B(p_input[16234]), .Z(n8370) );
  AND U12555 ( .A(p_input[6234]), .B(p_input[36234]), .Z(n8369) );
  AND U12556 ( .A(n8371), .B(n8372), .Z(o[6233]) );
  AND U12557 ( .A(p_input[26233]), .B(p_input[16233]), .Z(n8372) );
  AND U12558 ( .A(p_input[6233]), .B(p_input[36233]), .Z(n8371) );
  AND U12559 ( .A(n8373), .B(n8374), .Z(o[6232]) );
  AND U12560 ( .A(p_input[26232]), .B(p_input[16232]), .Z(n8374) );
  AND U12561 ( .A(p_input[6232]), .B(p_input[36232]), .Z(n8373) );
  AND U12562 ( .A(n8375), .B(n8376), .Z(o[6231]) );
  AND U12563 ( .A(p_input[26231]), .B(p_input[16231]), .Z(n8376) );
  AND U12564 ( .A(p_input[6231]), .B(p_input[36231]), .Z(n8375) );
  AND U12565 ( .A(n8377), .B(n8378), .Z(o[6230]) );
  AND U12566 ( .A(p_input[26230]), .B(p_input[16230]), .Z(n8378) );
  AND U12567 ( .A(p_input[6230]), .B(p_input[36230]), .Z(n8377) );
  AND U12568 ( .A(n8379), .B(n8380), .Z(o[622]) );
  AND U12569 ( .A(p_input[20622]), .B(p_input[10622]), .Z(n8380) );
  AND U12570 ( .A(p_input[622]), .B(p_input[30622]), .Z(n8379) );
  AND U12571 ( .A(n8381), .B(n8382), .Z(o[6229]) );
  AND U12572 ( .A(p_input[26229]), .B(p_input[16229]), .Z(n8382) );
  AND U12573 ( .A(p_input[6229]), .B(p_input[36229]), .Z(n8381) );
  AND U12574 ( .A(n8383), .B(n8384), .Z(o[6228]) );
  AND U12575 ( .A(p_input[26228]), .B(p_input[16228]), .Z(n8384) );
  AND U12576 ( .A(p_input[6228]), .B(p_input[36228]), .Z(n8383) );
  AND U12577 ( .A(n8385), .B(n8386), .Z(o[6227]) );
  AND U12578 ( .A(p_input[26227]), .B(p_input[16227]), .Z(n8386) );
  AND U12579 ( .A(p_input[6227]), .B(p_input[36227]), .Z(n8385) );
  AND U12580 ( .A(n8387), .B(n8388), .Z(o[6226]) );
  AND U12581 ( .A(p_input[26226]), .B(p_input[16226]), .Z(n8388) );
  AND U12582 ( .A(p_input[6226]), .B(p_input[36226]), .Z(n8387) );
  AND U12583 ( .A(n8389), .B(n8390), .Z(o[6225]) );
  AND U12584 ( .A(p_input[26225]), .B(p_input[16225]), .Z(n8390) );
  AND U12585 ( .A(p_input[6225]), .B(p_input[36225]), .Z(n8389) );
  AND U12586 ( .A(n8391), .B(n8392), .Z(o[6224]) );
  AND U12587 ( .A(p_input[26224]), .B(p_input[16224]), .Z(n8392) );
  AND U12588 ( .A(p_input[6224]), .B(p_input[36224]), .Z(n8391) );
  AND U12589 ( .A(n8393), .B(n8394), .Z(o[6223]) );
  AND U12590 ( .A(p_input[26223]), .B(p_input[16223]), .Z(n8394) );
  AND U12591 ( .A(p_input[6223]), .B(p_input[36223]), .Z(n8393) );
  AND U12592 ( .A(n8395), .B(n8396), .Z(o[6222]) );
  AND U12593 ( .A(p_input[26222]), .B(p_input[16222]), .Z(n8396) );
  AND U12594 ( .A(p_input[6222]), .B(p_input[36222]), .Z(n8395) );
  AND U12595 ( .A(n8397), .B(n8398), .Z(o[6221]) );
  AND U12596 ( .A(p_input[26221]), .B(p_input[16221]), .Z(n8398) );
  AND U12597 ( .A(p_input[6221]), .B(p_input[36221]), .Z(n8397) );
  AND U12598 ( .A(n8399), .B(n8400), .Z(o[6220]) );
  AND U12599 ( .A(p_input[26220]), .B(p_input[16220]), .Z(n8400) );
  AND U12600 ( .A(p_input[6220]), .B(p_input[36220]), .Z(n8399) );
  AND U12601 ( .A(n8401), .B(n8402), .Z(o[621]) );
  AND U12602 ( .A(p_input[20621]), .B(p_input[10621]), .Z(n8402) );
  AND U12603 ( .A(p_input[621]), .B(p_input[30621]), .Z(n8401) );
  AND U12604 ( .A(n8403), .B(n8404), .Z(o[6219]) );
  AND U12605 ( .A(p_input[26219]), .B(p_input[16219]), .Z(n8404) );
  AND U12606 ( .A(p_input[6219]), .B(p_input[36219]), .Z(n8403) );
  AND U12607 ( .A(n8405), .B(n8406), .Z(o[6218]) );
  AND U12608 ( .A(p_input[26218]), .B(p_input[16218]), .Z(n8406) );
  AND U12609 ( .A(p_input[6218]), .B(p_input[36218]), .Z(n8405) );
  AND U12610 ( .A(n8407), .B(n8408), .Z(o[6217]) );
  AND U12611 ( .A(p_input[26217]), .B(p_input[16217]), .Z(n8408) );
  AND U12612 ( .A(p_input[6217]), .B(p_input[36217]), .Z(n8407) );
  AND U12613 ( .A(n8409), .B(n8410), .Z(o[6216]) );
  AND U12614 ( .A(p_input[26216]), .B(p_input[16216]), .Z(n8410) );
  AND U12615 ( .A(p_input[6216]), .B(p_input[36216]), .Z(n8409) );
  AND U12616 ( .A(n8411), .B(n8412), .Z(o[6215]) );
  AND U12617 ( .A(p_input[26215]), .B(p_input[16215]), .Z(n8412) );
  AND U12618 ( .A(p_input[6215]), .B(p_input[36215]), .Z(n8411) );
  AND U12619 ( .A(n8413), .B(n8414), .Z(o[6214]) );
  AND U12620 ( .A(p_input[26214]), .B(p_input[16214]), .Z(n8414) );
  AND U12621 ( .A(p_input[6214]), .B(p_input[36214]), .Z(n8413) );
  AND U12622 ( .A(n8415), .B(n8416), .Z(o[6213]) );
  AND U12623 ( .A(p_input[26213]), .B(p_input[16213]), .Z(n8416) );
  AND U12624 ( .A(p_input[6213]), .B(p_input[36213]), .Z(n8415) );
  AND U12625 ( .A(n8417), .B(n8418), .Z(o[6212]) );
  AND U12626 ( .A(p_input[26212]), .B(p_input[16212]), .Z(n8418) );
  AND U12627 ( .A(p_input[6212]), .B(p_input[36212]), .Z(n8417) );
  AND U12628 ( .A(n8419), .B(n8420), .Z(o[6211]) );
  AND U12629 ( .A(p_input[26211]), .B(p_input[16211]), .Z(n8420) );
  AND U12630 ( .A(p_input[6211]), .B(p_input[36211]), .Z(n8419) );
  AND U12631 ( .A(n8421), .B(n8422), .Z(o[6210]) );
  AND U12632 ( .A(p_input[26210]), .B(p_input[16210]), .Z(n8422) );
  AND U12633 ( .A(p_input[6210]), .B(p_input[36210]), .Z(n8421) );
  AND U12634 ( .A(n8423), .B(n8424), .Z(o[620]) );
  AND U12635 ( .A(p_input[20620]), .B(p_input[10620]), .Z(n8424) );
  AND U12636 ( .A(p_input[620]), .B(p_input[30620]), .Z(n8423) );
  AND U12637 ( .A(n8425), .B(n8426), .Z(o[6209]) );
  AND U12638 ( .A(p_input[26209]), .B(p_input[16209]), .Z(n8426) );
  AND U12639 ( .A(p_input[6209]), .B(p_input[36209]), .Z(n8425) );
  AND U12640 ( .A(n8427), .B(n8428), .Z(o[6208]) );
  AND U12641 ( .A(p_input[26208]), .B(p_input[16208]), .Z(n8428) );
  AND U12642 ( .A(p_input[6208]), .B(p_input[36208]), .Z(n8427) );
  AND U12643 ( .A(n8429), .B(n8430), .Z(o[6207]) );
  AND U12644 ( .A(p_input[26207]), .B(p_input[16207]), .Z(n8430) );
  AND U12645 ( .A(p_input[6207]), .B(p_input[36207]), .Z(n8429) );
  AND U12646 ( .A(n8431), .B(n8432), .Z(o[6206]) );
  AND U12647 ( .A(p_input[26206]), .B(p_input[16206]), .Z(n8432) );
  AND U12648 ( .A(p_input[6206]), .B(p_input[36206]), .Z(n8431) );
  AND U12649 ( .A(n8433), .B(n8434), .Z(o[6205]) );
  AND U12650 ( .A(p_input[26205]), .B(p_input[16205]), .Z(n8434) );
  AND U12651 ( .A(p_input[6205]), .B(p_input[36205]), .Z(n8433) );
  AND U12652 ( .A(n8435), .B(n8436), .Z(o[6204]) );
  AND U12653 ( .A(p_input[26204]), .B(p_input[16204]), .Z(n8436) );
  AND U12654 ( .A(p_input[6204]), .B(p_input[36204]), .Z(n8435) );
  AND U12655 ( .A(n8437), .B(n8438), .Z(o[6203]) );
  AND U12656 ( .A(p_input[26203]), .B(p_input[16203]), .Z(n8438) );
  AND U12657 ( .A(p_input[6203]), .B(p_input[36203]), .Z(n8437) );
  AND U12658 ( .A(n8439), .B(n8440), .Z(o[6202]) );
  AND U12659 ( .A(p_input[26202]), .B(p_input[16202]), .Z(n8440) );
  AND U12660 ( .A(p_input[6202]), .B(p_input[36202]), .Z(n8439) );
  AND U12661 ( .A(n8441), .B(n8442), .Z(o[6201]) );
  AND U12662 ( .A(p_input[26201]), .B(p_input[16201]), .Z(n8442) );
  AND U12663 ( .A(p_input[6201]), .B(p_input[36201]), .Z(n8441) );
  AND U12664 ( .A(n8443), .B(n8444), .Z(o[6200]) );
  AND U12665 ( .A(p_input[26200]), .B(p_input[16200]), .Z(n8444) );
  AND U12666 ( .A(p_input[6200]), .B(p_input[36200]), .Z(n8443) );
  AND U12667 ( .A(n8445), .B(n8446), .Z(o[61]) );
  AND U12668 ( .A(p_input[20061]), .B(p_input[10061]), .Z(n8446) );
  AND U12669 ( .A(p_input[61]), .B(p_input[30061]), .Z(n8445) );
  AND U12670 ( .A(n8447), .B(n8448), .Z(o[619]) );
  AND U12671 ( .A(p_input[20619]), .B(p_input[10619]), .Z(n8448) );
  AND U12672 ( .A(p_input[619]), .B(p_input[30619]), .Z(n8447) );
  AND U12673 ( .A(n8449), .B(n8450), .Z(o[6199]) );
  AND U12674 ( .A(p_input[26199]), .B(p_input[16199]), .Z(n8450) );
  AND U12675 ( .A(p_input[6199]), .B(p_input[36199]), .Z(n8449) );
  AND U12676 ( .A(n8451), .B(n8452), .Z(o[6198]) );
  AND U12677 ( .A(p_input[26198]), .B(p_input[16198]), .Z(n8452) );
  AND U12678 ( .A(p_input[6198]), .B(p_input[36198]), .Z(n8451) );
  AND U12679 ( .A(n8453), .B(n8454), .Z(o[6197]) );
  AND U12680 ( .A(p_input[26197]), .B(p_input[16197]), .Z(n8454) );
  AND U12681 ( .A(p_input[6197]), .B(p_input[36197]), .Z(n8453) );
  AND U12682 ( .A(n8455), .B(n8456), .Z(o[6196]) );
  AND U12683 ( .A(p_input[26196]), .B(p_input[16196]), .Z(n8456) );
  AND U12684 ( .A(p_input[6196]), .B(p_input[36196]), .Z(n8455) );
  AND U12685 ( .A(n8457), .B(n8458), .Z(o[6195]) );
  AND U12686 ( .A(p_input[26195]), .B(p_input[16195]), .Z(n8458) );
  AND U12687 ( .A(p_input[6195]), .B(p_input[36195]), .Z(n8457) );
  AND U12688 ( .A(n8459), .B(n8460), .Z(o[6194]) );
  AND U12689 ( .A(p_input[26194]), .B(p_input[16194]), .Z(n8460) );
  AND U12690 ( .A(p_input[6194]), .B(p_input[36194]), .Z(n8459) );
  AND U12691 ( .A(n8461), .B(n8462), .Z(o[6193]) );
  AND U12692 ( .A(p_input[26193]), .B(p_input[16193]), .Z(n8462) );
  AND U12693 ( .A(p_input[6193]), .B(p_input[36193]), .Z(n8461) );
  AND U12694 ( .A(n8463), .B(n8464), .Z(o[6192]) );
  AND U12695 ( .A(p_input[26192]), .B(p_input[16192]), .Z(n8464) );
  AND U12696 ( .A(p_input[6192]), .B(p_input[36192]), .Z(n8463) );
  AND U12697 ( .A(n8465), .B(n8466), .Z(o[6191]) );
  AND U12698 ( .A(p_input[26191]), .B(p_input[16191]), .Z(n8466) );
  AND U12699 ( .A(p_input[6191]), .B(p_input[36191]), .Z(n8465) );
  AND U12700 ( .A(n8467), .B(n8468), .Z(o[6190]) );
  AND U12701 ( .A(p_input[26190]), .B(p_input[16190]), .Z(n8468) );
  AND U12702 ( .A(p_input[6190]), .B(p_input[36190]), .Z(n8467) );
  AND U12703 ( .A(n8469), .B(n8470), .Z(o[618]) );
  AND U12704 ( .A(p_input[20618]), .B(p_input[10618]), .Z(n8470) );
  AND U12705 ( .A(p_input[618]), .B(p_input[30618]), .Z(n8469) );
  AND U12706 ( .A(n8471), .B(n8472), .Z(o[6189]) );
  AND U12707 ( .A(p_input[26189]), .B(p_input[16189]), .Z(n8472) );
  AND U12708 ( .A(p_input[6189]), .B(p_input[36189]), .Z(n8471) );
  AND U12709 ( .A(n8473), .B(n8474), .Z(o[6188]) );
  AND U12710 ( .A(p_input[26188]), .B(p_input[16188]), .Z(n8474) );
  AND U12711 ( .A(p_input[6188]), .B(p_input[36188]), .Z(n8473) );
  AND U12712 ( .A(n8475), .B(n8476), .Z(o[6187]) );
  AND U12713 ( .A(p_input[26187]), .B(p_input[16187]), .Z(n8476) );
  AND U12714 ( .A(p_input[6187]), .B(p_input[36187]), .Z(n8475) );
  AND U12715 ( .A(n8477), .B(n8478), .Z(o[6186]) );
  AND U12716 ( .A(p_input[26186]), .B(p_input[16186]), .Z(n8478) );
  AND U12717 ( .A(p_input[6186]), .B(p_input[36186]), .Z(n8477) );
  AND U12718 ( .A(n8479), .B(n8480), .Z(o[6185]) );
  AND U12719 ( .A(p_input[26185]), .B(p_input[16185]), .Z(n8480) );
  AND U12720 ( .A(p_input[6185]), .B(p_input[36185]), .Z(n8479) );
  AND U12721 ( .A(n8481), .B(n8482), .Z(o[6184]) );
  AND U12722 ( .A(p_input[26184]), .B(p_input[16184]), .Z(n8482) );
  AND U12723 ( .A(p_input[6184]), .B(p_input[36184]), .Z(n8481) );
  AND U12724 ( .A(n8483), .B(n8484), .Z(o[6183]) );
  AND U12725 ( .A(p_input[26183]), .B(p_input[16183]), .Z(n8484) );
  AND U12726 ( .A(p_input[6183]), .B(p_input[36183]), .Z(n8483) );
  AND U12727 ( .A(n8485), .B(n8486), .Z(o[6182]) );
  AND U12728 ( .A(p_input[26182]), .B(p_input[16182]), .Z(n8486) );
  AND U12729 ( .A(p_input[6182]), .B(p_input[36182]), .Z(n8485) );
  AND U12730 ( .A(n8487), .B(n8488), .Z(o[6181]) );
  AND U12731 ( .A(p_input[26181]), .B(p_input[16181]), .Z(n8488) );
  AND U12732 ( .A(p_input[6181]), .B(p_input[36181]), .Z(n8487) );
  AND U12733 ( .A(n8489), .B(n8490), .Z(o[6180]) );
  AND U12734 ( .A(p_input[26180]), .B(p_input[16180]), .Z(n8490) );
  AND U12735 ( .A(p_input[6180]), .B(p_input[36180]), .Z(n8489) );
  AND U12736 ( .A(n8491), .B(n8492), .Z(o[617]) );
  AND U12737 ( .A(p_input[20617]), .B(p_input[10617]), .Z(n8492) );
  AND U12738 ( .A(p_input[617]), .B(p_input[30617]), .Z(n8491) );
  AND U12739 ( .A(n8493), .B(n8494), .Z(o[6179]) );
  AND U12740 ( .A(p_input[26179]), .B(p_input[16179]), .Z(n8494) );
  AND U12741 ( .A(p_input[6179]), .B(p_input[36179]), .Z(n8493) );
  AND U12742 ( .A(n8495), .B(n8496), .Z(o[6178]) );
  AND U12743 ( .A(p_input[26178]), .B(p_input[16178]), .Z(n8496) );
  AND U12744 ( .A(p_input[6178]), .B(p_input[36178]), .Z(n8495) );
  AND U12745 ( .A(n8497), .B(n8498), .Z(o[6177]) );
  AND U12746 ( .A(p_input[26177]), .B(p_input[16177]), .Z(n8498) );
  AND U12747 ( .A(p_input[6177]), .B(p_input[36177]), .Z(n8497) );
  AND U12748 ( .A(n8499), .B(n8500), .Z(o[6176]) );
  AND U12749 ( .A(p_input[26176]), .B(p_input[16176]), .Z(n8500) );
  AND U12750 ( .A(p_input[6176]), .B(p_input[36176]), .Z(n8499) );
  AND U12751 ( .A(n8501), .B(n8502), .Z(o[6175]) );
  AND U12752 ( .A(p_input[26175]), .B(p_input[16175]), .Z(n8502) );
  AND U12753 ( .A(p_input[6175]), .B(p_input[36175]), .Z(n8501) );
  AND U12754 ( .A(n8503), .B(n8504), .Z(o[6174]) );
  AND U12755 ( .A(p_input[26174]), .B(p_input[16174]), .Z(n8504) );
  AND U12756 ( .A(p_input[6174]), .B(p_input[36174]), .Z(n8503) );
  AND U12757 ( .A(n8505), .B(n8506), .Z(o[6173]) );
  AND U12758 ( .A(p_input[26173]), .B(p_input[16173]), .Z(n8506) );
  AND U12759 ( .A(p_input[6173]), .B(p_input[36173]), .Z(n8505) );
  AND U12760 ( .A(n8507), .B(n8508), .Z(o[6172]) );
  AND U12761 ( .A(p_input[26172]), .B(p_input[16172]), .Z(n8508) );
  AND U12762 ( .A(p_input[6172]), .B(p_input[36172]), .Z(n8507) );
  AND U12763 ( .A(n8509), .B(n8510), .Z(o[6171]) );
  AND U12764 ( .A(p_input[26171]), .B(p_input[16171]), .Z(n8510) );
  AND U12765 ( .A(p_input[6171]), .B(p_input[36171]), .Z(n8509) );
  AND U12766 ( .A(n8511), .B(n8512), .Z(o[6170]) );
  AND U12767 ( .A(p_input[26170]), .B(p_input[16170]), .Z(n8512) );
  AND U12768 ( .A(p_input[6170]), .B(p_input[36170]), .Z(n8511) );
  AND U12769 ( .A(n8513), .B(n8514), .Z(o[616]) );
  AND U12770 ( .A(p_input[20616]), .B(p_input[10616]), .Z(n8514) );
  AND U12771 ( .A(p_input[616]), .B(p_input[30616]), .Z(n8513) );
  AND U12772 ( .A(n8515), .B(n8516), .Z(o[6169]) );
  AND U12773 ( .A(p_input[26169]), .B(p_input[16169]), .Z(n8516) );
  AND U12774 ( .A(p_input[6169]), .B(p_input[36169]), .Z(n8515) );
  AND U12775 ( .A(n8517), .B(n8518), .Z(o[6168]) );
  AND U12776 ( .A(p_input[26168]), .B(p_input[16168]), .Z(n8518) );
  AND U12777 ( .A(p_input[6168]), .B(p_input[36168]), .Z(n8517) );
  AND U12778 ( .A(n8519), .B(n8520), .Z(o[6167]) );
  AND U12779 ( .A(p_input[26167]), .B(p_input[16167]), .Z(n8520) );
  AND U12780 ( .A(p_input[6167]), .B(p_input[36167]), .Z(n8519) );
  AND U12781 ( .A(n8521), .B(n8522), .Z(o[6166]) );
  AND U12782 ( .A(p_input[26166]), .B(p_input[16166]), .Z(n8522) );
  AND U12783 ( .A(p_input[6166]), .B(p_input[36166]), .Z(n8521) );
  AND U12784 ( .A(n8523), .B(n8524), .Z(o[6165]) );
  AND U12785 ( .A(p_input[26165]), .B(p_input[16165]), .Z(n8524) );
  AND U12786 ( .A(p_input[6165]), .B(p_input[36165]), .Z(n8523) );
  AND U12787 ( .A(n8525), .B(n8526), .Z(o[6164]) );
  AND U12788 ( .A(p_input[26164]), .B(p_input[16164]), .Z(n8526) );
  AND U12789 ( .A(p_input[6164]), .B(p_input[36164]), .Z(n8525) );
  AND U12790 ( .A(n8527), .B(n8528), .Z(o[6163]) );
  AND U12791 ( .A(p_input[26163]), .B(p_input[16163]), .Z(n8528) );
  AND U12792 ( .A(p_input[6163]), .B(p_input[36163]), .Z(n8527) );
  AND U12793 ( .A(n8529), .B(n8530), .Z(o[6162]) );
  AND U12794 ( .A(p_input[26162]), .B(p_input[16162]), .Z(n8530) );
  AND U12795 ( .A(p_input[6162]), .B(p_input[36162]), .Z(n8529) );
  AND U12796 ( .A(n8531), .B(n8532), .Z(o[6161]) );
  AND U12797 ( .A(p_input[26161]), .B(p_input[16161]), .Z(n8532) );
  AND U12798 ( .A(p_input[6161]), .B(p_input[36161]), .Z(n8531) );
  AND U12799 ( .A(n8533), .B(n8534), .Z(o[6160]) );
  AND U12800 ( .A(p_input[26160]), .B(p_input[16160]), .Z(n8534) );
  AND U12801 ( .A(p_input[6160]), .B(p_input[36160]), .Z(n8533) );
  AND U12802 ( .A(n8535), .B(n8536), .Z(o[615]) );
  AND U12803 ( .A(p_input[20615]), .B(p_input[10615]), .Z(n8536) );
  AND U12804 ( .A(p_input[615]), .B(p_input[30615]), .Z(n8535) );
  AND U12805 ( .A(n8537), .B(n8538), .Z(o[6159]) );
  AND U12806 ( .A(p_input[26159]), .B(p_input[16159]), .Z(n8538) );
  AND U12807 ( .A(p_input[6159]), .B(p_input[36159]), .Z(n8537) );
  AND U12808 ( .A(n8539), .B(n8540), .Z(o[6158]) );
  AND U12809 ( .A(p_input[26158]), .B(p_input[16158]), .Z(n8540) );
  AND U12810 ( .A(p_input[6158]), .B(p_input[36158]), .Z(n8539) );
  AND U12811 ( .A(n8541), .B(n8542), .Z(o[6157]) );
  AND U12812 ( .A(p_input[26157]), .B(p_input[16157]), .Z(n8542) );
  AND U12813 ( .A(p_input[6157]), .B(p_input[36157]), .Z(n8541) );
  AND U12814 ( .A(n8543), .B(n8544), .Z(o[6156]) );
  AND U12815 ( .A(p_input[26156]), .B(p_input[16156]), .Z(n8544) );
  AND U12816 ( .A(p_input[6156]), .B(p_input[36156]), .Z(n8543) );
  AND U12817 ( .A(n8545), .B(n8546), .Z(o[6155]) );
  AND U12818 ( .A(p_input[26155]), .B(p_input[16155]), .Z(n8546) );
  AND U12819 ( .A(p_input[6155]), .B(p_input[36155]), .Z(n8545) );
  AND U12820 ( .A(n8547), .B(n8548), .Z(o[6154]) );
  AND U12821 ( .A(p_input[26154]), .B(p_input[16154]), .Z(n8548) );
  AND U12822 ( .A(p_input[6154]), .B(p_input[36154]), .Z(n8547) );
  AND U12823 ( .A(n8549), .B(n8550), .Z(o[6153]) );
  AND U12824 ( .A(p_input[26153]), .B(p_input[16153]), .Z(n8550) );
  AND U12825 ( .A(p_input[6153]), .B(p_input[36153]), .Z(n8549) );
  AND U12826 ( .A(n8551), .B(n8552), .Z(o[6152]) );
  AND U12827 ( .A(p_input[26152]), .B(p_input[16152]), .Z(n8552) );
  AND U12828 ( .A(p_input[6152]), .B(p_input[36152]), .Z(n8551) );
  AND U12829 ( .A(n8553), .B(n8554), .Z(o[6151]) );
  AND U12830 ( .A(p_input[26151]), .B(p_input[16151]), .Z(n8554) );
  AND U12831 ( .A(p_input[6151]), .B(p_input[36151]), .Z(n8553) );
  AND U12832 ( .A(n8555), .B(n8556), .Z(o[6150]) );
  AND U12833 ( .A(p_input[26150]), .B(p_input[16150]), .Z(n8556) );
  AND U12834 ( .A(p_input[6150]), .B(p_input[36150]), .Z(n8555) );
  AND U12835 ( .A(n8557), .B(n8558), .Z(o[614]) );
  AND U12836 ( .A(p_input[20614]), .B(p_input[10614]), .Z(n8558) );
  AND U12837 ( .A(p_input[614]), .B(p_input[30614]), .Z(n8557) );
  AND U12838 ( .A(n8559), .B(n8560), .Z(o[6149]) );
  AND U12839 ( .A(p_input[26149]), .B(p_input[16149]), .Z(n8560) );
  AND U12840 ( .A(p_input[6149]), .B(p_input[36149]), .Z(n8559) );
  AND U12841 ( .A(n8561), .B(n8562), .Z(o[6148]) );
  AND U12842 ( .A(p_input[26148]), .B(p_input[16148]), .Z(n8562) );
  AND U12843 ( .A(p_input[6148]), .B(p_input[36148]), .Z(n8561) );
  AND U12844 ( .A(n8563), .B(n8564), .Z(o[6147]) );
  AND U12845 ( .A(p_input[26147]), .B(p_input[16147]), .Z(n8564) );
  AND U12846 ( .A(p_input[6147]), .B(p_input[36147]), .Z(n8563) );
  AND U12847 ( .A(n8565), .B(n8566), .Z(o[6146]) );
  AND U12848 ( .A(p_input[26146]), .B(p_input[16146]), .Z(n8566) );
  AND U12849 ( .A(p_input[6146]), .B(p_input[36146]), .Z(n8565) );
  AND U12850 ( .A(n8567), .B(n8568), .Z(o[6145]) );
  AND U12851 ( .A(p_input[26145]), .B(p_input[16145]), .Z(n8568) );
  AND U12852 ( .A(p_input[6145]), .B(p_input[36145]), .Z(n8567) );
  AND U12853 ( .A(n8569), .B(n8570), .Z(o[6144]) );
  AND U12854 ( .A(p_input[26144]), .B(p_input[16144]), .Z(n8570) );
  AND U12855 ( .A(p_input[6144]), .B(p_input[36144]), .Z(n8569) );
  AND U12856 ( .A(n8571), .B(n8572), .Z(o[6143]) );
  AND U12857 ( .A(p_input[26143]), .B(p_input[16143]), .Z(n8572) );
  AND U12858 ( .A(p_input[6143]), .B(p_input[36143]), .Z(n8571) );
  AND U12859 ( .A(n8573), .B(n8574), .Z(o[6142]) );
  AND U12860 ( .A(p_input[26142]), .B(p_input[16142]), .Z(n8574) );
  AND U12861 ( .A(p_input[6142]), .B(p_input[36142]), .Z(n8573) );
  AND U12862 ( .A(n8575), .B(n8576), .Z(o[6141]) );
  AND U12863 ( .A(p_input[26141]), .B(p_input[16141]), .Z(n8576) );
  AND U12864 ( .A(p_input[6141]), .B(p_input[36141]), .Z(n8575) );
  AND U12865 ( .A(n8577), .B(n8578), .Z(o[6140]) );
  AND U12866 ( .A(p_input[26140]), .B(p_input[16140]), .Z(n8578) );
  AND U12867 ( .A(p_input[6140]), .B(p_input[36140]), .Z(n8577) );
  AND U12868 ( .A(n8579), .B(n8580), .Z(o[613]) );
  AND U12869 ( .A(p_input[20613]), .B(p_input[10613]), .Z(n8580) );
  AND U12870 ( .A(p_input[613]), .B(p_input[30613]), .Z(n8579) );
  AND U12871 ( .A(n8581), .B(n8582), .Z(o[6139]) );
  AND U12872 ( .A(p_input[26139]), .B(p_input[16139]), .Z(n8582) );
  AND U12873 ( .A(p_input[6139]), .B(p_input[36139]), .Z(n8581) );
  AND U12874 ( .A(n8583), .B(n8584), .Z(o[6138]) );
  AND U12875 ( .A(p_input[26138]), .B(p_input[16138]), .Z(n8584) );
  AND U12876 ( .A(p_input[6138]), .B(p_input[36138]), .Z(n8583) );
  AND U12877 ( .A(n8585), .B(n8586), .Z(o[6137]) );
  AND U12878 ( .A(p_input[26137]), .B(p_input[16137]), .Z(n8586) );
  AND U12879 ( .A(p_input[6137]), .B(p_input[36137]), .Z(n8585) );
  AND U12880 ( .A(n8587), .B(n8588), .Z(o[6136]) );
  AND U12881 ( .A(p_input[26136]), .B(p_input[16136]), .Z(n8588) );
  AND U12882 ( .A(p_input[6136]), .B(p_input[36136]), .Z(n8587) );
  AND U12883 ( .A(n8589), .B(n8590), .Z(o[6135]) );
  AND U12884 ( .A(p_input[26135]), .B(p_input[16135]), .Z(n8590) );
  AND U12885 ( .A(p_input[6135]), .B(p_input[36135]), .Z(n8589) );
  AND U12886 ( .A(n8591), .B(n8592), .Z(o[6134]) );
  AND U12887 ( .A(p_input[26134]), .B(p_input[16134]), .Z(n8592) );
  AND U12888 ( .A(p_input[6134]), .B(p_input[36134]), .Z(n8591) );
  AND U12889 ( .A(n8593), .B(n8594), .Z(o[6133]) );
  AND U12890 ( .A(p_input[26133]), .B(p_input[16133]), .Z(n8594) );
  AND U12891 ( .A(p_input[6133]), .B(p_input[36133]), .Z(n8593) );
  AND U12892 ( .A(n8595), .B(n8596), .Z(o[6132]) );
  AND U12893 ( .A(p_input[26132]), .B(p_input[16132]), .Z(n8596) );
  AND U12894 ( .A(p_input[6132]), .B(p_input[36132]), .Z(n8595) );
  AND U12895 ( .A(n8597), .B(n8598), .Z(o[6131]) );
  AND U12896 ( .A(p_input[26131]), .B(p_input[16131]), .Z(n8598) );
  AND U12897 ( .A(p_input[6131]), .B(p_input[36131]), .Z(n8597) );
  AND U12898 ( .A(n8599), .B(n8600), .Z(o[6130]) );
  AND U12899 ( .A(p_input[26130]), .B(p_input[16130]), .Z(n8600) );
  AND U12900 ( .A(p_input[6130]), .B(p_input[36130]), .Z(n8599) );
  AND U12901 ( .A(n8601), .B(n8602), .Z(o[612]) );
  AND U12902 ( .A(p_input[20612]), .B(p_input[10612]), .Z(n8602) );
  AND U12903 ( .A(p_input[612]), .B(p_input[30612]), .Z(n8601) );
  AND U12904 ( .A(n8603), .B(n8604), .Z(o[6129]) );
  AND U12905 ( .A(p_input[26129]), .B(p_input[16129]), .Z(n8604) );
  AND U12906 ( .A(p_input[6129]), .B(p_input[36129]), .Z(n8603) );
  AND U12907 ( .A(n8605), .B(n8606), .Z(o[6128]) );
  AND U12908 ( .A(p_input[26128]), .B(p_input[16128]), .Z(n8606) );
  AND U12909 ( .A(p_input[6128]), .B(p_input[36128]), .Z(n8605) );
  AND U12910 ( .A(n8607), .B(n8608), .Z(o[6127]) );
  AND U12911 ( .A(p_input[26127]), .B(p_input[16127]), .Z(n8608) );
  AND U12912 ( .A(p_input[6127]), .B(p_input[36127]), .Z(n8607) );
  AND U12913 ( .A(n8609), .B(n8610), .Z(o[6126]) );
  AND U12914 ( .A(p_input[26126]), .B(p_input[16126]), .Z(n8610) );
  AND U12915 ( .A(p_input[6126]), .B(p_input[36126]), .Z(n8609) );
  AND U12916 ( .A(n8611), .B(n8612), .Z(o[6125]) );
  AND U12917 ( .A(p_input[26125]), .B(p_input[16125]), .Z(n8612) );
  AND U12918 ( .A(p_input[6125]), .B(p_input[36125]), .Z(n8611) );
  AND U12919 ( .A(n8613), .B(n8614), .Z(o[6124]) );
  AND U12920 ( .A(p_input[26124]), .B(p_input[16124]), .Z(n8614) );
  AND U12921 ( .A(p_input[6124]), .B(p_input[36124]), .Z(n8613) );
  AND U12922 ( .A(n8615), .B(n8616), .Z(o[6123]) );
  AND U12923 ( .A(p_input[26123]), .B(p_input[16123]), .Z(n8616) );
  AND U12924 ( .A(p_input[6123]), .B(p_input[36123]), .Z(n8615) );
  AND U12925 ( .A(n8617), .B(n8618), .Z(o[6122]) );
  AND U12926 ( .A(p_input[26122]), .B(p_input[16122]), .Z(n8618) );
  AND U12927 ( .A(p_input[6122]), .B(p_input[36122]), .Z(n8617) );
  AND U12928 ( .A(n8619), .B(n8620), .Z(o[6121]) );
  AND U12929 ( .A(p_input[26121]), .B(p_input[16121]), .Z(n8620) );
  AND U12930 ( .A(p_input[6121]), .B(p_input[36121]), .Z(n8619) );
  AND U12931 ( .A(n8621), .B(n8622), .Z(o[6120]) );
  AND U12932 ( .A(p_input[26120]), .B(p_input[16120]), .Z(n8622) );
  AND U12933 ( .A(p_input[6120]), .B(p_input[36120]), .Z(n8621) );
  AND U12934 ( .A(n8623), .B(n8624), .Z(o[611]) );
  AND U12935 ( .A(p_input[20611]), .B(p_input[10611]), .Z(n8624) );
  AND U12936 ( .A(p_input[611]), .B(p_input[30611]), .Z(n8623) );
  AND U12937 ( .A(n8625), .B(n8626), .Z(o[6119]) );
  AND U12938 ( .A(p_input[26119]), .B(p_input[16119]), .Z(n8626) );
  AND U12939 ( .A(p_input[6119]), .B(p_input[36119]), .Z(n8625) );
  AND U12940 ( .A(n8627), .B(n8628), .Z(o[6118]) );
  AND U12941 ( .A(p_input[26118]), .B(p_input[16118]), .Z(n8628) );
  AND U12942 ( .A(p_input[6118]), .B(p_input[36118]), .Z(n8627) );
  AND U12943 ( .A(n8629), .B(n8630), .Z(o[6117]) );
  AND U12944 ( .A(p_input[26117]), .B(p_input[16117]), .Z(n8630) );
  AND U12945 ( .A(p_input[6117]), .B(p_input[36117]), .Z(n8629) );
  AND U12946 ( .A(n8631), .B(n8632), .Z(o[6116]) );
  AND U12947 ( .A(p_input[26116]), .B(p_input[16116]), .Z(n8632) );
  AND U12948 ( .A(p_input[6116]), .B(p_input[36116]), .Z(n8631) );
  AND U12949 ( .A(n8633), .B(n8634), .Z(o[6115]) );
  AND U12950 ( .A(p_input[26115]), .B(p_input[16115]), .Z(n8634) );
  AND U12951 ( .A(p_input[6115]), .B(p_input[36115]), .Z(n8633) );
  AND U12952 ( .A(n8635), .B(n8636), .Z(o[6114]) );
  AND U12953 ( .A(p_input[26114]), .B(p_input[16114]), .Z(n8636) );
  AND U12954 ( .A(p_input[6114]), .B(p_input[36114]), .Z(n8635) );
  AND U12955 ( .A(n8637), .B(n8638), .Z(o[6113]) );
  AND U12956 ( .A(p_input[26113]), .B(p_input[16113]), .Z(n8638) );
  AND U12957 ( .A(p_input[6113]), .B(p_input[36113]), .Z(n8637) );
  AND U12958 ( .A(n8639), .B(n8640), .Z(o[6112]) );
  AND U12959 ( .A(p_input[26112]), .B(p_input[16112]), .Z(n8640) );
  AND U12960 ( .A(p_input[6112]), .B(p_input[36112]), .Z(n8639) );
  AND U12961 ( .A(n8641), .B(n8642), .Z(o[6111]) );
  AND U12962 ( .A(p_input[26111]), .B(p_input[16111]), .Z(n8642) );
  AND U12963 ( .A(p_input[6111]), .B(p_input[36111]), .Z(n8641) );
  AND U12964 ( .A(n8643), .B(n8644), .Z(o[6110]) );
  AND U12965 ( .A(p_input[26110]), .B(p_input[16110]), .Z(n8644) );
  AND U12966 ( .A(p_input[6110]), .B(p_input[36110]), .Z(n8643) );
  AND U12967 ( .A(n8645), .B(n8646), .Z(o[610]) );
  AND U12968 ( .A(p_input[20610]), .B(p_input[10610]), .Z(n8646) );
  AND U12969 ( .A(p_input[610]), .B(p_input[30610]), .Z(n8645) );
  AND U12970 ( .A(n8647), .B(n8648), .Z(o[6109]) );
  AND U12971 ( .A(p_input[26109]), .B(p_input[16109]), .Z(n8648) );
  AND U12972 ( .A(p_input[6109]), .B(p_input[36109]), .Z(n8647) );
  AND U12973 ( .A(n8649), .B(n8650), .Z(o[6108]) );
  AND U12974 ( .A(p_input[26108]), .B(p_input[16108]), .Z(n8650) );
  AND U12975 ( .A(p_input[6108]), .B(p_input[36108]), .Z(n8649) );
  AND U12976 ( .A(n8651), .B(n8652), .Z(o[6107]) );
  AND U12977 ( .A(p_input[26107]), .B(p_input[16107]), .Z(n8652) );
  AND U12978 ( .A(p_input[6107]), .B(p_input[36107]), .Z(n8651) );
  AND U12979 ( .A(n8653), .B(n8654), .Z(o[6106]) );
  AND U12980 ( .A(p_input[26106]), .B(p_input[16106]), .Z(n8654) );
  AND U12981 ( .A(p_input[6106]), .B(p_input[36106]), .Z(n8653) );
  AND U12982 ( .A(n8655), .B(n8656), .Z(o[6105]) );
  AND U12983 ( .A(p_input[26105]), .B(p_input[16105]), .Z(n8656) );
  AND U12984 ( .A(p_input[6105]), .B(p_input[36105]), .Z(n8655) );
  AND U12985 ( .A(n8657), .B(n8658), .Z(o[6104]) );
  AND U12986 ( .A(p_input[26104]), .B(p_input[16104]), .Z(n8658) );
  AND U12987 ( .A(p_input[6104]), .B(p_input[36104]), .Z(n8657) );
  AND U12988 ( .A(n8659), .B(n8660), .Z(o[6103]) );
  AND U12989 ( .A(p_input[26103]), .B(p_input[16103]), .Z(n8660) );
  AND U12990 ( .A(p_input[6103]), .B(p_input[36103]), .Z(n8659) );
  AND U12991 ( .A(n8661), .B(n8662), .Z(o[6102]) );
  AND U12992 ( .A(p_input[26102]), .B(p_input[16102]), .Z(n8662) );
  AND U12993 ( .A(p_input[6102]), .B(p_input[36102]), .Z(n8661) );
  AND U12994 ( .A(n8663), .B(n8664), .Z(o[6101]) );
  AND U12995 ( .A(p_input[26101]), .B(p_input[16101]), .Z(n8664) );
  AND U12996 ( .A(p_input[6101]), .B(p_input[36101]), .Z(n8663) );
  AND U12997 ( .A(n8665), .B(n8666), .Z(o[6100]) );
  AND U12998 ( .A(p_input[26100]), .B(p_input[16100]), .Z(n8666) );
  AND U12999 ( .A(p_input[6100]), .B(p_input[36100]), .Z(n8665) );
  AND U13000 ( .A(n8667), .B(n8668), .Z(o[60]) );
  AND U13001 ( .A(p_input[20060]), .B(p_input[10060]), .Z(n8668) );
  AND U13002 ( .A(p_input[60]), .B(p_input[30060]), .Z(n8667) );
  AND U13003 ( .A(n8669), .B(n8670), .Z(o[609]) );
  AND U13004 ( .A(p_input[20609]), .B(p_input[10609]), .Z(n8670) );
  AND U13005 ( .A(p_input[609]), .B(p_input[30609]), .Z(n8669) );
  AND U13006 ( .A(n8671), .B(n8672), .Z(o[6099]) );
  AND U13007 ( .A(p_input[26099]), .B(p_input[16099]), .Z(n8672) );
  AND U13008 ( .A(p_input[6099]), .B(p_input[36099]), .Z(n8671) );
  AND U13009 ( .A(n8673), .B(n8674), .Z(o[6098]) );
  AND U13010 ( .A(p_input[26098]), .B(p_input[16098]), .Z(n8674) );
  AND U13011 ( .A(p_input[6098]), .B(p_input[36098]), .Z(n8673) );
  AND U13012 ( .A(n8675), .B(n8676), .Z(o[6097]) );
  AND U13013 ( .A(p_input[26097]), .B(p_input[16097]), .Z(n8676) );
  AND U13014 ( .A(p_input[6097]), .B(p_input[36097]), .Z(n8675) );
  AND U13015 ( .A(n8677), .B(n8678), .Z(o[6096]) );
  AND U13016 ( .A(p_input[26096]), .B(p_input[16096]), .Z(n8678) );
  AND U13017 ( .A(p_input[6096]), .B(p_input[36096]), .Z(n8677) );
  AND U13018 ( .A(n8679), .B(n8680), .Z(o[6095]) );
  AND U13019 ( .A(p_input[26095]), .B(p_input[16095]), .Z(n8680) );
  AND U13020 ( .A(p_input[6095]), .B(p_input[36095]), .Z(n8679) );
  AND U13021 ( .A(n8681), .B(n8682), .Z(o[6094]) );
  AND U13022 ( .A(p_input[26094]), .B(p_input[16094]), .Z(n8682) );
  AND U13023 ( .A(p_input[6094]), .B(p_input[36094]), .Z(n8681) );
  AND U13024 ( .A(n8683), .B(n8684), .Z(o[6093]) );
  AND U13025 ( .A(p_input[26093]), .B(p_input[16093]), .Z(n8684) );
  AND U13026 ( .A(p_input[6093]), .B(p_input[36093]), .Z(n8683) );
  AND U13027 ( .A(n8685), .B(n8686), .Z(o[6092]) );
  AND U13028 ( .A(p_input[26092]), .B(p_input[16092]), .Z(n8686) );
  AND U13029 ( .A(p_input[6092]), .B(p_input[36092]), .Z(n8685) );
  AND U13030 ( .A(n8687), .B(n8688), .Z(o[6091]) );
  AND U13031 ( .A(p_input[26091]), .B(p_input[16091]), .Z(n8688) );
  AND U13032 ( .A(p_input[6091]), .B(p_input[36091]), .Z(n8687) );
  AND U13033 ( .A(n8689), .B(n8690), .Z(o[6090]) );
  AND U13034 ( .A(p_input[26090]), .B(p_input[16090]), .Z(n8690) );
  AND U13035 ( .A(p_input[6090]), .B(p_input[36090]), .Z(n8689) );
  AND U13036 ( .A(n8691), .B(n8692), .Z(o[608]) );
  AND U13037 ( .A(p_input[20608]), .B(p_input[10608]), .Z(n8692) );
  AND U13038 ( .A(p_input[608]), .B(p_input[30608]), .Z(n8691) );
  AND U13039 ( .A(n8693), .B(n8694), .Z(o[6089]) );
  AND U13040 ( .A(p_input[26089]), .B(p_input[16089]), .Z(n8694) );
  AND U13041 ( .A(p_input[6089]), .B(p_input[36089]), .Z(n8693) );
  AND U13042 ( .A(n8695), .B(n8696), .Z(o[6088]) );
  AND U13043 ( .A(p_input[26088]), .B(p_input[16088]), .Z(n8696) );
  AND U13044 ( .A(p_input[6088]), .B(p_input[36088]), .Z(n8695) );
  AND U13045 ( .A(n8697), .B(n8698), .Z(o[6087]) );
  AND U13046 ( .A(p_input[26087]), .B(p_input[16087]), .Z(n8698) );
  AND U13047 ( .A(p_input[6087]), .B(p_input[36087]), .Z(n8697) );
  AND U13048 ( .A(n8699), .B(n8700), .Z(o[6086]) );
  AND U13049 ( .A(p_input[26086]), .B(p_input[16086]), .Z(n8700) );
  AND U13050 ( .A(p_input[6086]), .B(p_input[36086]), .Z(n8699) );
  AND U13051 ( .A(n8701), .B(n8702), .Z(o[6085]) );
  AND U13052 ( .A(p_input[26085]), .B(p_input[16085]), .Z(n8702) );
  AND U13053 ( .A(p_input[6085]), .B(p_input[36085]), .Z(n8701) );
  AND U13054 ( .A(n8703), .B(n8704), .Z(o[6084]) );
  AND U13055 ( .A(p_input[26084]), .B(p_input[16084]), .Z(n8704) );
  AND U13056 ( .A(p_input[6084]), .B(p_input[36084]), .Z(n8703) );
  AND U13057 ( .A(n8705), .B(n8706), .Z(o[6083]) );
  AND U13058 ( .A(p_input[26083]), .B(p_input[16083]), .Z(n8706) );
  AND U13059 ( .A(p_input[6083]), .B(p_input[36083]), .Z(n8705) );
  AND U13060 ( .A(n8707), .B(n8708), .Z(o[6082]) );
  AND U13061 ( .A(p_input[26082]), .B(p_input[16082]), .Z(n8708) );
  AND U13062 ( .A(p_input[6082]), .B(p_input[36082]), .Z(n8707) );
  AND U13063 ( .A(n8709), .B(n8710), .Z(o[6081]) );
  AND U13064 ( .A(p_input[26081]), .B(p_input[16081]), .Z(n8710) );
  AND U13065 ( .A(p_input[6081]), .B(p_input[36081]), .Z(n8709) );
  AND U13066 ( .A(n8711), .B(n8712), .Z(o[6080]) );
  AND U13067 ( .A(p_input[26080]), .B(p_input[16080]), .Z(n8712) );
  AND U13068 ( .A(p_input[6080]), .B(p_input[36080]), .Z(n8711) );
  AND U13069 ( .A(n8713), .B(n8714), .Z(o[607]) );
  AND U13070 ( .A(p_input[20607]), .B(p_input[10607]), .Z(n8714) );
  AND U13071 ( .A(p_input[607]), .B(p_input[30607]), .Z(n8713) );
  AND U13072 ( .A(n8715), .B(n8716), .Z(o[6079]) );
  AND U13073 ( .A(p_input[26079]), .B(p_input[16079]), .Z(n8716) );
  AND U13074 ( .A(p_input[6079]), .B(p_input[36079]), .Z(n8715) );
  AND U13075 ( .A(n8717), .B(n8718), .Z(o[6078]) );
  AND U13076 ( .A(p_input[26078]), .B(p_input[16078]), .Z(n8718) );
  AND U13077 ( .A(p_input[6078]), .B(p_input[36078]), .Z(n8717) );
  AND U13078 ( .A(n8719), .B(n8720), .Z(o[6077]) );
  AND U13079 ( .A(p_input[26077]), .B(p_input[16077]), .Z(n8720) );
  AND U13080 ( .A(p_input[6077]), .B(p_input[36077]), .Z(n8719) );
  AND U13081 ( .A(n8721), .B(n8722), .Z(o[6076]) );
  AND U13082 ( .A(p_input[26076]), .B(p_input[16076]), .Z(n8722) );
  AND U13083 ( .A(p_input[6076]), .B(p_input[36076]), .Z(n8721) );
  AND U13084 ( .A(n8723), .B(n8724), .Z(o[6075]) );
  AND U13085 ( .A(p_input[26075]), .B(p_input[16075]), .Z(n8724) );
  AND U13086 ( .A(p_input[6075]), .B(p_input[36075]), .Z(n8723) );
  AND U13087 ( .A(n8725), .B(n8726), .Z(o[6074]) );
  AND U13088 ( .A(p_input[26074]), .B(p_input[16074]), .Z(n8726) );
  AND U13089 ( .A(p_input[6074]), .B(p_input[36074]), .Z(n8725) );
  AND U13090 ( .A(n8727), .B(n8728), .Z(o[6073]) );
  AND U13091 ( .A(p_input[26073]), .B(p_input[16073]), .Z(n8728) );
  AND U13092 ( .A(p_input[6073]), .B(p_input[36073]), .Z(n8727) );
  AND U13093 ( .A(n8729), .B(n8730), .Z(o[6072]) );
  AND U13094 ( .A(p_input[26072]), .B(p_input[16072]), .Z(n8730) );
  AND U13095 ( .A(p_input[6072]), .B(p_input[36072]), .Z(n8729) );
  AND U13096 ( .A(n8731), .B(n8732), .Z(o[6071]) );
  AND U13097 ( .A(p_input[26071]), .B(p_input[16071]), .Z(n8732) );
  AND U13098 ( .A(p_input[6071]), .B(p_input[36071]), .Z(n8731) );
  AND U13099 ( .A(n8733), .B(n8734), .Z(o[6070]) );
  AND U13100 ( .A(p_input[26070]), .B(p_input[16070]), .Z(n8734) );
  AND U13101 ( .A(p_input[6070]), .B(p_input[36070]), .Z(n8733) );
  AND U13102 ( .A(n8735), .B(n8736), .Z(o[606]) );
  AND U13103 ( .A(p_input[20606]), .B(p_input[10606]), .Z(n8736) );
  AND U13104 ( .A(p_input[606]), .B(p_input[30606]), .Z(n8735) );
  AND U13105 ( .A(n8737), .B(n8738), .Z(o[6069]) );
  AND U13106 ( .A(p_input[26069]), .B(p_input[16069]), .Z(n8738) );
  AND U13107 ( .A(p_input[6069]), .B(p_input[36069]), .Z(n8737) );
  AND U13108 ( .A(n8739), .B(n8740), .Z(o[6068]) );
  AND U13109 ( .A(p_input[26068]), .B(p_input[16068]), .Z(n8740) );
  AND U13110 ( .A(p_input[6068]), .B(p_input[36068]), .Z(n8739) );
  AND U13111 ( .A(n8741), .B(n8742), .Z(o[6067]) );
  AND U13112 ( .A(p_input[26067]), .B(p_input[16067]), .Z(n8742) );
  AND U13113 ( .A(p_input[6067]), .B(p_input[36067]), .Z(n8741) );
  AND U13114 ( .A(n8743), .B(n8744), .Z(o[6066]) );
  AND U13115 ( .A(p_input[26066]), .B(p_input[16066]), .Z(n8744) );
  AND U13116 ( .A(p_input[6066]), .B(p_input[36066]), .Z(n8743) );
  AND U13117 ( .A(n8745), .B(n8746), .Z(o[6065]) );
  AND U13118 ( .A(p_input[26065]), .B(p_input[16065]), .Z(n8746) );
  AND U13119 ( .A(p_input[6065]), .B(p_input[36065]), .Z(n8745) );
  AND U13120 ( .A(n8747), .B(n8748), .Z(o[6064]) );
  AND U13121 ( .A(p_input[26064]), .B(p_input[16064]), .Z(n8748) );
  AND U13122 ( .A(p_input[6064]), .B(p_input[36064]), .Z(n8747) );
  AND U13123 ( .A(n8749), .B(n8750), .Z(o[6063]) );
  AND U13124 ( .A(p_input[26063]), .B(p_input[16063]), .Z(n8750) );
  AND U13125 ( .A(p_input[6063]), .B(p_input[36063]), .Z(n8749) );
  AND U13126 ( .A(n8751), .B(n8752), .Z(o[6062]) );
  AND U13127 ( .A(p_input[26062]), .B(p_input[16062]), .Z(n8752) );
  AND U13128 ( .A(p_input[6062]), .B(p_input[36062]), .Z(n8751) );
  AND U13129 ( .A(n8753), .B(n8754), .Z(o[6061]) );
  AND U13130 ( .A(p_input[26061]), .B(p_input[16061]), .Z(n8754) );
  AND U13131 ( .A(p_input[6061]), .B(p_input[36061]), .Z(n8753) );
  AND U13132 ( .A(n8755), .B(n8756), .Z(o[6060]) );
  AND U13133 ( .A(p_input[26060]), .B(p_input[16060]), .Z(n8756) );
  AND U13134 ( .A(p_input[6060]), .B(p_input[36060]), .Z(n8755) );
  AND U13135 ( .A(n8757), .B(n8758), .Z(o[605]) );
  AND U13136 ( .A(p_input[20605]), .B(p_input[10605]), .Z(n8758) );
  AND U13137 ( .A(p_input[605]), .B(p_input[30605]), .Z(n8757) );
  AND U13138 ( .A(n8759), .B(n8760), .Z(o[6059]) );
  AND U13139 ( .A(p_input[26059]), .B(p_input[16059]), .Z(n8760) );
  AND U13140 ( .A(p_input[6059]), .B(p_input[36059]), .Z(n8759) );
  AND U13141 ( .A(n8761), .B(n8762), .Z(o[6058]) );
  AND U13142 ( .A(p_input[26058]), .B(p_input[16058]), .Z(n8762) );
  AND U13143 ( .A(p_input[6058]), .B(p_input[36058]), .Z(n8761) );
  AND U13144 ( .A(n8763), .B(n8764), .Z(o[6057]) );
  AND U13145 ( .A(p_input[26057]), .B(p_input[16057]), .Z(n8764) );
  AND U13146 ( .A(p_input[6057]), .B(p_input[36057]), .Z(n8763) );
  AND U13147 ( .A(n8765), .B(n8766), .Z(o[6056]) );
  AND U13148 ( .A(p_input[26056]), .B(p_input[16056]), .Z(n8766) );
  AND U13149 ( .A(p_input[6056]), .B(p_input[36056]), .Z(n8765) );
  AND U13150 ( .A(n8767), .B(n8768), .Z(o[6055]) );
  AND U13151 ( .A(p_input[26055]), .B(p_input[16055]), .Z(n8768) );
  AND U13152 ( .A(p_input[6055]), .B(p_input[36055]), .Z(n8767) );
  AND U13153 ( .A(n8769), .B(n8770), .Z(o[6054]) );
  AND U13154 ( .A(p_input[26054]), .B(p_input[16054]), .Z(n8770) );
  AND U13155 ( .A(p_input[6054]), .B(p_input[36054]), .Z(n8769) );
  AND U13156 ( .A(n8771), .B(n8772), .Z(o[6053]) );
  AND U13157 ( .A(p_input[26053]), .B(p_input[16053]), .Z(n8772) );
  AND U13158 ( .A(p_input[6053]), .B(p_input[36053]), .Z(n8771) );
  AND U13159 ( .A(n8773), .B(n8774), .Z(o[6052]) );
  AND U13160 ( .A(p_input[26052]), .B(p_input[16052]), .Z(n8774) );
  AND U13161 ( .A(p_input[6052]), .B(p_input[36052]), .Z(n8773) );
  AND U13162 ( .A(n8775), .B(n8776), .Z(o[6051]) );
  AND U13163 ( .A(p_input[26051]), .B(p_input[16051]), .Z(n8776) );
  AND U13164 ( .A(p_input[6051]), .B(p_input[36051]), .Z(n8775) );
  AND U13165 ( .A(n8777), .B(n8778), .Z(o[6050]) );
  AND U13166 ( .A(p_input[26050]), .B(p_input[16050]), .Z(n8778) );
  AND U13167 ( .A(p_input[6050]), .B(p_input[36050]), .Z(n8777) );
  AND U13168 ( .A(n8779), .B(n8780), .Z(o[604]) );
  AND U13169 ( .A(p_input[20604]), .B(p_input[10604]), .Z(n8780) );
  AND U13170 ( .A(p_input[604]), .B(p_input[30604]), .Z(n8779) );
  AND U13171 ( .A(n8781), .B(n8782), .Z(o[6049]) );
  AND U13172 ( .A(p_input[26049]), .B(p_input[16049]), .Z(n8782) );
  AND U13173 ( .A(p_input[6049]), .B(p_input[36049]), .Z(n8781) );
  AND U13174 ( .A(n8783), .B(n8784), .Z(o[6048]) );
  AND U13175 ( .A(p_input[26048]), .B(p_input[16048]), .Z(n8784) );
  AND U13176 ( .A(p_input[6048]), .B(p_input[36048]), .Z(n8783) );
  AND U13177 ( .A(n8785), .B(n8786), .Z(o[6047]) );
  AND U13178 ( .A(p_input[26047]), .B(p_input[16047]), .Z(n8786) );
  AND U13179 ( .A(p_input[6047]), .B(p_input[36047]), .Z(n8785) );
  AND U13180 ( .A(n8787), .B(n8788), .Z(o[6046]) );
  AND U13181 ( .A(p_input[26046]), .B(p_input[16046]), .Z(n8788) );
  AND U13182 ( .A(p_input[6046]), .B(p_input[36046]), .Z(n8787) );
  AND U13183 ( .A(n8789), .B(n8790), .Z(o[6045]) );
  AND U13184 ( .A(p_input[26045]), .B(p_input[16045]), .Z(n8790) );
  AND U13185 ( .A(p_input[6045]), .B(p_input[36045]), .Z(n8789) );
  AND U13186 ( .A(n8791), .B(n8792), .Z(o[6044]) );
  AND U13187 ( .A(p_input[26044]), .B(p_input[16044]), .Z(n8792) );
  AND U13188 ( .A(p_input[6044]), .B(p_input[36044]), .Z(n8791) );
  AND U13189 ( .A(n8793), .B(n8794), .Z(o[6043]) );
  AND U13190 ( .A(p_input[26043]), .B(p_input[16043]), .Z(n8794) );
  AND U13191 ( .A(p_input[6043]), .B(p_input[36043]), .Z(n8793) );
  AND U13192 ( .A(n8795), .B(n8796), .Z(o[6042]) );
  AND U13193 ( .A(p_input[26042]), .B(p_input[16042]), .Z(n8796) );
  AND U13194 ( .A(p_input[6042]), .B(p_input[36042]), .Z(n8795) );
  AND U13195 ( .A(n8797), .B(n8798), .Z(o[6041]) );
  AND U13196 ( .A(p_input[26041]), .B(p_input[16041]), .Z(n8798) );
  AND U13197 ( .A(p_input[6041]), .B(p_input[36041]), .Z(n8797) );
  AND U13198 ( .A(n8799), .B(n8800), .Z(o[6040]) );
  AND U13199 ( .A(p_input[26040]), .B(p_input[16040]), .Z(n8800) );
  AND U13200 ( .A(p_input[6040]), .B(p_input[36040]), .Z(n8799) );
  AND U13201 ( .A(n8801), .B(n8802), .Z(o[603]) );
  AND U13202 ( .A(p_input[20603]), .B(p_input[10603]), .Z(n8802) );
  AND U13203 ( .A(p_input[603]), .B(p_input[30603]), .Z(n8801) );
  AND U13204 ( .A(n8803), .B(n8804), .Z(o[6039]) );
  AND U13205 ( .A(p_input[26039]), .B(p_input[16039]), .Z(n8804) );
  AND U13206 ( .A(p_input[6039]), .B(p_input[36039]), .Z(n8803) );
  AND U13207 ( .A(n8805), .B(n8806), .Z(o[6038]) );
  AND U13208 ( .A(p_input[26038]), .B(p_input[16038]), .Z(n8806) );
  AND U13209 ( .A(p_input[6038]), .B(p_input[36038]), .Z(n8805) );
  AND U13210 ( .A(n8807), .B(n8808), .Z(o[6037]) );
  AND U13211 ( .A(p_input[26037]), .B(p_input[16037]), .Z(n8808) );
  AND U13212 ( .A(p_input[6037]), .B(p_input[36037]), .Z(n8807) );
  AND U13213 ( .A(n8809), .B(n8810), .Z(o[6036]) );
  AND U13214 ( .A(p_input[26036]), .B(p_input[16036]), .Z(n8810) );
  AND U13215 ( .A(p_input[6036]), .B(p_input[36036]), .Z(n8809) );
  AND U13216 ( .A(n8811), .B(n8812), .Z(o[6035]) );
  AND U13217 ( .A(p_input[26035]), .B(p_input[16035]), .Z(n8812) );
  AND U13218 ( .A(p_input[6035]), .B(p_input[36035]), .Z(n8811) );
  AND U13219 ( .A(n8813), .B(n8814), .Z(o[6034]) );
  AND U13220 ( .A(p_input[26034]), .B(p_input[16034]), .Z(n8814) );
  AND U13221 ( .A(p_input[6034]), .B(p_input[36034]), .Z(n8813) );
  AND U13222 ( .A(n8815), .B(n8816), .Z(o[6033]) );
  AND U13223 ( .A(p_input[26033]), .B(p_input[16033]), .Z(n8816) );
  AND U13224 ( .A(p_input[6033]), .B(p_input[36033]), .Z(n8815) );
  AND U13225 ( .A(n8817), .B(n8818), .Z(o[6032]) );
  AND U13226 ( .A(p_input[26032]), .B(p_input[16032]), .Z(n8818) );
  AND U13227 ( .A(p_input[6032]), .B(p_input[36032]), .Z(n8817) );
  AND U13228 ( .A(n8819), .B(n8820), .Z(o[6031]) );
  AND U13229 ( .A(p_input[26031]), .B(p_input[16031]), .Z(n8820) );
  AND U13230 ( .A(p_input[6031]), .B(p_input[36031]), .Z(n8819) );
  AND U13231 ( .A(n8821), .B(n8822), .Z(o[6030]) );
  AND U13232 ( .A(p_input[26030]), .B(p_input[16030]), .Z(n8822) );
  AND U13233 ( .A(p_input[6030]), .B(p_input[36030]), .Z(n8821) );
  AND U13234 ( .A(n8823), .B(n8824), .Z(o[602]) );
  AND U13235 ( .A(p_input[20602]), .B(p_input[10602]), .Z(n8824) );
  AND U13236 ( .A(p_input[602]), .B(p_input[30602]), .Z(n8823) );
  AND U13237 ( .A(n8825), .B(n8826), .Z(o[6029]) );
  AND U13238 ( .A(p_input[26029]), .B(p_input[16029]), .Z(n8826) );
  AND U13239 ( .A(p_input[6029]), .B(p_input[36029]), .Z(n8825) );
  AND U13240 ( .A(n8827), .B(n8828), .Z(o[6028]) );
  AND U13241 ( .A(p_input[26028]), .B(p_input[16028]), .Z(n8828) );
  AND U13242 ( .A(p_input[6028]), .B(p_input[36028]), .Z(n8827) );
  AND U13243 ( .A(n8829), .B(n8830), .Z(o[6027]) );
  AND U13244 ( .A(p_input[26027]), .B(p_input[16027]), .Z(n8830) );
  AND U13245 ( .A(p_input[6027]), .B(p_input[36027]), .Z(n8829) );
  AND U13246 ( .A(n8831), .B(n8832), .Z(o[6026]) );
  AND U13247 ( .A(p_input[26026]), .B(p_input[16026]), .Z(n8832) );
  AND U13248 ( .A(p_input[6026]), .B(p_input[36026]), .Z(n8831) );
  AND U13249 ( .A(n8833), .B(n8834), .Z(o[6025]) );
  AND U13250 ( .A(p_input[26025]), .B(p_input[16025]), .Z(n8834) );
  AND U13251 ( .A(p_input[6025]), .B(p_input[36025]), .Z(n8833) );
  AND U13252 ( .A(n8835), .B(n8836), .Z(o[6024]) );
  AND U13253 ( .A(p_input[26024]), .B(p_input[16024]), .Z(n8836) );
  AND U13254 ( .A(p_input[6024]), .B(p_input[36024]), .Z(n8835) );
  AND U13255 ( .A(n8837), .B(n8838), .Z(o[6023]) );
  AND U13256 ( .A(p_input[26023]), .B(p_input[16023]), .Z(n8838) );
  AND U13257 ( .A(p_input[6023]), .B(p_input[36023]), .Z(n8837) );
  AND U13258 ( .A(n8839), .B(n8840), .Z(o[6022]) );
  AND U13259 ( .A(p_input[26022]), .B(p_input[16022]), .Z(n8840) );
  AND U13260 ( .A(p_input[6022]), .B(p_input[36022]), .Z(n8839) );
  AND U13261 ( .A(n8841), .B(n8842), .Z(o[6021]) );
  AND U13262 ( .A(p_input[26021]), .B(p_input[16021]), .Z(n8842) );
  AND U13263 ( .A(p_input[6021]), .B(p_input[36021]), .Z(n8841) );
  AND U13264 ( .A(n8843), .B(n8844), .Z(o[6020]) );
  AND U13265 ( .A(p_input[26020]), .B(p_input[16020]), .Z(n8844) );
  AND U13266 ( .A(p_input[6020]), .B(p_input[36020]), .Z(n8843) );
  AND U13267 ( .A(n8845), .B(n8846), .Z(o[601]) );
  AND U13268 ( .A(p_input[20601]), .B(p_input[10601]), .Z(n8846) );
  AND U13269 ( .A(p_input[601]), .B(p_input[30601]), .Z(n8845) );
  AND U13270 ( .A(n8847), .B(n8848), .Z(o[6019]) );
  AND U13271 ( .A(p_input[26019]), .B(p_input[16019]), .Z(n8848) );
  AND U13272 ( .A(p_input[6019]), .B(p_input[36019]), .Z(n8847) );
  AND U13273 ( .A(n8849), .B(n8850), .Z(o[6018]) );
  AND U13274 ( .A(p_input[26018]), .B(p_input[16018]), .Z(n8850) );
  AND U13275 ( .A(p_input[6018]), .B(p_input[36018]), .Z(n8849) );
  AND U13276 ( .A(n8851), .B(n8852), .Z(o[6017]) );
  AND U13277 ( .A(p_input[26017]), .B(p_input[16017]), .Z(n8852) );
  AND U13278 ( .A(p_input[6017]), .B(p_input[36017]), .Z(n8851) );
  AND U13279 ( .A(n8853), .B(n8854), .Z(o[6016]) );
  AND U13280 ( .A(p_input[26016]), .B(p_input[16016]), .Z(n8854) );
  AND U13281 ( .A(p_input[6016]), .B(p_input[36016]), .Z(n8853) );
  AND U13282 ( .A(n8855), .B(n8856), .Z(o[6015]) );
  AND U13283 ( .A(p_input[26015]), .B(p_input[16015]), .Z(n8856) );
  AND U13284 ( .A(p_input[6015]), .B(p_input[36015]), .Z(n8855) );
  AND U13285 ( .A(n8857), .B(n8858), .Z(o[6014]) );
  AND U13286 ( .A(p_input[26014]), .B(p_input[16014]), .Z(n8858) );
  AND U13287 ( .A(p_input[6014]), .B(p_input[36014]), .Z(n8857) );
  AND U13288 ( .A(n8859), .B(n8860), .Z(o[6013]) );
  AND U13289 ( .A(p_input[26013]), .B(p_input[16013]), .Z(n8860) );
  AND U13290 ( .A(p_input[6013]), .B(p_input[36013]), .Z(n8859) );
  AND U13291 ( .A(n8861), .B(n8862), .Z(o[6012]) );
  AND U13292 ( .A(p_input[26012]), .B(p_input[16012]), .Z(n8862) );
  AND U13293 ( .A(p_input[6012]), .B(p_input[36012]), .Z(n8861) );
  AND U13294 ( .A(n8863), .B(n8864), .Z(o[6011]) );
  AND U13295 ( .A(p_input[26011]), .B(p_input[16011]), .Z(n8864) );
  AND U13296 ( .A(p_input[6011]), .B(p_input[36011]), .Z(n8863) );
  AND U13297 ( .A(n8865), .B(n8866), .Z(o[6010]) );
  AND U13298 ( .A(p_input[26010]), .B(p_input[16010]), .Z(n8866) );
  AND U13299 ( .A(p_input[6010]), .B(p_input[36010]), .Z(n8865) );
  AND U13300 ( .A(n8867), .B(n8868), .Z(o[600]) );
  AND U13301 ( .A(p_input[20600]), .B(p_input[10600]), .Z(n8868) );
  AND U13302 ( .A(p_input[600]), .B(p_input[30600]), .Z(n8867) );
  AND U13303 ( .A(n8869), .B(n8870), .Z(o[6009]) );
  AND U13304 ( .A(p_input[26009]), .B(p_input[16009]), .Z(n8870) );
  AND U13305 ( .A(p_input[6009]), .B(p_input[36009]), .Z(n8869) );
  AND U13306 ( .A(n8871), .B(n8872), .Z(o[6008]) );
  AND U13307 ( .A(p_input[26008]), .B(p_input[16008]), .Z(n8872) );
  AND U13308 ( .A(p_input[6008]), .B(p_input[36008]), .Z(n8871) );
  AND U13309 ( .A(n8873), .B(n8874), .Z(o[6007]) );
  AND U13310 ( .A(p_input[26007]), .B(p_input[16007]), .Z(n8874) );
  AND U13311 ( .A(p_input[6007]), .B(p_input[36007]), .Z(n8873) );
  AND U13312 ( .A(n8875), .B(n8876), .Z(o[6006]) );
  AND U13313 ( .A(p_input[26006]), .B(p_input[16006]), .Z(n8876) );
  AND U13314 ( .A(p_input[6006]), .B(p_input[36006]), .Z(n8875) );
  AND U13315 ( .A(n8877), .B(n8878), .Z(o[6005]) );
  AND U13316 ( .A(p_input[26005]), .B(p_input[16005]), .Z(n8878) );
  AND U13317 ( .A(p_input[6005]), .B(p_input[36005]), .Z(n8877) );
  AND U13318 ( .A(n8879), .B(n8880), .Z(o[6004]) );
  AND U13319 ( .A(p_input[26004]), .B(p_input[16004]), .Z(n8880) );
  AND U13320 ( .A(p_input[6004]), .B(p_input[36004]), .Z(n8879) );
  AND U13321 ( .A(n8881), .B(n8882), .Z(o[6003]) );
  AND U13322 ( .A(p_input[26003]), .B(p_input[16003]), .Z(n8882) );
  AND U13323 ( .A(p_input[6003]), .B(p_input[36003]), .Z(n8881) );
  AND U13324 ( .A(n8883), .B(n8884), .Z(o[6002]) );
  AND U13325 ( .A(p_input[26002]), .B(p_input[16002]), .Z(n8884) );
  AND U13326 ( .A(p_input[6002]), .B(p_input[36002]), .Z(n8883) );
  AND U13327 ( .A(n8885), .B(n8886), .Z(o[6001]) );
  AND U13328 ( .A(p_input[26001]), .B(p_input[16001]), .Z(n8886) );
  AND U13329 ( .A(p_input[6001]), .B(p_input[36001]), .Z(n8885) );
  AND U13330 ( .A(n8887), .B(n8888), .Z(o[6000]) );
  AND U13331 ( .A(p_input[26000]), .B(p_input[16000]), .Z(n8888) );
  AND U13332 ( .A(p_input[6000]), .B(p_input[36000]), .Z(n8887) );
  AND U13333 ( .A(n8889), .B(n8890), .Z(o[5]) );
  AND U13334 ( .A(p_input[20005]), .B(p_input[10005]), .Z(n8890) );
  AND U13335 ( .A(p_input[5]), .B(p_input[30005]), .Z(n8889) );
  AND U13336 ( .A(n8891), .B(n8892), .Z(o[59]) );
  AND U13337 ( .A(p_input[20059]), .B(p_input[10059]), .Z(n8892) );
  AND U13338 ( .A(p_input[59]), .B(p_input[30059]), .Z(n8891) );
  AND U13339 ( .A(n8893), .B(n8894), .Z(o[599]) );
  AND U13340 ( .A(p_input[20599]), .B(p_input[10599]), .Z(n8894) );
  AND U13341 ( .A(p_input[599]), .B(p_input[30599]), .Z(n8893) );
  AND U13342 ( .A(n8895), .B(n8896), .Z(o[5999]) );
  AND U13343 ( .A(p_input[25999]), .B(p_input[15999]), .Z(n8896) );
  AND U13344 ( .A(p_input[5999]), .B(p_input[35999]), .Z(n8895) );
  AND U13345 ( .A(n8897), .B(n8898), .Z(o[5998]) );
  AND U13346 ( .A(p_input[25998]), .B(p_input[15998]), .Z(n8898) );
  AND U13347 ( .A(p_input[5998]), .B(p_input[35998]), .Z(n8897) );
  AND U13348 ( .A(n8899), .B(n8900), .Z(o[5997]) );
  AND U13349 ( .A(p_input[25997]), .B(p_input[15997]), .Z(n8900) );
  AND U13350 ( .A(p_input[5997]), .B(p_input[35997]), .Z(n8899) );
  AND U13351 ( .A(n8901), .B(n8902), .Z(o[5996]) );
  AND U13352 ( .A(p_input[25996]), .B(p_input[15996]), .Z(n8902) );
  AND U13353 ( .A(p_input[5996]), .B(p_input[35996]), .Z(n8901) );
  AND U13354 ( .A(n8903), .B(n8904), .Z(o[5995]) );
  AND U13355 ( .A(p_input[25995]), .B(p_input[15995]), .Z(n8904) );
  AND U13356 ( .A(p_input[5995]), .B(p_input[35995]), .Z(n8903) );
  AND U13357 ( .A(n8905), .B(n8906), .Z(o[5994]) );
  AND U13358 ( .A(p_input[25994]), .B(p_input[15994]), .Z(n8906) );
  AND U13359 ( .A(p_input[5994]), .B(p_input[35994]), .Z(n8905) );
  AND U13360 ( .A(n8907), .B(n8908), .Z(o[5993]) );
  AND U13361 ( .A(p_input[25993]), .B(p_input[15993]), .Z(n8908) );
  AND U13362 ( .A(p_input[5993]), .B(p_input[35993]), .Z(n8907) );
  AND U13363 ( .A(n8909), .B(n8910), .Z(o[5992]) );
  AND U13364 ( .A(p_input[25992]), .B(p_input[15992]), .Z(n8910) );
  AND U13365 ( .A(p_input[5992]), .B(p_input[35992]), .Z(n8909) );
  AND U13366 ( .A(n8911), .B(n8912), .Z(o[5991]) );
  AND U13367 ( .A(p_input[25991]), .B(p_input[15991]), .Z(n8912) );
  AND U13368 ( .A(p_input[5991]), .B(p_input[35991]), .Z(n8911) );
  AND U13369 ( .A(n8913), .B(n8914), .Z(o[5990]) );
  AND U13370 ( .A(p_input[25990]), .B(p_input[15990]), .Z(n8914) );
  AND U13371 ( .A(p_input[5990]), .B(p_input[35990]), .Z(n8913) );
  AND U13372 ( .A(n8915), .B(n8916), .Z(o[598]) );
  AND U13373 ( .A(p_input[20598]), .B(p_input[10598]), .Z(n8916) );
  AND U13374 ( .A(p_input[598]), .B(p_input[30598]), .Z(n8915) );
  AND U13375 ( .A(n8917), .B(n8918), .Z(o[5989]) );
  AND U13376 ( .A(p_input[25989]), .B(p_input[15989]), .Z(n8918) );
  AND U13377 ( .A(p_input[5989]), .B(p_input[35989]), .Z(n8917) );
  AND U13378 ( .A(n8919), .B(n8920), .Z(o[5988]) );
  AND U13379 ( .A(p_input[25988]), .B(p_input[15988]), .Z(n8920) );
  AND U13380 ( .A(p_input[5988]), .B(p_input[35988]), .Z(n8919) );
  AND U13381 ( .A(n8921), .B(n8922), .Z(o[5987]) );
  AND U13382 ( .A(p_input[25987]), .B(p_input[15987]), .Z(n8922) );
  AND U13383 ( .A(p_input[5987]), .B(p_input[35987]), .Z(n8921) );
  AND U13384 ( .A(n8923), .B(n8924), .Z(o[5986]) );
  AND U13385 ( .A(p_input[25986]), .B(p_input[15986]), .Z(n8924) );
  AND U13386 ( .A(p_input[5986]), .B(p_input[35986]), .Z(n8923) );
  AND U13387 ( .A(n8925), .B(n8926), .Z(o[5985]) );
  AND U13388 ( .A(p_input[25985]), .B(p_input[15985]), .Z(n8926) );
  AND U13389 ( .A(p_input[5985]), .B(p_input[35985]), .Z(n8925) );
  AND U13390 ( .A(n8927), .B(n8928), .Z(o[5984]) );
  AND U13391 ( .A(p_input[25984]), .B(p_input[15984]), .Z(n8928) );
  AND U13392 ( .A(p_input[5984]), .B(p_input[35984]), .Z(n8927) );
  AND U13393 ( .A(n8929), .B(n8930), .Z(o[5983]) );
  AND U13394 ( .A(p_input[25983]), .B(p_input[15983]), .Z(n8930) );
  AND U13395 ( .A(p_input[5983]), .B(p_input[35983]), .Z(n8929) );
  AND U13396 ( .A(n8931), .B(n8932), .Z(o[5982]) );
  AND U13397 ( .A(p_input[25982]), .B(p_input[15982]), .Z(n8932) );
  AND U13398 ( .A(p_input[5982]), .B(p_input[35982]), .Z(n8931) );
  AND U13399 ( .A(n8933), .B(n8934), .Z(o[5981]) );
  AND U13400 ( .A(p_input[25981]), .B(p_input[15981]), .Z(n8934) );
  AND U13401 ( .A(p_input[5981]), .B(p_input[35981]), .Z(n8933) );
  AND U13402 ( .A(n8935), .B(n8936), .Z(o[5980]) );
  AND U13403 ( .A(p_input[25980]), .B(p_input[15980]), .Z(n8936) );
  AND U13404 ( .A(p_input[5980]), .B(p_input[35980]), .Z(n8935) );
  AND U13405 ( .A(n8937), .B(n8938), .Z(o[597]) );
  AND U13406 ( .A(p_input[20597]), .B(p_input[10597]), .Z(n8938) );
  AND U13407 ( .A(p_input[597]), .B(p_input[30597]), .Z(n8937) );
  AND U13408 ( .A(n8939), .B(n8940), .Z(o[5979]) );
  AND U13409 ( .A(p_input[25979]), .B(p_input[15979]), .Z(n8940) );
  AND U13410 ( .A(p_input[5979]), .B(p_input[35979]), .Z(n8939) );
  AND U13411 ( .A(n8941), .B(n8942), .Z(o[5978]) );
  AND U13412 ( .A(p_input[25978]), .B(p_input[15978]), .Z(n8942) );
  AND U13413 ( .A(p_input[5978]), .B(p_input[35978]), .Z(n8941) );
  AND U13414 ( .A(n8943), .B(n8944), .Z(o[5977]) );
  AND U13415 ( .A(p_input[25977]), .B(p_input[15977]), .Z(n8944) );
  AND U13416 ( .A(p_input[5977]), .B(p_input[35977]), .Z(n8943) );
  AND U13417 ( .A(n8945), .B(n8946), .Z(o[5976]) );
  AND U13418 ( .A(p_input[25976]), .B(p_input[15976]), .Z(n8946) );
  AND U13419 ( .A(p_input[5976]), .B(p_input[35976]), .Z(n8945) );
  AND U13420 ( .A(n8947), .B(n8948), .Z(o[5975]) );
  AND U13421 ( .A(p_input[25975]), .B(p_input[15975]), .Z(n8948) );
  AND U13422 ( .A(p_input[5975]), .B(p_input[35975]), .Z(n8947) );
  AND U13423 ( .A(n8949), .B(n8950), .Z(o[5974]) );
  AND U13424 ( .A(p_input[25974]), .B(p_input[15974]), .Z(n8950) );
  AND U13425 ( .A(p_input[5974]), .B(p_input[35974]), .Z(n8949) );
  AND U13426 ( .A(n8951), .B(n8952), .Z(o[5973]) );
  AND U13427 ( .A(p_input[25973]), .B(p_input[15973]), .Z(n8952) );
  AND U13428 ( .A(p_input[5973]), .B(p_input[35973]), .Z(n8951) );
  AND U13429 ( .A(n8953), .B(n8954), .Z(o[5972]) );
  AND U13430 ( .A(p_input[25972]), .B(p_input[15972]), .Z(n8954) );
  AND U13431 ( .A(p_input[5972]), .B(p_input[35972]), .Z(n8953) );
  AND U13432 ( .A(n8955), .B(n8956), .Z(o[5971]) );
  AND U13433 ( .A(p_input[25971]), .B(p_input[15971]), .Z(n8956) );
  AND U13434 ( .A(p_input[5971]), .B(p_input[35971]), .Z(n8955) );
  AND U13435 ( .A(n8957), .B(n8958), .Z(o[5970]) );
  AND U13436 ( .A(p_input[25970]), .B(p_input[15970]), .Z(n8958) );
  AND U13437 ( .A(p_input[5970]), .B(p_input[35970]), .Z(n8957) );
  AND U13438 ( .A(n8959), .B(n8960), .Z(o[596]) );
  AND U13439 ( .A(p_input[20596]), .B(p_input[10596]), .Z(n8960) );
  AND U13440 ( .A(p_input[596]), .B(p_input[30596]), .Z(n8959) );
  AND U13441 ( .A(n8961), .B(n8962), .Z(o[5969]) );
  AND U13442 ( .A(p_input[25969]), .B(p_input[15969]), .Z(n8962) );
  AND U13443 ( .A(p_input[5969]), .B(p_input[35969]), .Z(n8961) );
  AND U13444 ( .A(n8963), .B(n8964), .Z(o[5968]) );
  AND U13445 ( .A(p_input[25968]), .B(p_input[15968]), .Z(n8964) );
  AND U13446 ( .A(p_input[5968]), .B(p_input[35968]), .Z(n8963) );
  AND U13447 ( .A(n8965), .B(n8966), .Z(o[5967]) );
  AND U13448 ( .A(p_input[25967]), .B(p_input[15967]), .Z(n8966) );
  AND U13449 ( .A(p_input[5967]), .B(p_input[35967]), .Z(n8965) );
  AND U13450 ( .A(n8967), .B(n8968), .Z(o[5966]) );
  AND U13451 ( .A(p_input[25966]), .B(p_input[15966]), .Z(n8968) );
  AND U13452 ( .A(p_input[5966]), .B(p_input[35966]), .Z(n8967) );
  AND U13453 ( .A(n8969), .B(n8970), .Z(o[5965]) );
  AND U13454 ( .A(p_input[25965]), .B(p_input[15965]), .Z(n8970) );
  AND U13455 ( .A(p_input[5965]), .B(p_input[35965]), .Z(n8969) );
  AND U13456 ( .A(n8971), .B(n8972), .Z(o[5964]) );
  AND U13457 ( .A(p_input[25964]), .B(p_input[15964]), .Z(n8972) );
  AND U13458 ( .A(p_input[5964]), .B(p_input[35964]), .Z(n8971) );
  AND U13459 ( .A(n8973), .B(n8974), .Z(o[5963]) );
  AND U13460 ( .A(p_input[25963]), .B(p_input[15963]), .Z(n8974) );
  AND U13461 ( .A(p_input[5963]), .B(p_input[35963]), .Z(n8973) );
  AND U13462 ( .A(n8975), .B(n8976), .Z(o[5962]) );
  AND U13463 ( .A(p_input[25962]), .B(p_input[15962]), .Z(n8976) );
  AND U13464 ( .A(p_input[5962]), .B(p_input[35962]), .Z(n8975) );
  AND U13465 ( .A(n8977), .B(n8978), .Z(o[5961]) );
  AND U13466 ( .A(p_input[25961]), .B(p_input[15961]), .Z(n8978) );
  AND U13467 ( .A(p_input[5961]), .B(p_input[35961]), .Z(n8977) );
  AND U13468 ( .A(n8979), .B(n8980), .Z(o[5960]) );
  AND U13469 ( .A(p_input[25960]), .B(p_input[15960]), .Z(n8980) );
  AND U13470 ( .A(p_input[5960]), .B(p_input[35960]), .Z(n8979) );
  AND U13471 ( .A(n8981), .B(n8982), .Z(o[595]) );
  AND U13472 ( .A(p_input[20595]), .B(p_input[10595]), .Z(n8982) );
  AND U13473 ( .A(p_input[595]), .B(p_input[30595]), .Z(n8981) );
  AND U13474 ( .A(n8983), .B(n8984), .Z(o[5959]) );
  AND U13475 ( .A(p_input[25959]), .B(p_input[15959]), .Z(n8984) );
  AND U13476 ( .A(p_input[5959]), .B(p_input[35959]), .Z(n8983) );
  AND U13477 ( .A(n8985), .B(n8986), .Z(o[5958]) );
  AND U13478 ( .A(p_input[25958]), .B(p_input[15958]), .Z(n8986) );
  AND U13479 ( .A(p_input[5958]), .B(p_input[35958]), .Z(n8985) );
  AND U13480 ( .A(n8987), .B(n8988), .Z(o[5957]) );
  AND U13481 ( .A(p_input[25957]), .B(p_input[15957]), .Z(n8988) );
  AND U13482 ( .A(p_input[5957]), .B(p_input[35957]), .Z(n8987) );
  AND U13483 ( .A(n8989), .B(n8990), .Z(o[5956]) );
  AND U13484 ( .A(p_input[25956]), .B(p_input[15956]), .Z(n8990) );
  AND U13485 ( .A(p_input[5956]), .B(p_input[35956]), .Z(n8989) );
  AND U13486 ( .A(n8991), .B(n8992), .Z(o[5955]) );
  AND U13487 ( .A(p_input[25955]), .B(p_input[15955]), .Z(n8992) );
  AND U13488 ( .A(p_input[5955]), .B(p_input[35955]), .Z(n8991) );
  AND U13489 ( .A(n8993), .B(n8994), .Z(o[5954]) );
  AND U13490 ( .A(p_input[25954]), .B(p_input[15954]), .Z(n8994) );
  AND U13491 ( .A(p_input[5954]), .B(p_input[35954]), .Z(n8993) );
  AND U13492 ( .A(n8995), .B(n8996), .Z(o[5953]) );
  AND U13493 ( .A(p_input[25953]), .B(p_input[15953]), .Z(n8996) );
  AND U13494 ( .A(p_input[5953]), .B(p_input[35953]), .Z(n8995) );
  AND U13495 ( .A(n8997), .B(n8998), .Z(o[5952]) );
  AND U13496 ( .A(p_input[25952]), .B(p_input[15952]), .Z(n8998) );
  AND U13497 ( .A(p_input[5952]), .B(p_input[35952]), .Z(n8997) );
  AND U13498 ( .A(n8999), .B(n9000), .Z(o[5951]) );
  AND U13499 ( .A(p_input[25951]), .B(p_input[15951]), .Z(n9000) );
  AND U13500 ( .A(p_input[5951]), .B(p_input[35951]), .Z(n8999) );
  AND U13501 ( .A(n9001), .B(n9002), .Z(o[5950]) );
  AND U13502 ( .A(p_input[25950]), .B(p_input[15950]), .Z(n9002) );
  AND U13503 ( .A(p_input[5950]), .B(p_input[35950]), .Z(n9001) );
  AND U13504 ( .A(n9003), .B(n9004), .Z(o[594]) );
  AND U13505 ( .A(p_input[20594]), .B(p_input[10594]), .Z(n9004) );
  AND U13506 ( .A(p_input[594]), .B(p_input[30594]), .Z(n9003) );
  AND U13507 ( .A(n9005), .B(n9006), .Z(o[5949]) );
  AND U13508 ( .A(p_input[25949]), .B(p_input[15949]), .Z(n9006) );
  AND U13509 ( .A(p_input[5949]), .B(p_input[35949]), .Z(n9005) );
  AND U13510 ( .A(n9007), .B(n9008), .Z(o[5948]) );
  AND U13511 ( .A(p_input[25948]), .B(p_input[15948]), .Z(n9008) );
  AND U13512 ( .A(p_input[5948]), .B(p_input[35948]), .Z(n9007) );
  AND U13513 ( .A(n9009), .B(n9010), .Z(o[5947]) );
  AND U13514 ( .A(p_input[25947]), .B(p_input[15947]), .Z(n9010) );
  AND U13515 ( .A(p_input[5947]), .B(p_input[35947]), .Z(n9009) );
  AND U13516 ( .A(n9011), .B(n9012), .Z(o[5946]) );
  AND U13517 ( .A(p_input[25946]), .B(p_input[15946]), .Z(n9012) );
  AND U13518 ( .A(p_input[5946]), .B(p_input[35946]), .Z(n9011) );
  AND U13519 ( .A(n9013), .B(n9014), .Z(o[5945]) );
  AND U13520 ( .A(p_input[25945]), .B(p_input[15945]), .Z(n9014) );
  AND U13521 ( .A(p_input[5945]), .B(p_input[35945]), .Z(n9013) );
  AND U13522 ( .A(n9015), .B(n9016), .Z(o[5944]) );
  AND U13523 ( .A(p_input[25944]), .B(p_input[15944]), .Z(n9016) );
  AND U13524 ( .A(p_input[5944]), .B(p_input[35944]), .Z(n9015) );
  AND U13525 ( .A(n9017), .B(n9018), .Z(o[5943]) );
  AND U13526 ( .A(p_input[25943]), .B(p_input[15943]), .Z(n9018) );
  AND U13527 ( .A(p_input[5943]), .B(p_input[35943]), .Z(n9017) );
  AND U13528 ( .A(n9019), .B(n9020), .Z(o[5942]) );
  AND U13529 ( .A(p_input[25942]), .B(p_input[15942]), .Z(n9020) );
  AND U13530 ( .A(p_input[5942]), .B(p_input[35942]), .Z(n9019) );
  AND U13531 ( .A(n9021), .B(n9022), .Z(o[5941]) );
  AND U13532 ( .A(p_input[25941]), .B(p_input[15941]), .Z(n9022) );
  AND U13533 ( .A(p_input[5941]), .B(p_input[35941]), .Z(n9021) );
  AND U13534 ( .A(n9023), .B(n9024), .Z(o[5940]) );
  AND U13535 ( .A(p_input[25940]), .B(p_input[15940]), .Z(n9024) );
  AND U13536 ( .A(p_input[5940]), .B(p_input[35940]), .Z(n9023) );
  AND U13537 ( .A(n9025), .B(n9026), .Z(o[593]) );
  AND U13538 ( .A(p_input[20593]), .B(p_input[10593]), .Z(n9026) );
  AND U13539 ( .A(p_input[593]), .B(p_input[30593]), .Z(n9025) );
  AND U13540 ( .A(n9027), .B(n9028), .Z(o[5939]) );
  AND U13541 ( .A(p_input[25939]), .B(p_input[15939]), .Z(n9028) );
  AND U13542 ( .A(p_input[5939]), .B(p_input[35939]), .Z(n9027) );
  AND U13543 ( .A(n9029), .B(n9030), .Z(o[5938]) );
  AND U13544 ( .A(p_input[25938]), .B(p_input[15938]), .Z(n9030) );
  AND U13545 ( .A(p_input[5938]), .B(p_input[35938]), .Z(n9029) );
  AND U13546 ( .A(n9031), .B(n9032), .Z(o[5937]) );
  AND U13547 ( .A(p_input[25937]), .B(p_input[15937]), .Z(n9032) );
  AND U13548 ( .A(p_input[5937]), .B(p_input[35937]), .Z(n9031) );
  AND U13549 ( .A(n9033), .B(n9034), .Z(o[5936]) );
  AND U13550 ( .A(p_input[25936]), .B(p_input[15936]), .Z(n9034) );
  AND U13551 ( .A(p_input[5936]), .B(p_input[35936]), .Z(n9033) );
  AND U13552 ( .A(n9035), .B(n9036), .Z(o[5935]) );
  AND U13553 ( .A(p_input[25935]), .B(p_input[15935]), .Z(n9036) );
  AND U13554 ( .A(p_input[5935]), .B(p_input[35935]), .Z(n9035) );
  AND U13555 ( .A(n9037), .B(n9038), .Z(o[5934]) );
  AND U13556 ( .A(p_input[25934]), .B(p_input[15934]), .Z(n9038) );
  AND U13557 ( .A(p_input[5934]), .B(p_input[35934]), .Z(n9037) );
  AND U13558 ( .A(n9039), .B(n9040), .Z(o[5933]) );
  AND U13559 ( .A(p_input[25933]), .B(p_input[15933]), .Z(n9040) );
  AND U13560 ( .A(p_input[5933]), .B(p_input[35933]), .Z(n9039) );
  AND U13561 ( .A(n9041), .B(n9042), .Z(o[5932]) );
  AND U13562 ( .A(p_input[25932]), .B(p_input[15932]), .Z(n9042) );
  AND U13563 ( .A(p_input[5932]), .B(p_input[35932]), .Z(n9041) );
  AND U13564 ( .A(n9043), .B(n9044), .Z(o[5931]) );
  AND U13565 ( .A(p_input[25931]), .B(p_input[15931]), .Z(n9044) );
  AND U13566 ( .A(p_input[5931]), .B(p_input[35931]), .Z(n9043) );
  AND U13567 ( .A(n9045), .B(n9046), .Z(o[5930]) );
  AND U13568 ( .A(p_input[25930]), .B(p_input[15930]), .Z(n9046) );
  AND U13569 ( .A(p_input[5930]), .B(p_input[35930]), .Z(n9045) );
  AND U13570 ( .A(n9047), .B(n9048), .Z(o[592]) );
  AND U13571 ( .A(p_input[20592]), .B(p_input[10592]), .Z(n9048) );
  AND U13572 ( .A(p_input[592]), .B(p_input[30592]), .Z(n9047) );
  AND U13573 ( .A(n9049), .B(n9050), .Z(o[5929]) );
  AND U13574 ( .A(p_input[25929]), .B(p_input[15929]), .Z(n9050) );
  AND U13575 ( .A(p_input[5929]), .B(p_input[35929]), .Z(n9049) );
  AND U13576 ( .A(n9051), .B(n9052), .Z(o[5928]) );
  AND U13577 ( .A(p_input[25928]), .B(p_input[15928]), .Z(n9052) );
  AND U13578 ( .A(p_input[5928]), .B(p_input[35928]), .Z(n9051) );
  AND U13579 ( .A(n9053), .B(n9054), .Z(o[5927]) );
  AND U13580 ( .A(p_input[25927]), .B(p_input[15927]), .Z(n9054) );
  AND U13581 ( .A(p_input[5927]), .B(p_input[35927]), .Z(n9053) );
  AND U13582 ( .A(n9055), .B(n9056), .Z(o[5926]) );
  AND U13583 ( .A(p_input[25926]), .B(p_input[15926]), .Z(n9056) );
  AND U13584 ( .A(p_input[5926]), .B(p_input[35926]), .Z(n9055) );
  AND U13585 ( .A(n9057), .B(n9058), .Z(o[5925]) );
  AND U13586 ( .A(p_input[25925]), .B(p_input[15925]), .Z(n9058) );
  AND U13587 ( .A(p_input[5925]), .B(p_input[35925]), .Z(n9057) );
  AND U13588 ( .A(n9059), .B(n9060), .Z(o[5924]) );
  AND U13589 ( .A(p_input[25924]), .B(p_input[15924]), .Z(n9060) );
  AND U13590 ( .A(p_input[5924]), .B(p_input[35924]), .Z(n9059) );
  AND U13591 ( .A(n9061), .B(n9062), .Z(o[5923]) );
  AND U13592 ( .A(p_input[25923]), .B(p_input[15923]), .Z(n9062) );
  AND U13593 ( .A(p_input[5923]), .B(p_input[35923]), .Z(n9061) );
  AND U13594 ( .A(n9063), .B(n9064), .Z(o[5922]) );
  AND U13595 ( .A(p_input[25922]), .B(p_input[15922]), .Z(n9064) );
  AND U13596 ( .A(p_input[5922]), .B(p_input[35922]), .Z(n9063) );
  AND U13597 ( .A(n9065), .B(n9066), .Z(o[5921]) );
  AND U13598 ( .A(p_input[25921]), .B(p_input[15921]), .Z(n9066) );
  AND U13599 ( .A(p_input[5921]), .B(p_input[35921]), .Z(n9065) );
  AND U13600 ( .A(n9067), .B(n9068), .Z(o[5920]) );
  AND U13601 ( .A(p_input[25920]), .B(p_input[15920]), .Z(n9068) );
  AND U13602 ( .A(p_input[5920]), .B(p_input[35920]), .Z(n9067) );
  AND U13603 ( .A(n9069), .B(n9070), .Z(o[591]) );
  AND U13604 ( .A(p_input[20591]), .B(p_input[10591]), .Z(n9070) );
  AND U13605 ( .A(p_input[591]), .B(p_input[30591]), .Z(n9069) );
  AND U13606 ( .A(n9071), .B(n9072), .Z(o[5919]) );
  AND U13607 ( .A(p_input[25919]), .B(p_input[15919]), .Z(n9072) );
  AND U13608 ( .A(p_input[5919]), .B(p_input[35919]), .Z(n9071) );
  AND U13609 ( .A(n9073), .B(n9074), .Z(o[5918]) );
  AND U13610 ( .A(p_input[25918]), .B(p_input[15918]), .Z(n9074) );
  AND U13611 ( .A(p_input[5918]), .B(p_input[35918]), .Z(n9073) );
  AND U13612 ( .A(n9075), .B(n9076), .Z(o[5917]) );
  AND U13613 ( .A(p_input[25917]), .B(p_input[15917]), .Z(n9076) );
  AND U13614 ( .A(p_input[5917]), .B(p_input[35917]), .Z(n9075) );
  AND U13615 ( .A(n9077), .B(n9078), .Z(o[5916]) );
  AND U13616 ( .A(p_input[25916]), .B(p_input[15916]), .Z(n9078) );
  AND U13617 ( .A(p_input[5916]), .B(p_input[35916]), .Z(n9077) );
  AND U13618 ( .A(n9079), .B(n9080), .Z(o[5915]) );
  AND U13619 ( .A(p_input[25915]), .B(p_input[15915]), .Z(n9080) );
  AND U13620 ( .A(p_input[5915]), .B(p_input[35915]), .Z(n9079) );
  AND U13621 ( .A(n9081), .B(n9082), .Z(o[5914]) );
  AND U13622 ( .A(p_input[25914]), .B(p_input[15914]), .Z(n9082) );
  AND U13623 ( .A(p_input[5914]), .B(p_input[35914]), .Z(n9081) );
  AND U13624 ( .A(n9083), .B(n9084), .Z(o[5913]) );
  AND U13625 ( .A(p_input[25913]), .B(p_input[15913]), .Z(n9084) );
  AND U13626 ( .A(p_input[5913]), .B(p_input[35913]), .Z(n9083) );
  AND U13627 ( .A(n9085), .B(n9086), .Z(o[5912]) );
  AND U13628 ( .A(p_input[25912]), .B(p_input[15912]), .Z(n9086) );
  AND U13629 ( .A(p_input[5912]), .B(p_input[35912]), .Z(n9085) );
  AND U13630 ( .A(n9087), .B(n9088), .Z(o[5911]) );
  AND U13631 ( .A(p_input[25911]), .B(p_input[15911]), .Z(n9088) );
  AND U13632 ( .A(p_input[5911]), .B(p_input[35911]), .Z(n9087) );
  AND U13633 ( .A(n9089), .B(n9090), .Z(o[5910]) );
  AND U13634 ( .A(p_input[25910]), .B(p_input[15910]), .Z(n9090) );
  AND U13635 ( .A(p_input[5910]), .B(p_input[35910]), .Z(n9089) );
  AND U13636 ( .A(n9091), .B(n9092), .Z(o[590]) );
  AND U13637 ( .A(p_input[20590]), .B(p_input[10590]), .Z(n9092) );
  AND U13638 ( .A(p_input[590]), .B(p_input[30590]), .Z(n9091) );
  AND U13639 ( .A(n9093), .B(n9094), .Z(o[5909]) );
  AND U13640 ( .A(p_input[25909]), .B(p_input[15909]), .Z(n9094) );
  AND U13641 ( .A(p_input[5909]), .B(p_input[35909]), .Z(n9093) );
  AND U13642 ( .A(n9095), .B(n9096), .Z(o[5908]) );
  AND U13643 ( .A(p_input[25908]), .B(p_input[15908]), .Z(n9096) );
  AND U13644 ( .A(p_input[5908]), .B(p_input[35908]), .Z(n9095) );
  AND U13645 ( .A(n9097), .B(n9098), .Z(o[5907]) );
  AND U13646 ( .A(p_input[25907]), .B(p_input[15907]), .Z(n9098) );
  AND U13647 ( .A(p_input[5907]), .B(p_input[35907]), .Z(n9097) );
  AND U13648 ( .A(n9099), .B(n9100), .Z(o[5906]) );
  AND U13649 ( .A(p_input[25906]), .B(p_input[15906]), .Z(n9100) );
  AND U13650 ( .A(p_input[5906]), .B(p_input[35906]), .Z(n9099) );
  AND U13651 ( .A(n9101), .B(n9102), .Z(o[5905]) );
  AND U13652 ( .A(p_input[25905]), .B(p_input[15905]), .Z(n9102) );
  AND U13653 ( .A(p_input[5905]), .B(p_input[35905]), .Z(n9101) );
  AND U13654 ( .A(n9103), .B(n9104), .Z(o[5904]) );
  AND U13655 ( .A(p_input[25904]), .B(p_input[15904]), .Z(n9104) );
  AND U13656 ( .A(p_input[5904]), .B(p_input[35904]), .Z(n9103) );
  AND U13657 ( .A(n9105), .B(n9106), .Z(o[5903]) );
  AND U13658 ( .A(p_input[25903]), .B(p_input[15903]), .Z(n9106) );
  AND U13659 ( .A(p_input[5903]), .B(p_input[35903]), .Z(n9105) );
  AND U13660 ( .A(n9107), .B(n9108), .Z(o[5902]) );
  AND U13661 ( .A(p_input[25902]), .B(p_input[15902]), .Z(n9108) );
  AND U13662 ( .A(p_input[5902]), .B(p_input[35902]), .Z(n9107) );
  AND U13663 ( .A(n9109), .B(n9110), .Z(o[5901]) );
  AND U13664 ( .A(p_input[25901]), .B(p_input[15901]), .Z(n9110) );
  AND U13665 ( .A(p_input[5901]), .B(p_input[35901]), .Z(n9109) );
  AND U13666 ( .A(n9111), .B(n9112), .Z(o[5900]) );
  AND U13667 ( .A(p_input[25900]), .B(p_input[15900]), .Z(n9112) );
  AND U13668 ( .A(p_input[5900]), .B(p_input[35900]), .Z(n9111) );
  AND U13669 ( .A(n9113), .B(n9114), .Z(o[58]) );
  AND U13670 ( .A(p_input[20058]), .B(p_input[10058]), .Z(n9114) );
  AND U13671 ( .A(p_input[58]), .B(p_input[30058]), .Z(n9113) );
  AND U13672 ( .A(n9115), .B(n9116), .Z(o[589]) );
  AND U13673 ( .A(p_input[20589]), .B(p_input[10589]), .Z(n9116) );
  AND U13674 ( .A(p_input[589]), .B(p_input[30589]), .Z(n9115) );
  AND U13675 ( .A(n9117), .B(n9118), .Z(o[5899]) );
  AND U13676 ( .A(p_input[25899]), .B(p_input[15899]), .Z(n9118) );
  AND U13677 ( .A(p_input[5899]), .B(p_input[35899]), .Z(n9117) );
  AND U13678 ( .A(n9119), .B(n9120), .Z(o[5898]) );
  AND U13679 ( .A(p_input[25898]), .B(p_input[15898]), .Z(n9120) );
  AND U13680 ( .A(p_input[5898]), .B(p_input[35898]), .Z(n9119) );
  AND U13681 ( .A(n9121), .B(n9122), .Z(o[5897]) );
  AND U13682 ( .A(p_input[25897]), .B(p_input[15897]), .Z(n9122) );
  AND U13683 ( .A(p_input[5897]), .B(p_input[35897]), .Z(n9121) );
  AND U13684 ( .A(n9123), .B(n9124), .Z(o[5896]) );
  AND U13685 ( .A(p_input[25896]), .B(p_input[15896]), .Z(n9124) );
  AND U13686 ( .A(p_input[5896]), .B(p_input[35896]), .Z(n9123) );
  AND U13687 ( .A(n9125), .B(n9126), .Z(o[5895]) );
  AND U13688 ( .A(p_input[25895]), .B(p_input[15895]), .Z(n9126) );
  AND U13689 ( .A(p_input[5895]), .B(p_input[35895]), .Z(n9125) );
  AND U13690 ( .A(n9127), .B(n9128), .Z(o[5894]) );
  AND U13691 ( .A(p_input[25894]), .B(p_input[15894]), .Z(n9128) );
  AND U13692 ( .A(p_input[5894]), .B(p_input[35894]), .Z(n9127) );
  AND U13693 ( .A(n9129), .B(n9130), .Z(o[5893]) );
  AND U13694 ( .A(p_input[25893]), .B(p_input[15893]), .Z(n9130) );
  AND U13695 ( .A(p_input[5893]), .B(p_input[35893]), .Z(n9129) );
  AND U13696 ( .A(n9131), .B(n9132), .Z(o[5892]) );
  AND U13697 ( .A(p_input[25892]), .B(p_input[15892]), .Z(n9132) );
  AND U13698 ( .A(p_input[5892]), .B(p_input[35892]), .Z(n9131) );
  AND U13699 ( .A(n9133), .B(n9134), .Z(o[5891]) );
  AND U13700 ( .A(p_input[25891]), .B(p_input[15891]), .Z(n9134) );
  AND U13701 ( .A(p_input[5891]), .B(p_input[35891]), .Z(n9133) );
  AND U13702 ( .A(n9135), .B(n9136), .Z(o[5890]) );
  AND U13703 ( .A(p_input[25890]), .B(p_input[15890]), .Z(n9136) );
  AND U13704 ( .A(p_input[5890]), .B(p_input[35890]), .Z(n9135) );
  AND U13705 ( .A(n9137), .B(n9138), .Z(o[588]) );
  AND U13706 ( .A(p_input[20588]), .B(p_input[10588]), .Z(n9138) );
  AND U13707 ( .A(p_input[588]), .B(p_input[30588]), .Z(n9137) );
  AND U13708 ( .A(n9139), .B(n9140), .Z(o[5889]) );
  AND U13709 ( .A(p_input[25889]), .B(p_input[15889]), .Z(n9140) );
  AND U13710 ( .A(p_input[5889]), .B(p_input[35889]), .Z(n9139) );
  AND U13711 ( .A(n9141), .B(n9142), .Z(o[5888]) );
  AND U13712 ( .A(p_input[25888]), .B(p_input[15888]), .Z(n9142) );
  AND U13713 ( .A(p_input[5888]), .B(p_input[35888]), .Z(n9141) );
  AND U13714 ( .A(n9143), .B(n9144), .Z(o[5887]) );
  AND U13715 ( .A(p_input[25887]), .B(p_input[15887]), .Z(n9144) );
  AND U13716 ( .A(p_input[5887]), .B(p_input[35887]), .Z(n9143) );
  AND U13717 ( .A(n9145), .B(n9146), .Z(o[5886]) );
  AND U13718 ( .A(p_input[25886]), .B(p_input[15886]), .Z(n9146) );
  AND U13719 ( .A(p_input[5886]), .B(p_input[35886]), .Z(n9145) );
  AND U13720 ( .A(n9147), .B(n9148), .Z(o[5885]) );
  AND U13721 ( .A(p_input[25885]), .B(p_input[15885]), .Z(n9148) );
  AND U13722 ( .A(p_input[5885]), .B(p_input[35885]), .Z(n9147) );
  AND U13723 ( .A(n9149), .B(n9150), .Z(o[5884]) );
  AND U13724 ( .A(p_input[25884]), .B(p_input[15884]), .Z(n9150) );
  AND U13725 ( .A(p_input[5884]), .B(p_input[35884]), .Z(n9149) );
  AND U13726 ( .A(n9151), .B(n9152), .Z(o[5883]) );
  AND U13727 ( .A(p_input[25883]), .B(p_input[15883]), .Z(n9152) );
  AND U13728 ( .A(p_input[5883]), .B(p_input[35883]), .Z(n9151) );
  AND U13729 ( .A(n9153), .B(n9154), .Z(o[5882]) );
  AND U13730 ( .A(p_input[25882]), .B(p_input[15882]), .Z(n9154) );
  AND U13731 ( .A(p_input[5882]), .B(p_input[35882]), .Z(n9153) );
  AND U13732 ( .A(n9155), .B(n9156), .Z(o[5881]) );
  AND U13733 ( .A(p_input[25881]), .B(p_input[15881]), .Z(n9156) );
  AND U13734 ( .A(p_input[5881]), .B(p_input[35881]), .Z(n9155) );
  AND U13735 ( .A(n9157), .B(n9158), .Z(o[5880]) );
  AND U13736 ( .A(p_input[25880]), .B(p_input[15880]), .Z(n9158) );
  AND U13737 ( .A(p_input[5880]), .B(p_input[35880]), .Z(n9157) );
  AND U13738 ( .A(n9159), .B(n9160), .Z(o[587]) );
  AND U13739 ( .A(p_input[20587]), .B(p_input[10587]), .Z(n9160) );
  AND U13740 ( .A(p_input[587]), .B(p_input[30587]), .Z(n9159) );
  AND U13741 ( .A(n9161), .B(n9162), .Z(o[5879]) );
  AND U13742 ( .A(p_input[25879]), .B(p_input[15879]), .Z(n9162) );
  AND U13743 ( .A(p_input[5879]), .B(p_input[35879]), .Z(n9161) );
  AND U13744 ( .A(n9163), .B(n9164), .Z(o[5878]) );
  AND U13745 ( .A(p_input[25878]), .B(p_input[15878]), .Z(n9164) );
  AND U13746 ( .A(p_input[5878]), .B(p_input[35878]), .Z(n9163) );
  AND U13747 ( .A(n9165), .B(n9166), .Z(o[5877]) );
  AND U13748 ( .A(p_input[25877]), .B(p_input[15877]), .Z(n9166) );
  AND U13749 ( .A(p_input[5877]), .B(p_input[35877]), .Z(n9165) );
  AND U13750 ( .A(n9167), .B(n9168), .Z(o[5876]) );
  AND U13751 ( .A(p_input[25876]), .B(p_input[15876]), .Z(n9168) );
  AND U13752 ( .A(p_input[5876]), .B(p_input[35876]), .Z(n9167) );
  AND U13753 ( .A(n9169), .B(n9170), .Z(o[5875]) );
  AND U13754 ( .A(p_input[25875]), .B(p_input[15875]), .Z(n9170) );
  AND U13755 ( .A(p_input[5875]), .B(p_input[35875]), .Z(n9169) );
  AND U13756 ( .A(n9171), .B(n9172), .Z(o[5874]) );
  AND U13757 ( .A(p_input[25874]), .B(p_input[15874]), .Z(n9172) );
  AND U13758 ( .A(p_input[5874]), .B(p_input[35874]), .Z(n9171) );
  AND U13759 ( .A(n9173), .B(n9174), .Z(o[5873]) );
  AND U13760 ( .A(p_input[25873]), .B(p_input[15873]), .Z(n9174) );
  AND U13761 ( .A(p_input[5873]), .B(p_input[35873]), .Z(n9173) );
  AND U13762 ( .A(n9175), .B(n9176), .Z(o[5872]) );
  AND U13763 ( .A(p_input[25872]), .B(p_input[15872]), .Z(n9176) );
  AND U13764 ( .A(p_input[5872]), .B(p_input[35872]), .Z(n9175) );
  AND U13765 ( .A(n9177), .B(n9178), .Z(o[5871]) );
  AND U13766 ( .A(p_input[25871]), .B(p_input[15871]), .Z(n9178) );
  AND U13767 ( .A(p_input[5871]), .B(p_input[35871]), .Z(n9177) );
  AND U13768 ( .A(n9179), .B(n9180), .Z(o[5870]) );
  AND U13769 ( .A(p_input[25870]), .B(p_input[15870]), .Z(n9180) );
  AND U13770 ( .A(p_input[5870]), .B(p_input[35870]), .Z(n9179) );
  AND U13771 ( .A(n9181), .B(n9182), .Z(o[586]) );
  AND U13772 ( .A(p_input[20586]), .B(p_input[10586]), .Z(n9182) );
  AND U13773 ( .A(p_input[586]), .B(p_input[30586]), .Z(n9181) );
  AND U13774 ( .A(n9183), .B(n9184), .Z(o[5869]) );
  AND U13775 ( .A(p_input[25869]), .B(p_input[15869]), .Z(n9184) );
  AND U13776 ( .A(p_input[5869]), .B(p_input[35869]), .Z(n9183) );
  AND U13777 ( .A(n9185), .B(n9186), .Z(o[5868]) );
  AND U13778 ( .A(p_input[25868]), .B(p_input[15868]), .Z(n9186) );
  AND U13779 ( .A(p_input[5868]), .B(p_input[35868]), .Z(n9185) );
  AND U13780 ( .A(n9187), .B(n9188), .Z(o[5867]) );
  AND U13781 ( .A(p_input[25867]), .B(p_input[15867]), .Z(n9188) );
  AND U13782 ( .A(p_input[5867]), .B(p_input[35867]), .Z(n9187) );
  AND U13783 ( .A(n9189), .B(n9190), .Z(o[5866]) );
  AND U13784 ( .A(p_input[25866]), .B(p_input[15866]), .Z(n9190) );
  AND U13785 ( .A(p_input[5866]), .B(p_input[35866]), .Z(n9189) );
  AND U13786 ( .A(n9191), .B(n9192), .Z(o[5865]) );
  AND U13787 ( .A(p_input[25865]), .B(p_input[15865]), .Z(n9192) );
  AND U13788 ( .A(p_input[5865]), .B(p_input[35865]), .Z(n9191) );
  AND U13789 ( .A(n9193), .B(n9194), .Z(o[5864]) );
  AND U13790 ( .A(p_input[25864]), .B(p_input[15864]), .Z(n9194) );
  AND U13791 ( .A(p_input[5864]), .B(p_input[35864]), .Z(n9193) );
  AND U13792 ( .A(n9195), .B(n9196), .Z(o[5863]) );
  AND U13793 ( .A(p_input[25863]), .B(p_input[15863]), .Z(n9196) );
  AND U13794 ( .A(p_input[5863]), .B(p_input[35863]), .Z(n9195) );
  AND U13795 ( .A(n9197), .B(n9198), .Z(o[5862]) );
  AND U13796 ( .A(p_input[25862]), .B(p_input[15862]), .Z(n9198) );
  AND U13797 ( .A(p_input[5862]), .B(p_input[35862]), .Z(n9197) );
  AND U13798 ( .A(n9199), .B(n9200), .Z(o[5861]) );
  AND U13799 ( .A(p_input[25861]), .B(p_input[15861]), .Z(n9200) );
  AND U13800 ( .A(p_input[5861]), .B(p_input[35861]), .Z(n9199) );
  AND U13801 ( .A(n9201), .B(n9202), .Z(o[5860]) );
  AND U13802 ( .A(p_input[25860]), .B(p_input[15860]), .Z(n9202) );
  AND U13803 ( .A(p_input[5860]), .B(p_input[35860]), .Z(n9201) );
  AND U13804 ( .A(n9203), .B(n9204), .Z(o[585]) );
  AND U13805 ( .A(p_input[20585]), .B(p_input[10585]), .Z(n9204) );
  AND U13806 ( .A(p_input[585]), .B(p_input[30585]), .Z(n9203) );
  AND U13807 ( .A(n9205), .B(n9206), .Z(o[5859]) );
  AND U13808 ( .A(p_input[25859]), .B(p_input[15859]), .Z(n9206) );
  AND U13809 ( .A(p_input[5859]), .B(p_input[35859]), .Z(n9205) );
  AND U13810 ( .A(n9207), .B(n9208), .Z(o[5858]) );
  AND U13811 ( .A(p_input[25858]), .B(p_input[15858]), .Z(n9208) );
  AND U13812 ( .A(p_input[5858]), .B(p_input[35858]), .Z(n9207) );
  AND U13813 ( .A(n9209), .B(n9210), .Z(o[5857]) );
  AND U13814 ( .A(p_input[25857]), .B(p_input[15857]), .Z(n9210) );
  AND U13815 ( .A(p_input[5857]), .B(p_input[35857]), .Z(n9209) );
  AND U13816 ( .A(n9211), .B(n9212), .Z(o[5856]) );
  AND U13817 ( .A(p_input[25856]), .B(p_input[15856]), .Z(n9212) );
  AND U13818 ( .A(p_input[5856]), .B(p_input[35856]), .Z(n9211) );
  AND U13819 ( .A(n9213), .B(n9214), .Z(o[5855]) );
  AND U13820 ( .A(p_input[25855]), .B(p_input[15855]), .Z(n9214) );
  AND U13821 ( .A(p_input[5855]), .B(p_input[35855]), .Z(n9213) );
  AND U13822 ( .A(n9215), .B(n9216), .Z(o[5854]) );
  AND U13823 ( .A(p_input[25854]), .B(p_input[15854]), .Z(n9216) );
  AND U13824 ( .A(p_input[5854]), .B(p_input[35854]), .Z(n9215) );
  AND U13825 ( .A(n9217), .B(n9218), .Z(o[5853]) );
  AND U13826 ( .A(p_input[25853]), .B(p_input[15853]), .Z(n9218) );
  AND U13827 ( .A(p_input[5853]), .B(p_input[35853]), .Z(n9217) );
  AND U13828 ( .A(n9219), .B(n9220), .Z(o[5852]) );
  AND U13829 ( .A(p_input[25852]), .B(p_input[15852]), .Z(n9220) );
  AND U13830 ( .A(p_input[5852]), .B(p_input[35852]), .Z(n9219) );
  AND U13831 ( .A(n9221), .B(n9222), .Z(o[5851]) );
  AND U13832 ( .A(p_input[25851]), .B(p_input[15851]), .Z(n9222) );
  AND U13833 ( .A(p_input[5851]), .B(p_input[35851]), .Z(n9221) );
  AND U13834 ( .A(n9223), .B(n9224), .Z(o[5850]) );
  AND U13835 ( .A(p_input[25850]), .B(p_input[15850]), .Z(n9224) );
  AND U13836 ( .A(p_input[5850]), .B(p_input[35850]), .Z(n9223) );
  AND U13837 ( .A(n9225), .B(n9226), .Z(o[584]) );
  AND U13838 ( .A(p_input[20584]), .B(p_input[10584]), .Z(n9226) );
  AND U13839 ( .A(p_input[584]), .B(p_input[30584]), .Z(n9225) );
  AND U13840 ( .A(n9227), .B(n9228), .Z(o[5849]) );
  AND U13841 ( .A(p_input[25849]), .B(p_input[15849]), .Z(n9228) );
  AND U13842 ( .A(p_input[5849]), .B(p_input[35849]), .Z(n9227) );
  AND U13843 ( .A(n9229), .B(n9230), .Z(o[5848]) );
  AND U13844 ( .A(p_input[25848]), .B(p_input[15848]), .Z(n9230) );
  AND U13845 ( .A(p_input[5848]), .B(p_input[35848]), .Z(n9229) );
  AND U13846 ( .A(n9231), .B(n9232), .Z(o[5847]) );
  AND U13847 ( .A(p_input[25847]), .B(p_input[15847]), .Z(n9232) );
  AND U13848 ( .A(p_input[5847]), .B(p_input[35847]), .Z(n9231) );
  AND U13849 ( .A(n9233), .B(n9234), .Z(o[5846]) );
  AND U13850 ( .A(p_input[25846]), .B(p_input[15846]), .Z(n9234) );
  AND U13851 ( .A(p_input[5846]), .B(p_input[35846]), .Z(n9233) );
  AND U13852 ( .A(n9235), .B(n9236), .Z(o[5845]) );
  AND U13853 ( .A(p_input[25845]), .B(p_input[15845]), .Z(n9236) );
  AND U13854 ( .A(p_input[5845]), .B(p_input[35845]), .Z(n9235) );
  AND U13855 ( .A(n9237), .B(n9238), .Z(o[5844]) );
  AND U13856 ( .A(p_input[25844]), .B(p_input[15844]), .Z(n9238) );
  AND U13857 ( .A(p_input[5844]), .B(p_input[35844]), .Z(n9237) );
  AND U13858 ( .A(n9239), .B(n9240), .Z(o[5843]) );
  AND U13859 ( .A(p_input[25843]), .B(p_input[15843]), .Z(n9240) );
  AND U13860 ( .A(p_input[5843]), .B(p_input[35843]), .Z(n9239) );
  AND U13861 ( .A(n9241), .B(n9242), .Z(o[5842]) );
  AND U13862 ( .A(p_input[25842]), .B(p_input[15842]), .Z(n9242) );
  AND U13863 ( .A(p_input[5842]), .B(p_input[35842]), .Z(n9241) );
  AND U13864 ( .A(n9243), .B(n9244), .Z(o[5841]) );
  AND U13865 ( .A(p_input[25841]), .B(p_input[15841]), .Z(n9244) );
  AND U13866 ( .A(p_input[5841]), .B(p_input[35841]), .Z(n9243) );
  AND U13867 ( .A(n9245), .B(n9246), .Z(o[5840]) );
  AND U13868 ( .A(p_input[25840]), .B(p_input[15840]), .Z(n9246) );
  AND U13869 ( .A(p_input[5840]), .B(p_input[35840]), .Z(n9245) );
  AND U13870 ( .A(n9247), .B(n9248), .Z(o[583]) );
  AND U13871 ( .A(p_input[20583]), .B(p_input[10583]), .Z(n9248) );
  AND U13872 ( .A(p_input[583]), .B(p_input[30583]), .Z(n9247) );
  AND U13873 ( .A(n9249), .B(n9250), .Z(o[5839]) );
  AND U13874 ( .A(p_input[25839]), .B(p_input[15839]), .Z(n9250) );
  AND U13875 ( .A(p_input[5839]), .B(p_input[35839]), .Z(n9249) );
  AND U13876 ( .A(n9251), .B(n9252), .Z(o[5838]) );
  AND U13877 ( .A(p_input[25838]), .B(p_input[15838]), .Z(n9252) );
  AND U13878 ( .A(p_input[5838]), .B(p_input[35838]), .Z(n9251) );
  AND U13879 ( .A(n9253), .B(n9254), .Z(o[5837]) );
  AND U13880 ( .A(p_input[25837]), .B(p_input[15837]), .Z(n9254) );
  AND U13881 ( .A(p_input[5837]), .B(p_input[35837]), .Z(n9253) );
  AND U13882 ( .A(n9255), .B(n9256), .Z(o[5836]) );
  AND U13883 ( .A(p_input[25836]), .B(p_input[15836]), .Z(n9256) );
  AND U13884 ( .A(p_input[5836]), .B(p_input[35836]), .Z(n9255) );
  AND U13885 ( .A(n9257), .B(n9258), .Z(o[5835]) );
  AND U13886 ( .A(p_input[25835]), .B(p_input[15835]), .Z(n9258) );
  AND U13887 ( .A(p_input[5835]), .B(p_input[35835]), .Z(n9257) );
  AND U13888 ( .A(n9259), .B(n9260), .Z(o[5834]) );
  AND U13889 ( .A(p_input[25834]), .B(p_input[15834]), .Z(n9260) );
  AND U13890 ( .A(p_input[5834]), .B(p_input[35834]), .Z(n9259) );
  AND U13891 ( .A(n9261), .B(n9262), .Z(o[5833]) );
  AND U13892 ( .A(p_input[25833]), .B(p_input[15833]), .Z(n9262) );
  AND U13893 ( .A(p_input[5833]), .B(p_input[35833]), .Z(n9261) );
  AND U13894 ( .A(n9263), .B(n9264), .Z(o[5832]) );
  AND U13895 ( .A(p_input[25832]), .B(p_input[15832]), .Z(n9264) );
  AND U13896 ( .A(p_input[5832]), .B(p_input[35832]), .Z(n9263) );
  AND U13897 ( .A(n9265), .B(n9266), .Z(o[5831]) );
  AND U13898 ( .A(p_input[25831]), .B(p_input[15831]), .Z(n9266) );
  AND U13899 ( .A(p_input[5831]), .B(p_input[35831]), .Z(n9265) );
  AND U13900 ( .A(n9267), .B(n9268), .Z(o[5830]) );
  AND U13901 ( .A(p_input[25830]), .B(p_input[15830]), .Z(n9268) );
  AND U13902 ( .A(p_input[5830]), .B(p_input[35830]), .Z(n9267) );
  AND U13903 ( .A(n9269), .B(n9270), .Z(o[582]) );
  AND U13904 ( .A(p_input[20582]), .B(p_input[10582]), .Z(n9270) );
  AND U13905 ( .A(p_input[582]), .B(p_input[30582]), .Z(n9269) );
  AND U13906 ( .A(n9271), .B(n9272), .Z(o[5829]) );
  AND U13907 ( .A(p_input[25829]), .B(p_input[15829]), .Z(n9272) );
  AND U13908 ( .A(p_input[5829]), .B(p_input[35829]), .Z(n9271) );
  AND U13909 ( .A(n9273), .B(n9274), .Z(o[5828]) );
  AND U13910 ( .A(p_input[25828]), .B(p_input[15828]), .Z(n9274) );
  AND U13911 ( .A(p_input[5828]), .B(p_input[35828]), .Z(n9273) );
  AND U13912 ( .A(n9275), .B(n9276), .Z(o[5827]) );
  AND U13913 ( .A(p_input[25827]), .B(p_input[15827]), .Z(n9276) );
  AND U13914 ( .A(p_input[5827]), .B(p_input[35827]), .Z(n9275) );
  AND U13915 ( .A(n9277), .B(n9278), .Z(o[5826]) );
  AND U13916 ( .A(p_input[25826]), .B(p_input[15826]), .Z(n9278) );
  AND U13917 ( .A(p_input[5826]), .B(p_input[35826]), .Z(n9277) );
  AND U13918 ( .A(n9279), .B(n9280), .Z(o[5825]) );
  AND U13919 ( .A(p_input[25825]), .B(p_input[15825]), .Z(n9280) );
  AND U13920 ( .A(p_input[5825]), .B(p_input[35825]), .Z(n9279) );
  AND U13921 ( .A(n9281), .B(n9282), .Z(o[5824]) );
  AND U13922 ( .A(p_input[25824]), .B(p_input[15824]), .Z(n9282) );
  AND U13923 ( .A(p_input[5824]), .B(p_input[35824]), .Z(n9281) );
  AND U13924 ( .A(n9283), .B(n9284), .Z(o[5823]) );
  AND U13925 ( .A(p_input[25823]), .B(p_input[15823]), .Z(n9284) );
  AND U13926 ( .A(p_input[5823]), .B(p_input[35823]), .Z(n9283) );
  AND U13927 ( .A(n9285), .B(n9286), .Z(o[5822]) );
  AND U13928 ( .A(p_input[25822]), .B(p_input[15822]), .Z(n9286) );
  AND U13929 ( .A(p_input[5822]), .B(p_input[35822]), .Z(n9285) );
  AND U13930 ( .A(n9287), .B(n9288), .Z(o[5821]) );
  AND U13931 ( .A(p_input[25821]), .B(p_input[15821]), .Z(n9288) );
  AND U13932 ( .A(p_input[5821]), .B(p_input[35821]), .Z(n9287) );
  AND U13933 ( .A(n9289), .B(n9290), .Z(o[5820]) );
  AND U13934 ( .A(p_input[25820]), .B(p_input[15820]), .Z(n9290) );
  AND U13935 ( .A(p_input[5820]), .B(p_input[35820]), .Z(n9289) );
  AND U13936 ( .A(n9291), .B(n9292), .Z(o[581]) );
  AND U13937 ( .A(p_input[20581]), .B(p_input[10581]), .Z(n9292) );
  AND U13938 ( .A(p_input[581]), .B(p_input[30581]), .Z(n9291) );
  AND U13939 ( .A(n9293), .B(n9294), .Z(o[5819]) );
  AND U13940 ( .A(p_input[25819]), .B(p_input[15819]), .Z(n9294) );
  AND U13941 ( .A(p_input[5819]), .B(p_input[35819]), .Z(n9293) );
  AND U13942 ( .A(n9295), .B(n9296), .Z(o[5818]) );
  AND U13943 ( .A(p_input[25818]), .B(p_input[15818]), .Z(n9296) );
  AND U13944 ( .A(p_input[5818]), .B(p_input[35818]), .Z(n9295) );
  AND U13945 ( .A(n9297), .B(n9298), .Z(o[5817]) );
  AND U13946 ( .A(p_input[25817]), .B(p_input[15817]), .Z(n9298) );
  AND U13947 ( .A(p_input[5817]), .B(p_input[35817]), .Z(n9297) );
  AND U13948 ( .A(n9299), .B(n9300), .Z(o[5816]) );
  AND U13949 ( .A(p_input[25816]), .B(p_input[15816]), .Z(n9300) );
  AND U13950 ( .A(p_input[5816]), .B(p_input[35816]), .Z(n9299) );
  AND U13951 ( .A(n9301), .B(n9302), .Z(o[5815]) );
  AND U13952 ( .A(p_input[25815]), .B(p_input[15815]), .Z(n9302) );
  AND U13953 ( .A(p_input[5815]), .B(p_input[35815]), .Z(n9301) );
  AND U13954 ( .A(n9303), .B(n9304), .Z(o[5814]) );
  AND U13955 ( .A(p_input[25814]), .B(p_input[15814]), .Z(n9304) );
  AND U13956 ( .A(p_input[5814]), .B(p_input[35814]), .Z(n9303) );
  AND U13957 ( .A(n9305), .B(n9306), .Z(o[5813]) );
  AND U13958 ( .A(p_input[25813]), .B(p_input[15813]), .Z(n9306) );
  AND U13959 ( .A(p_input[5813]), .B(p_input[35813]), .Z(n9305) );
  AND U13960 ( .A(n9307), .B(n9308), .Z(o[5812]) );
  AND U13961 ( .A(p_input[25812]), .B(p_input[15812]), .Z(n9308) );
  AND U13962 ( .A(p_input[5812]), .B(p_input[35812]), .Z(n9307) );
  AND U13963 ( .A(n9309), .B(n9310), .Z(o[5811]) );
  AND U13964 ( .A(p_input[25811]), .B(p_input[15811]), .Z(n9310) );
  AND U13965 ( .A(p_input[5811]), .B(p_input[35811]), .Z(n9309) );
  AND U13966 ( .A(n9311), .B(n9312), .Z(o[5810]) );
  AND U13967 ( .A(p_input[25810]), .B(p_input[15810]), .Z(n9312) );
  AND U13968 ( .A(p_input[5810]), .B(p_input[35810]), .Z(n9311) );
  AND U13969 ( .A(n9313), .B(n9314), .Z(o[580]) );
  AND U13970 ( .A(p_input[20580]), .B(p_input[10580]), .Z(n9314) );
  AND U13971 ( .A(p_input[580]), .B(p_input[30580]), .Z(n9313) );
  AND U13972 ( .A(n9315), .B(n9316), .Z(o[5809]) );
  AND U13973 ( .A(p_input[25809]), .B(p_input[15809]), .Z(n9316) );
  AND U13974 ( .A(p_input[5809]), .B(p_input[35809]), .Z(n9315) );
  AND U13975 ( .A(n9317), .B(n9318), .Z(o[5808]) );
  AND U13976 ( .A(p_input[25808]), .B(p_input[15808]), .Z(n9318) );
  AND U13977 ( .A(p_input[5808]), .B(p_input[35808]), .Z(n9317) );
  AND U13978 ( .A(n9319), .B(n9320), .Z(o[5807]) );
  AND U13979 ( .A(p_input[25807]), .B(p_input[15807]), .Z(n9320) );
  AND U13980 ( .A(p_input[5807]), .B(p_input[35807]), .Z(n9319) );
  AND U13981 ( .A(n9321), .B(n9322), .Z(o[5806]) );
  AND U13982 ( .A(p_input[25806]), .B(p_input[15806]), .Z(n9322) );
  AND U13983 ( .A(p_input[5806]), .B(p_input[35806]), .Z(n9321) );
  AND U13984 ( .A(n9323), .B(n9324), .Z(o[5805]) );
  AND U13985 ( .A(p_input[25805]), .B(p_input[15805]), .Z(n9324) );
  AND U13986 ( .A(p_input[5805]), .B(p_input[35805]), .Z(n9323) );
  AND U13987 ( .A(n9325), .B(n9326), .Z(o[5804]) );
  AND U13988 ( .A(p_input[25804]), .B(p_input[15804]), .Z(n9326) );
  AND U13989 ( .A(p_input[5804]), .B(p_input[35804]), .Z(n9325) );
  AND U13990 ( .A(n9327), .B(n9328), .Z(o[5803]) );
  AND U13991 ( .A(p_input[25803]), .B(p_input[15803]), .Z(n9328) );
  AND U13992 ( .A(p_input[5803]), .B(p_input[35803]), .Z(n9327) );
  AND U13993 ( .A(n9329), .B(n9330), .Z(o[5802]) );
  AND U13994 ( .A(p_input[25802]), .B(p_input[15802]), .Z(n9330) );
  AND U13995 ( .A(p_input[5802]), .B(p_input[35802]), .Z(n9329) );
  AND U13996 ( .A(n9331), .B(n9332), .Z(o[5801]) );
  AND U13997 ( .A(p_input[25801]), .B(p_input[15801]), .Z(n9332) );
  AND U13998 ( .A(p_input[5801]), .B(p_input[35801]), .Z(n9331) );
  AND U13999 ( .A(n9333), .B(n9334), .Z(o[5800]) );
  AND U14000 ( .A(p_input[25800]), .B(p_input[15800]), .Z(n9334) );
  AND U14001 ( .A(p_input[5800]), .B(p_input[35800]), .Z(n9333) );
  AND U14002 ( .A(n9335), .B(n9336), .Z(o[57]) );
  AND U14003 ( .A(p_input[20057]), .B(p_input[10057]), .Z(n9336) );
  AND U14004 ( .A(p_input[57]), .B(p_input[30057]), .Z(n9335) );
  AND U14005 ( .A(n9337), .B(n9338), .Z(o[579]) );
  AND U14006 ( .A(p_input[20579]), .B(p_input[10579]), .Z(n9338) );
  AND U14007 ( .A(p_input[579]), .B(p_input[30579]), .Z(n9337) );
  AND U14008 ( .A(n9339), .B(n9340), .Z(o[5799]) );
  AND U14009 ( .A(p_input[25799]), .B(p_input[15799]), .Z(n9340) );
  AND U14010 ( .A(p_input[5799]), .B(p_input[35799]), .Z(n9339) );
  AND U14011 ( .A(n9341), .B(n9342), .Z(o[5798]) );
  AND U14012 ( .A(p_input[25798]), .B(p_input[15798]), .Z(n9342) );
  AND U14013 ( .A(p_input[5798]), .B(p_input[35798]), .Z(n9341) );
  AND U14014 ( .A(n9343), .B(n9344), .Z(o[5797]) );
  AND U14015 ( .A(p_input[25797]), .B(p_input[15797]), .Z(n9344) );
  AND U14016 ( .A(p_input[5797]), .B(p_input[35797]), .Z(n9343) );
  AND U14017 ( .A(n9345), .B(n9346), .Z(o[5796]) );
  AND U14018 ( .A(p_input[25796]), .B(p_input[15796]), .Z(n9346) );
  AND U14019 ( .A(p_input[5796]), .B(p_input[35796]), .Z(n9345) );
  AND U14020 ( .A(n9347), .B(n9348), .Z(o[5795]) );
  AND U14021 ( .A(p_input[25795]), .B(p_input[15795]), .Z(n9348) );
  AND U14022 ( .A(p_input[5795]), .B(p_input[35795]), .Z(n9347) );
  AND U14023 ( .A(n9349), .B(n9350), .Z(o[5794]) );
  AND U14024 ( .A(p_input[25794]), .B(p_input[15794]), .Z(n9350) );
  AND U14025 ( .A(p_input[5794]), .B(p_input[35794]), .Z(n9349) );
  AND U14026 ( .A(n9351), .B(n9352), .Z(o[5793]) );
  AND U14027 ( .A(p_input[25793]), .B(p_input[15793]), .Z(n9352) );
  AND U14028 ( .A(p_input[5793]), .B(p_input[35793]), .Z(n9351) );
  AND U14029 ( .A(n9353), .B(n9354), .Z(o[5792]) );
  AND U14030 ( .A(p_input[25792]), .B(p_input[15792]), .Z(n9354) );
  AND U14031 ( .A(p_input[5792]), .B(p_input[35792]), .Z(n9353) );
  AND U14032 ( .A(n9355), .B(n9356), .Z(o[5791]) );
  AND U14033 ( .A(p_input[25791]), .B(p_input[15791]), .Z(n9356) );
  AND U14034 ( .A(p_input[5791]), .B(p_input[35791]), .Z(n9355) );
  AND U14035 ( .A(n9357), .B(n9358), .Z(o[5790]) );
  AND U14036 ( .A(p_input[25790]), .B(p_input[15790]), .Z(n9358) );
  AND U14037 ( .A(p_input[5790]), .B(p_input[35790]), .Z(n9357) );
  AND U14038 ( .A(n9359), .B(n9360), .Z(o[578]) );
  AND U14039 ( .A(p_input[20578]), .B(p_input[10578]), .Z(n9360) );
  AND U14040 ( .A(p_input[578]), .B(p_input[30578]), .Z(n9359) );
  AND U14041 ( .A(n9361), .B(n9362), .Z(o[5789]) );
  AND U14042 ( .A(p_input[25789]), .B(p_input[15789]), .Z(n9362) );
  AND U14043 ( .A(p_input[5789]), .B(p_input[35789]), .Z(n9361) );
  AND U14044 ( .A(n9363), .B(n9364), .Z(o[5788]) );
  AND U14045 ( .A(p_input[25788]), .B(p_input[15788]), .Z(n9364) );
  AND U14046 ( .A(p_input[5788]), .B(p_input[35788]), .Z(n9363) );
  AND U14047 ( .A(n9365), .B(n9366), .Z(o[5787]) );
  AND U14048 ( .A(p_input[25787]), .B(p_input[15787]), .Z(n9366) );
  AND U14049 ( .A(p_input[5787]), .B(p_input[35787]), .Z(n9365) );
  AND U14050 ( .A(n9367), .B(n9368), .Z(o[5786]) );
  AND U14051 ( .A(p_input[25786]), .B(p_input[15786]), .Z(n9368) );
  AND U14052 ( .A(p_input[5786]), .B(p_input[35786]), .Z(n9367) );
  AND U14053 ( .A(n9369), .B(n9370), .Z(o[5785]) );
  AND U14054 ( .A(p_input[25785]), .B(p_input[15785]), .Z(n9370) );
  AND U14055 ( .A(p_input[5785]), .B(p_input[35785]), .Z(n9369) );
  AND U14056 ( .A(n9371), .B(n9372), .Z(o[5784]) );
  AND U14057 ( .A(p_input[25784]), .B(p_input[15784]), .Z(n9372) );
  AND U14058 ( .A(p_input[5784]), .B(p_input[35784]), .Z(n9371) );
  AND U14059 ( .A(n9373), .B(n9374), .Z(o[5783]) );
  AND U14060 ( .A(p_input[25783]), .B(p_input[15783]), .Z(n9374) );
  AND U14061 ( .A(p_input[5783]), .B(p_input[35783]), .Z(n9373) );
  AND U14062 ( .A(n9375), .B(n9376), .Z(o[5782]) );
  AND U14063 ( .A(p_input[25782]), .B(p_input[15782]), .Z(n9376) );
  AND U14064 ( .A(p_input[5782]), .B(p_input[35782]), .Z(n9375) );
  AND U14065 ( .A(n9377), .B(n9378), .Z(o[5781]) );
  AND U14066 ( .A(p_input[25781]), .B(p_input[15781]), .Z(n9378) );
  AND U14067 ( .A(p_input[5781]), .B(p_input[35781]), .Z(n9377) );
  AND U14068 ( .A(n9379), .B(n9380), .Z(o[5780]) );
  AND U14069 ( .A(p_input[25780]), .B(p_input[15780]), .Z(n9380) );
  AND U14070 ( .A(p_input[5780]), .B(p_input[35780]), .Z(n9379) );
  AND U14071 ( .A(n9381), .B(n9382), .Z(o[577]) );
  AND U14072 ( .A(p_input[20577]), .B(p_input[10577]), .Z(n9382) );
  AND U14073 ( .A(p_input[577]), .B(p_input[30577]), .Z(n9381) );
  AND U14074 ( .A(n9383), .B(n9384), .Z(o[5779]) );
  AND U14075 ( .A(p_input[25779]), .B(p_input[15779]), .Z(n9384) );
  AND U14076 ( .A(p_input[5779]), .B(p_input[35779]), .Z(n9383) );
  AND U14077 ( .A(n9385), .B(n9386), .Z(o[5778]) );
  AND U14078 ( .A(p_input[25778]), .B(p_input[15778]), .Z(n9386) );
  AND U14079 ( .A(p_input[5778]), .B(p_input[35778]), .Z(n9385) );
  AND U14080 ( .A(n9387), .B(n9388), .Z(o[5777]) );
  AND U14081 ( .A(p_input[25777]), .B(p_input[15777]), .Z(n9388) );
  AND U14082 ( .A(p_input[5777]), .B(p_input[35777]), .Z(n9387) );
  AND U14083 ( .A(n9389), .B(n9390), .Z(o[5776]) );
  AND U14084 ( .A(p_input[25776]), .B(p_input[15776]), .Z(n9390) );
  AND U14085 ( .A(p_input[5776]), .B(p_input[35776]), .Z(n9389) );
  AND U14086 ( .A(n9391), .B(n9392), .Z(o[5775]) );
  AND U14087 ( .A(p_input[25775]), .B(p_input[15775]), .Z(n9392) );
  AND U14088 ( .A(p_input[5775]), .B(p_input[35775]), .Z(n9391) );
  AND U14089 ( .A(n9393), .B(n9394), .Z(o[5774]) );
  AND U14090 ( .A(p_input[25774]), .B(p_input[15774]), .Z(n9394) );
  AND U14091 ( .A(p_input[5774]), .B(p_input[35774]), .Z(n9393) );
  AND U14092 ( .A(n9395), .B(n9396), .Z(o[5773]) );
  AND U14093 ( .A(p_input[25773]), .B(p_input[15773]), .Z(n9396) );
  AND U14094 ( .A(p_input[5773]), .B(p_input[35773]), .Z(n9395) );
  AND U14095 ( .A(n9397), .B(n9398), .Z(o[5772]) );
  AND U14096 ( .A(p_input[25772]), .B(p_input[15772]), .Z(n9398) );
  AND U14097 ( .A(p_input[5772]), .B(p_input[35772]), .Z(n9397) );
  AND U14098 ( .A(n9399), .B(n9400), .Z(o[5771]) );
  AND U14099 ( .A(p_input[25771]), .B(p_input[15771]), .Z(n9400) );
  AND U14100 ( .A(p_input[5771]), .B(p_input[35771]), .Z(n9399) );
  AND U14101 ( .A(n9401), .B(n9402), .Z(o[5770]) );
  AND U14102 ( .A(p_input[25770]), .B(p_input[15770]), .Z(n9402) );
  AND U14103 ( .A(p_input[5770]), .B(p_input[35770]), .Z(n9401) );
  AND U14104 ( .A(n9403), .B(n9404), .Z(o[576]) );
  AND U14105 ( .A(p_input[20576]), .B(p_input[10576]), .Z(n9404) );
  AND U14106 ( .A(p_input[576]), .B(p_input[30576]), .Z(n9403) );
  AND U14107 ( .A(n9405), .B(n9406), .Z(o[5769]) );
  AND U14108 ( .A(p_input[25769]), .B(p_input[15769]), .Z(n9406) );
  AND U14109 ( .A(p_input[5769]), .B(p_input[35769]), .Z(n9405) );
  AND U14110 ( .A(n9407), .B(n9408), .Z(o[5768]) );
  AND U14111 ( .A(p_input[25768]), .B(p_input[15768]), .Z(n9408) );
  AND U14112 ( .A(p_input[5768]), .B(p_input[35768]), .Z(n9407) );
  AND U14113 ( .A(n9409), .B(n9410), .Z(o[5767]) );
  AND U14114 ( .A(p_input[25767]), .B(p_input[15767]), .Z(n9410) );
  AND U14115 ( .A(p_input[5767]), .B(p_input[35767]), .Z(n9409) );
  AND U14116 ( .A(n9411), .B(n9412), .Z(o[5766]) );
  AND U14117 ( .A(p_input[25766]), .B(p_input[15766]), .Z(n9412) );
  AND U14118 ( .A(p_input[5766]), .B(p_input[35766]), .Z(n9411) );
  AND U14119 ( .A(n9413), .B(n9414), .Z(o[5765]) );
  AND U14120 ( .A(p_input[25765]), .B(p_input[15765]), .Z(n9414) );
  AND U14121 ( .A(p_input[5765]), .B(p_input[35765]), .Z(n9413) );
  AND U14122 ( .A(n9415), .B(n9416), .Z(o[5764]) );
  AND U14123 ( .A(p_input[25764]), .B(p_input[15764]), .Z(n9416) );
  AND U14124 ( .A(p_input[5764]), .B(p_input[35764]), .Z(n9415) );
  AND U14125 ( .A(n9417), .B(n9418), .Z(o[5763]) );
  AND U14126 ( .A(p_input[25763]), .B(p_input[15763]), .Z(n9418) );
  AND U14127 ( .A(p_input[5763]), .B(p_input[35763]), .Z(n9417) );
  AND U14128 ( .A(n9419), .B(n9420), .Z(o[5762]) );
  AND U14129 ( .A(p_input[25762]), .B(p_input[15762]), .Z(n9420) );
  AND U14130 ( .A(p_input[5762]), .B(p_input[35762]), .Z(n9419) );
  AND U14131 ( .A(n9421), .B(n9422), .Z(o[5761]) );
  AND U14132 ( .A(p_input[25761]), .B(p_input[15761]), .Z(n9422) );
  AND U14133 ( .A(p_input[5761]), .B(p_input[35761]), .Z(n9421) );
  AND U14134 ( .A(n9423), .B(n9424), .Z(o[5760]) );
  AND U14135 ( .A(p_input[25760]), .B(p_input[15760]), .Z(n9424) );
  AND U14136 ( .A(p_input[5760]), .B(p_input[35760]), .Z(n9423) );
  AND U14137 ( .A(n9425), .B(n9426), .Z(o[575]) );
  AND U14138 ( .A(p_input[20575]), .B(p_input[10575]), .Z(n9426) );
  AND U14139 ( .A(p_input[575]), .B(p_input[30575]), .Z(n9425) );
  AND U14140 ( .A(n9427), .B(n9428), .Z(o[5759]) );
  AND U14141 ( .A(p_input[25759]), .B(p_input[15759]), .Z(n9428) );
  AND U14142 ( .A(p_input[5759]), .B(p_input[35759]), .Z(n9427) );
  AND U14143 ( .A(n9429), .B(n9430), .Z(o[5758]) );
  AND U14144 ( .A(p_input[25758]), .B(p_input[15758]), .Z(n9430) );
  AND U14145 ( .A(p_input[5758]), .B(p_input[35758]), .Z(n9429) );
  AND U14146 ( .A(n9431), .B(n9432), .Z(o[5757]) );
  AND U14147 ( .A(p_input[25757]), .B(p_input[15757]), .Z(n9432) );
  AND U14148 ( .A(p_input[5757]), .B(p_input[35757]), .Z(n9431) );
  AND U14149 ( .A(n9433), .B(n9434), .Z(o[5756]) );
  AND U14150 ( .A(p_input[25756]), .B(p_input[15756]), .Z(n9434) );
  AND U14151 ( .A(p_input[5756]), .B(p_input[35756]), .Z(n9433) );
  AND U14152 ( .A(n9435), .B(n9436), .Z(o[5755]) );
  AND U14153 ( .A(p_input[25755]), .B(p_input[15755]), .Z(n9436) );
  AND U14154 ( .A(p_input[5755]), .B(p_input[35755]), .Z(n9435) );
  AND U14155 ( .A(n9437), .B(n9438), .Z(o[5754]) );
  AND U14156 ( .A(p_input[25754]), .B(p_input[15754]), .Z(n9438) );
  AND U14157 ( .A(p_input[5754]), .B(p_input[35754]), .Z(n9437) );
  AND U14158 ( .A(n9439), .B(n9440), .Z(o[5753]) );
  AND U14159 ( .A(p_input[25753]), .B(p_input[15753]), .Z(n9440) );
  AND U14160 ( .A(p_input[5753]), .B(p_input[35753]), .Z(n9439) );
  AND U14161 ( .A(n9441), .B(n9442), .Z(o[5752]) );
  AND U14162 ( .A(p_input[25752]), .B(p_input[15752]), .Z(n9442) );
  AND U14163 ( .A(p_input[5752]), .B(p_input[35752]), .Z(n9441) );
  AND U14164 ( .A(n9443), .B(n9444), .Z(o[5751]) );
  AND U14165 ( .A(p_input[25751]), .B(p_input[15751]), .Z(n9444) );
  AND U14166 ( .A(p_input[5751]), .B(p_input[35751]), .Z(n9443) );
  AND U14167 ( .A(n9445), .B(n9446), .Z(o[5750]) );
  AND U14168 ( .A(p_input[25750]), .B(p_input[15750]), .Z(n9446) );
  AND U14169 ( .A(p_input[5750]), .B(p_input[35750]), .Z(n9445) );
  AND U14170 ( .A(n9447), .B(n9448), .Z(o[574]) );
  AND U14171 ( .A(p_input[20574]), .B(p_input[10574]), .Z(n9448) );
  AND U14172 ( .A(p_input[574]), .B(p_input[30574]), .Z(n9447) );
  AND U14173 ( .A(n9449), .B(n9450), .Z(o[5749]) );
  AND U14174 ( .A(p_input[25749]), .B(p_input[15749]), .Z(n9450) );
  AND U14175 ( .A(p_input[5749]), .B(p_input[35749]), .Z(n9449) );
  AND U14176 ( .A(n9451), .B(n9452), .Z(o[5748]) );
  AND U14177 ( .A(p_input[25748]), .B(p_input[15748]), .Z(n9452) );
  AND U14178 ( .A(p_input[5748]), .B(p_input[35748]), .Z(n9451) );
  AND U14179 ( .A(n9453), .B(n9454), .Z(o[5747]) );
  AND U14180 ( .A(p_input[25747]), .B(p_input[15747]), .Z(n9454) );
  AND U14181 ( .A(p_input[5747]), .B(p_input[35747]), .Z(n9453) );
  AND U14182 ( .A(n9455), .B(n9456), .Z(o[5746]) );
  AND U14183 ( .A(p_input[25746]), .B(p_input[15746]), .Z(n9456) );
  AND U14184 ( .A(p_input[5746]), .B(p_input[35746]), .Z(n9455) );
  AND U14185 ( .A(n9457), .B(n9458), .Z(o[5745]) );
  AND U14186 ( .A(p_input[25745]), .B(p_input[15745]), .Z(n9458) );
  AND U14187 ( .A(p_input[5745]), .B(p_input[35745]), .Z(n9457) );
  AND U14188 ( .A(n9459), .B(n9460), .Z(o[5744]) );
  AND U14189 ( .A(p_input[25744]), .B(p_input[15744]), .Z(n9460) );
  AND U14190 ( .A(p_input[5744]), .B(p_input[35744]), .Z(n9459) );
  AND U14191 ( .A(n9461), .B(n9462), .Z(o[5743]) );
  AND U14192 ( .A(p_input[25743]), .B(p_input[15743]), .Z(n9462) );
  AND U14193 ( .A(p_input[5743]), .B(p_input[35743]), .Z(n9461) );
  AND U14194 ( .A(n9463), .B(n9464), .Z(o[5742]) );
  AND U14195 ( .A(p_input[25742]), .B(p_input[15742]), .Z(n9464) );
  AND U14196 ( .A(p_input[5742]), .B(p_input[35742]), .Z(n9463) );
  AND U14197 ( .A(n9465), .B(n9466), .Z(o[5741]) );
  AND U14198 ( .A(p_input[25741]), .B(p_input[15741]), .Z(n9466) );
  AND U14199 ( .A(p_input[5741]), .B(p_input[35741]), .Z(n9465) );
  AND U14200 ( .A(n9467), .B(n9468), .Z(o[5740]) );
  AND U14201 ( .A(p_input[25740]), .B(p_input[15740]), .Z(n9468) );
  AND U14202 ( .A(p_input[5740]), .B(p_input[35740]), .Z(n9467) );
  AND U14203 ( .A(n9469), .B(n9470), .Z(o[573]) );
  AND U14204 ( .A(p_input[20573]), .B(p_input[10573]), .Z(n9470) );
  AND U14205 ( .A(p_input[573]), .B(p_input[30573]), .Z(n9469) );
  AND U14206 ( .A(n9471), .B(n9472), .Z(o[5739]) );
  AND U14207 ( .A(p_input[25739]), .B(p_input[15739]), .Z(n9472) );
  AND U14208 ( .A(p_input[5739]), .B(p_input[35739]), .Z(n9471) );
  AND U14209 ( .A(n9473), .B(n9474), .Z(o[5738]) );
  AND U14210 ( .A(p_input[25738]), .B(p_input[15738]), .Z(n9474) );
  AND U14211 ( .A(p_input[5738]), .B(p_input[35738]), .Z(n9473) );
  AND U14212 ( .A(n9475), .B(n9476), .Z(o[5737]) );
  AND U14213 ( .A(p_input[25737]), .B(p_input[15737]), .Z(n9476) );
  AND U14214 ( .A(p_input[5737]), .B(p_input[35737]), .Z(n9475) );
  AND U14215 ( .A(n9477), .B(n9478), .Z(o[5736]) );
  AND U14216 ( .A(p_input[25736]), .B(p_input[15736]), .Z(n9478) );
  AND U14217 ( .A(p_input[5736]), .B(p_input[35736]), .Z(n9477) );
  AND U14218 ( .A(n9479), .B(n9480), .Z(o[5735]) );
  AND U14219 ( .A(p_input[25735]), .B(p_input[15735]), .Z(n9480) );
  AND U14220 ( .A(p_input[5735]), .B(p_input[35735]), .Z(n9479) );
  AND U14221 ( .A(n9481), .B(n9482), .Z(o[5734]) );
  AND U14222 ( .A(p_input[25734]), .B(p_input[15734]), .Z(n9482) );
  AND U14223 ( .A(p_input[5734]), .B(p_input[35734]), .Z(n9481) );
  AND U14224 ( .A(n9483), .B(n9484), .Z(o[5733]) );
  AND U14225 ( .A(p_input[25733]), .B(p_input[15733]), .Z(n9484) );
  AND U14226 ( .A(p_input[5733]), .B(p_input[35733]), .Z(n9483) );
  AND U14227 ( .A(n9485), .B(n9486), .Z(o[5732]) );
  AND U14228 ( .A(p_input[25732]), .B(p_input[15732]), .Z(n9486) );
  AND U14229 ( .A(p_input[5732]), .B(p_input[35732]), .Z(n9485) );
  AND U14230 ( .A(n9487), .B(n9488), .Z(o[5731]) );
  AND U14231 ( .A(p_input[25731]), .B(p_input[15731]), .Z(n9488) );
  AND U14232 ( .A(p_input[5731]), .B(p_input[35731]), .Z(n9487) );
  AND U14233 ( .A(n9489), .B(n9490), .Z(o[5730]) );
  AND U14234 ( .A(p_input[25730]), .B(p_input[15730]), .Z(n9490) );
  AND U14235 ( .A(p_input[5730]), .B(p_input[35730]), .Z(n9489) );
  AND U14236 ( .A(n9491), .B(n9492), .Z(o[572]) );
  AND U14237 ( .A(p_input[20572]), .B(p_input[10572]), .Z(n9492) );
  AND U14238 ( .A(p_input[572]), .B(p_input[30572]), .Z(n9491) );
  AND U14239 ( .A(n9493), .B(n9494), .Z(o[5729]) );
  AND U14240 ( .A(p_input[25729]), .B(p_input[15729]), .Z(n9494) );
  AND U14241 ( .A(p_input[5729]), .B(p_input[35729]), .Z(n9493) );
  AND U14242 ( .A(n9495), .B(n9496), .Z(o[5728]) );
  AND U14243 ( .A(p_input[25728]), .B(p_input[15728]), .Z(n9496) );
  AND U14244 ( .A(p_input[5728]), .B(p_input[35728]), .Z(n9495) );
  AND U14245 ( .A(n9497), .B(n9498), .Z(o[5727]) );
  AND U14246 ( .A(p_input[25727]), .B(p_input[15727]), .Z(n9498) );
  AND U14247 ( .A(p_input[5727]), .B(p_input[35727]), .Z(n9497) );
  AND U14248 ( .A(n9499), .B(n9500), .Z(o[5726]) );
  AND U14249 ( .A(p_input[25726]), .B(p_input[15726]), .Z(n9500) );
  AND U14250 ( .A(p_input[5726]), .B(p_input[35726]), .Z(n9499) );
  AND U14251 ( .A(n9501), .B(n9502), .Z(o[5725]) );
  AND U14252 ( .A(p_input[25725]), .B(p_input[15725]), .Z(n9502) );
  AND U14253 ( .A(p_input[5725]), .B(p_input[35725]), .Z(n9501) );
  AND U14254 ( .A(n9503), .B(n9504), .Z(o[5724]) );
  AND U14255 ( .A(p_input[25724]), .B(p_input[15724]), .Z(n9504) );
  AND U14256 ( .A(p_input[5724]), .B(p_input[35724]), .Z(n9503) );
  AND U14257 ( .A(n9505), .B(n9506), .Z(o[5723]) );
  AND U14258 ( .A(p_input[25723]), .B(p_input[15723]), .Z(n9506) );
  AND U14259 ( .A(p_input[5723]), .B(p_input[35723]), .Z(n9505) );
  AND U14260 ( .A(n9507), .B(n9508), .Z(o[5722]) );
  AND U14261 ( .A(p_input[25722]), .B(p_input[15722]), .Z(n9508) );
  AND U14262 ( .A(p_input[5722]), .B(p_input[35722]), .Z(n9507) );
  AND U14263 ( .A(n9509), .B(n9510), .Z(o[5721]) );
  AND U14264 ( .A(p_input[25721]), .B(p_input[15721]), .Z(n9510) );
  AND U14265 ( .A(p_input[5721]), .B(p_input[35721]), .Z(n9509) );
  AND U14266 ( .A(n9511), .B(n9512), .Z(o[5720]) );
  AND U14267 ( .A(p_input[25720]), .B(p_input[15720]), .Z(n9512) );
  AND U14268 ( .A(p_input[5720]), .B(p_input[35720]), .Z(n9511) );
  AND U14269 ( .A(n9513), .B(n9514), .Z(o[571]) );
  AND U14270 ( .A(p_input[20571]), .B(p_input[10571]), .Z(n9514) );
  AND U14271 ( .A(p_input[571]), .B(p_input[30571]), .Z(n9513) );
  AND U14272 ( .A(n9515), .B(n9516), .Z(o[5719]) );
  AND U14273 ( .A(p_input[25719]), .B(p_input[15719]), .Z(n9516) );
  AND U14274 ( .A(p_input[5719]), .B(p_input[35719]), .Z(n9515) );
  AND U14275 ( .A(n9517), .B(n9518), .Z(o[5718]) );
  AND U14276 ( .A(p_input[25718]), .B(p_input[15718]), .Z(n9518) );
  AND U14277 ( .A(p_input[5718]), .B(p_input[35718]), .Z(n9517) );
  AND U14278 ( .A(n9519), .B(n9520), .Z(o[5717]) );
  AND U14279 ( .A(p_input[25717]), .B(p_input[15717]), .Z(n9520) );
  AND U14280 ( .A(p_input[5717]), .B(p_input[35717]), .Z(n9519) );
  AND U14281 ( .A(n9521), .B(n9522), .Z(o[5716]) );
  AND U14282 ( .A(p_input[25716]), .B(p_input[15716]), .Z(n9522) );
  AND U14283 ( .A(p_input[5716]), .B(p_input[35716]), .Z(n9521) );
  AND U14284 ( .A(n9523), .B(n9524), .Z(o[5715]) );
  AND U14285 ( .A(p_input[25715]), .B(p_input[15715]), .Z(n9524) );
  AND U14286 ( .A(p_input[5715]), .B(p_input[35715]), .Z(n9523) );
  AND U14287 ( .A(n9525), .B(n9526), .Z(o[5714]) );
  AND U14288 ( .A(p_input[25714]), .B(p_input[15714]), .Z(n9526) );
  AND U14289 ( .A(p_input[5714]), .B(p_input[35714]), .Z(n9525) );
  AND U14290 ( .A(n9527), .B(n9528), .Z(o[5713]) );
  AND U14291 ( .A(p_input[25713]), .B(p_input[15713]), .Z(n9528) );
  AND U14292 ( .A(p_input[5713]), .B(p_input[35713]), .Z(n9527) );
  AND U14293 ( .A(n9529), .B(n9530), .Z(o[5712]) );
  AND U14294 ( .A(p_input[25712]), .B(p_input[15712]), .Z(n9530) );
  AND U14295 ( .A(p_input[5712]), .B(p_input[35712]), .Z(n9529) );
  AND U14296 ( .A(n9531), .B(n9532), .Z(o[5711]) );
  AND U14297 ( .A(p_input[25711]), .B(p_input[15711]), .Z(n9532) );
  AND U14298 ( .A(p_input[5711]), .B(p_input[35711]), .Z(n9531) );
  AND U14299 ( .A(n9533), .B(n9534), .Z(o[5710]) );
  AND U14300 ( .A(p_input[25710]), .B(p_input[15710]), .Z(n9534) );
  AND U14301 ( .A(p_input[5710]), .B(p_input[35710]), .Z(n9533) );
  AND U14302 ( .A(n9535), .B(n9536), .Z(o[570]) );
  AND U14303 ( .A(p_input[20570]), .B(p_input[10570]), .Z(n9536) );
  AND U14304 ( .A(p_input[570]), .B(p_input[30570]), .Z(n9535) );
  AND U14305 ( .A(n9537), .B(n9538), .Z(o[5709]) );
  AND U14306 ( .A(p_input[25709]), .B(p_input[15709]), .Z(n9538) );
  AND U14307 ( .A(p_input[5709]), .B(p_input[35709]), .Z(n9537) );
  AND U14308 ( .A(n9539), .B(n9540), .Z(o[5708]) );
  AND U14309 ( .A(p_input[25708]), .B(p_input[15708]), .Z(n9540) );
  AND U14310 ( .A(p_input[5708]), .B(p_input[35708]), .Z(n9539) );
  AND U14311 ( .A(n9541), .B(n9542), .Z(o[5707]) );
  AND U14312 ( .A(p_input[25707]), .B(p_input[15707]), .Z(n9542) );
  AND U14313 ( .A(p_input[5707]), .B(p_input[35707]), .Z(n9541) );
  AND U14314 ( .A(n9543), .B(n9544), .Z(o[5706]) );
  AND U14315 ( .A(p_input[25706]), .B(p_input[15706]), .Z(n9544) );
  AND U14316 ( .A(p_input[5706]), .B(p_input[35706]), .Z(n9543) );
  AND U14317 ( .A(n9545), .B(n9546), .Z(o[5705]) );
  AND U14318 ( .A(p_input[25705]), .B(p_input[15705]), .Z(n9546) );
  AND U14319 ( .A(p_input[5705]), .B(p_input[35705]), .Z(n9545) );
  AND U14320 ( .A(n9547), .B(n9548), .Z(o[5704]) );
  AND U14321 ( .A(p_input[25704]), .B(p_input[15704]), .Z(n9548) );
  AND U14322 ( .A(p_input[5704]), .B(p_input[35704]), .Z(n9547) );
  AND U14323 ( .A(n9549), .B(n9550), .Z(o[5703]) );
  AND U14324 ( .A(p_input[25703]), .B(p_input[15703]), .Z(n9550) );
  AND U14325 ( .A(p_input[5703]), .B(p_input[35703]), .Z(n9549) );
  AND U14326 ( .A(n9551), .B(n9552), .Z(o[5702]) );
  AND U14327 ( .A(p_input[25702]), .B(p_input[15702]), .Z(n9552) );
  AND U14328 ( .A(p_input[5702]), .B(p_input[35702]), .Z(n9551) );
  AND U14329 ( .A(n9553), .B(n9554), .Z(o[5701]) );
  AND U14330 ( .A(p_input[25701]), .B(p_input[15701]), .Z(n9554) );
  AND U14331 ( .A(p_input[5701]), .B(p_input[35701]), .Z(n9553) );
  AND U14332 ( .A(n9555), .B(n9556), .Z(o[5700]) );
  AND U14333 ( .A(p_input[25700]), .B(p_input[15700]), .Z(n9556) );
  AND U14334 ( .A(p_input[5700]), .B(p_input[35700]), .Z(n9555) );
  AND U14335 ( .A(n9557), .B(n9558), .Z(o[56]) );
  AND U14336 ( .A(p_input[20056]), .B(p_input[10056]), .Z(n9558) );
  AND U14337 ( .A(p_input[56]), .B(p_input[30056]), .Z(n9557) );
  AND U14338 ( .A(n9559), .B(n9560), .Z(o[569]) );
  AND U14339 ( .A(p_input[20569]), .B(p_input[10569]), .Z(n9560) );
  AND U14340 ( .A(p_input[569]), .B(p_input[30569]), .Z(n9559) );
  AND U14341 ( .A(n9561), .B(n9562), .Z(o[5699]) );
  AND U14342 ( .A(p_input[25699]), .B(p_input[15699]), .Z(n9562) );
  AND U14343 ( .A(p_input[5699]), .B(p_input[35699]), .Z(n9561) );
  AND U14344 ( .A(n9563), .B(n9564), .Z(o[5698]) );
  AND U14345 ( .A(p_input[25698]), .B(p_input[15698]), .Z(n9564) );
  AND U14346 ( .A(p_input[5698]), .B(p_input[35698]), .Z(n9563) );
  AND U14347 ( .A(n9565), .B(n9566), .Z(o[5697]) );
  AND U14348 ( .A(p_input[25697]), .B(p_input[15697]), .Z(n9566) );
  AND U14349 ( .A(p_input[5697]), .B(p_input[35697]), .Z(n9565) );
  AND U14350 ( .A(n9567), .B(n9568), .Z(o[5696]) );
  AND U14351 ( .A(p_input[25696]), .B(p_input[15696]), .Z(n9568) );
  AND U14352 ( .A(p_input[5696]), .B(p_input[35696]), .Z(n9567) );
  AND U14353 ( .A(n9569), .B(n9570), .Z(o[5695]) );
  AND U14354 ( .A(p_input[25695]), .B(p_input[15695]), .Z(n9570) );
  AND U14355 ( .A(p_input[5695]), .B(p_input[35695]), .Z(n9569) );
  AND U14356 ( .A(n9571), .B(n9572), .Z(o[5694]) );
  AND U14357 ( .A(p_input[25694]), .B(p_input[15694]), .Z(n9572) );
  AND U14358 ( .A(p_input[5694]), .B(p_input[35694]), .Z(n9571) );
  AND U14359 ( .A(n9573), .B(n9574), .Z(o[5693]) );
  AND U14360 ( .A(p_input[25693]), .B(p_input[15693]), .Z(n9574) );
  AND U14361 ( .A(p_input[5693]), .B(p_input[35693]), .Z(n9573) );
  AND U14362 ( .A(n9575), .B(n9576), .Z(o[5692]) );
  AND U14363 ( .A(p_input[25692]), .B(p_input[15692]), .Z(n9576) );
  AND U14364 ( .A(p_input[5692]), .B(p_input[35692]), .Z(n9575) );
  AND U14365 ( .A(n9577), .B(n9578), .Z(o[5691]) );
  AND U14366 ( .A(p_input[25691]), .B(p_input[15691]), .Z(n9578) );
  AND U14367 ( .A(p_input[5691]), .B(p_input[35691]), .Z(n9577) );
  AND U14368 ( .A(n9579), .B(n9580), .Z(o[5690]) );
  AND U14369 ( .A(p_input[25690]), .B(p_input[15690]), .Z(n9580) );
  AND U14370 ( .A(p_input[5690]), .B(p_input[35690]), .Z(n9579) );
  AND U14371 ( .A(n9581), .B(n9582), .Z(o[568]) );
  AND U14372 ( .A(p_input[20568]), .B(p_input[10568]), .Z(n9582) );
  AND U14373 ( .A(p_input[568]), .B(p_input[30568]), .Z(n9581) );
  AND U14374 ( .A(n9583), .B(n9584), .Z(o[5689]) );
  AND U14375 ( .A(p_input[25689]), .B(p_input[15689]), .Z(n9584) );
  AND U14376 ( .A(p_input[5689]), .B(p_input[35689]), .Z(n9583) );
  AND U14377 ( .A(n9585), .B(n9586), .Z(o[5688]) );
  AND U14378 ( .A(p_input[25688]), .B(p_input[15688]), .Z(n9586) );
  AND U14379 ( .A(p_input[5688]), .B(p_input[35688]), .Z(n9585) );
  AND U14380 ( .A(n9587), .B(n9588), .Z(o[5687]) );
  AND U14381 ( .A(p_input[25687]), .B(p_input[15687]), .Z(n9588) );
  AND U14382 ( .A(p_input[5687]), .B(p_input[35687]), .Z(n9587) );
  AND U14383 ( .A(n9589), .B(n9590), .Z(o[5686]) );
  AND U14384 ( .A(p_input[25686]), .B(p_input[15686]), .Z(n9590) );
  AND U14385 ( .A(p_input[5686]), .B(p_input[35686]), .Z(n9589) );
  AND U14386 ( .A(n9591), .B(n9592), .Z(o[5685]) );
  AND U14387 ( .A(p_input[25685]), .B(p_input[15685]), .Z(n9592) );
  AND U14388 ( .A(p_input[5685]), .B(p_input[35685]), .Z(n9591) );
  AND U14389 ( .A(n9593), .B(n9594), .Z(o[5684]) );
  AND U14390 ( .A(p_input[25684]), .B(p_input[15684]), .Z(n9594) );
  AND U14391 ( .A(p_input[5684]), .B(p_input[35684]), .Z(n9593) );
  AND U14392 ( .A(n9595), .B(n9596), .Z(o[5683]) );
  AND U14393 ( .A(p_input[25683]), .B(p_input[15683]), .Z(n9596) );
  AND U14394 ( .A(p_input[5683]), .B(p_input[35683]), .Z(n9595) );
  AND U14395 ( .A(n9597), .B(n9598), .Z(o[5682]) );
  AND U14396 ( .A(p_input[25682]), .B(p_input[15682]), .Z(n9598) );
  AND U14397 ( .A(p_input[5682]), .B(p_input[35682]), .Z(n9597) );
  AND U14398 ( .A(n9599), .B(n9600), .Z(o[5681]) );
  AND U14399 ( .A(p_input[25681]), .B(p_input[15681]), .Z(n9600) );
  AND U14400 ( .A(p_input[5681]), .B(p_input[35681]), .Z(n9599) );
  AND U14401 ( .A(n9601), .B(n9602), .Z(o[5680]) );
  AND U14402 ( .A(p_input[25680]), .B(p_input[15680]), .Z(n9602) );
  AND U14403 ( .A(p_input[5680]), .B(p_input[35680]), .Z(n9601) );
  AND U14404 ( .A(n9603), .B(n9604), .Z(o[567]) );
  AND U14405 ( .A(p_input[20567]), .B(p_input[10567]), .Z(n9604) );
  AND U14406 ( .A(p_input[567]), .B(p_input[30567]), .Z(n9603) );
  AND U14407 ( .A(n9605), .B(n9606), .Z(o[5679]) );
  AND U14408 ( .A(p_input[25679]), .B(p_input[15679]), .Z(n9606) );
  AND U14409 ( .A(p_input[5679]), .B(p_input[35679]), .Z(n9605) );
  AND U14410 ( .A(n9607), .B(n9608), .Z(o[5678]) );
  AND U14411 ( .A(p_input[25678]), .B(p_input[15678]), .Z(n9608) );
  AND U14412 ( .A(p_input[5678]), .B(p_input[35678]), .Z(n9607) );
  AND U14413 ( .A(n9609), .B(n9610), .Z(o[5677]) );
  AND U14414 ( .A(p_input[25677]), .B(p_input[15677]), .Z(n9610) );
  AND U14415 ( .A(p_input[5677]), .B(p_input[35677]), .Z(n9609) );
  AND U14416 ( .A(n9611), .B(n9612), .Z(o[5676]) );
  AND U14417 ( .A(p_input[25676]), .B(p_input[15676]), .Z(n9612) );
  AND U14418 ( .A(p_input[5676]), .B(p_input[35676]), .Z(n9611) );
  AND U14419 ( .A(n9613), .B(n9614), .Z(o[5675]) );
  AND U14420 ( .A(p_input[25675]), .B(p_input[15675]), .Z(n9614) );
  AND U14421 ( .A(p_input[5675]), .B(p_input[35675]), .Z(n9613) );
  AND U14422 ( .A(n9615), .B(n9616), .Z(o[5674]) );
  AND U14423 ( .A(p_input[25674]), .B(p_input[15674]), .Z(n9616) );
  AND U14424 ( .A(p_input[5674]), .B(p_input[35674]), .Z(n9615) );
  AND U14425 ( .A(n9617), .B(n9618), .Z(o[5673]) );
  AND U14426 ( .A(p_input[25673]), .B(p_input[15673]), .Z(n9618) );
  AND U14427 ( .A(p_input[5673]), .B(p_input[35673]), .Z(n9617) );
  AND U14428 ( .A(n9619), .B(n9620), .Z(o[5672]) );
  AND U14429 ( .A(p_input[25672]), .B(p_input[15672]), .Z(n9620) );
  AND U14430 ( .A(p_input[5672]), .B(p_input[35672]), .Z(n9619) );
  AND U14431 ( .A(n9621), .B(n9622), .Z(o[5671]) );
  AND U14432 ( .A(p_input[25671]), .B(p_input[15671]), .Z(n9622) );
  AND U14433 ( .A(p_input[5671]), .B(p_input[35671]), .Z(n9621) );
  AND U14434 ( .A(n9623), .B(n9624), .Z(o[5670]) );
  AND U14435 ( .A(p_input[25670]), .B(p_input[15670]), .Z(n9624) );
  AND U14436 ( .A(p_input[5670]), .B(p_input[35670]), .Z(n9623) );
  AND U14437 ( .A(n9625), .B(n9626), .Z(o[566]) );
  AND U14438 ( .A(p_input[20566]), .B(p_input[10566]), .Z(n9626) );
  AND U14439 ( .A(p_input[566]), .B(p_input[30566]), .Z(n9625) );
  AND U14440 ( .A(n9627), .B(n9628), .Z(o[5669]) );
  AND U14441 ( .A(p_input[25669]), .B(p_input[15669]), .Z(n9628) );
  AND U14442 ( .A(p_input[5669]), .B(p_input[35669]), .Z(n9627) );
  AND U14443 ( .A(n9629), .B(n9630), .Z(o[5668]) );
  AND U14444 ( .A(p_input[25668]), .B(p_input[15668]), .Z(n9630) );
  AND U14445 ( .A(p_input[5668]), .B(p_input[35668]), .Z(n9629) );
  AND U14446 ( .A(n9631), .B(n9632), .Z(o[5667]) );
  AND U14447 ( .A(p_input[25667]), .B(p_input[15667]), .Z(n9632) );
  AND U14448 ( .A(p_input[5667]), .B(p_input[35667]), .Z(n9631) );
  AND U14449 ( .A(n9633), .B(n9634), .Z(o[5666]) );
  AND U14450 ( .A(p_input[25666]), .B(p_input[15666]), .Z(n9634) );
  AND U14451 ( .A(p_input[5666]), .B(p_input[35666]), .Z(n9633) );
  AND U14452 ( .A(n9635), .B(n9636), .Z(o[5665]) );
  AND U14453 ( .A(p_input[25665]), .B(p_input[15665]), .Z(n9636) );
  AND U14454 ( .A(p_input[5665]), .B(p_input[35665]), .Z(n9635) );
  AND U14455 ( .A(n9637), .B(n9638), .Z(o[5664]) );
  AND U14456 ( .A(p_input[25664]), .B(p_input[15664]), .Z(n9638) );
  AND U14457 ( .A(p_input[5664]), .B(p_input[35664]), .Z(n9637) );
  AND U14458 ( .A(n9639), .B(n9640), .Z(o[5663]) );
  AND U14459 ( .A(p_input[25663]), .B(p_input[15663]), .Z(n9640) );
  AND U14460 ( .A(p_input[5663]), .B(p_input[35663]), .Z(n9639) );
  AND U14461 ( .A(n9641), .B(n9642), .Z(o[5662]) );
  AND U14462 ( .A(p_input[25662]), .B(p_input[15662]), .Z(n9642) );
  AND U14463 ( .A(p_input[5662]), .B(p_input[35662]), .Z(n9641) );
  AND U14464 ( .A(n9643), .B(n9644), .Z(o[5661]) );
  AND U14465 ( .A(p_input[25661]), .B(p_input[15661]), .Z(n9644) );
  AND U14466 ( .A(p_input[5661]), .B(p_input[35661]), .Z(n9643) );
  AND U14467 ( .A(n9645), .B(n9646), .Z(o[5660]) );
  AND U14468 ( .A(p_input[25660]), .B(p_input[15660]), .Z(n9646) );
  AND U14469 ( .A(p_input[5660]), .B(p_input[35660]), .Z(n9645) );
  AND U14470 ( .A(n9647), .B(n9648), .Z(o[565]) );
  AND U14471 ( .A(p_input[20565]), .B(p_input[10565]), .Z(n9648) );
  AND U14472 ( .A(p_input[565]), .B(p_input[30565]), .Z(n9647) );
  AND U14473 ( .A(n9649), .B(n9650), .Z(o[5659]) );
  AND U14474 ( .A(p_input[25659]), .B(p_input[15659]), .Z(n9650) );
  AND U14475 ( .A(p_input[5659]), .B(p_input[35659]), .Z(n9649) );
  AND U14476 ( .A(n9651), .B(n9652), .Z(o[5658]) );
  AND U14477 ( .A(p_input[25658]), .B(p_input[15658]), .Z(n9652) );
  AND U14478 ( .A(p_input[5658]), .B(p_input[35658]), .Z(n9651) );
  AND U14479 ( .A(n9653), .B(n9654), .Z(o[5657]) );
  AND U14480 ( .A(p_input[25657]), .B(p_input[15657]), .Z(n9654) );
  AND U14481 ( .A(p_input[5657]), .B(p_input[35657]), .Z(n9653) );
  AND U14482 ( .A(n9655), .B(n9656), .Z(o[5656]) );
  AND U14483 ( .A(p_input[25656]), .B(p_input[15656]), .Z(n9656) );
  AND U14484 ( .A(p_input[5656]), .B(p_input[35656]), .Z(n9655) );
  AND U14485 ( .A(n9657), .B(n9658), .Z(o[5655]) );
  AND U14486 ( .A(p_input[25655]), .B(p_input[15655]), .Z(n9658) );
  AND U14487 ( .A(p_input[5655]), .B(p_input[35655]), .Z(n9657) );
  AND U14488 ( .A(n9659), .B(n9660), .Z(o[5654]) );
  AND U14489 ( .A(p_input[25654]), .B(p_input[15654]), .Z(n9660) );
  AND U14490 ( .A(p_input[5654]), .B(p_input[35654]), .Z(n9659) );
  AND U14491 ( .A(n9661), .B(n9662), .Z(o[5653]) );
  AND U14492 ( .A(p_input[25653]), .B(p_input[15653]), .Z(n9662) );
  AND U14493 ( .A(p_input[5653]), .B(p_input[35653]), .Z(n9661) );
  AND U14494 ( .A(n9663), .B(n9664), .Z(o[5652]) );
  AND U14495 ( .A(p_input[25652]), .B(p_input[15652]), .Z(n9664) );
  AND U14496 ( .A(p_input[5652]), .B(p_input[35652]), .Z(n9663) );
  AND U14497 ( .A(n9665), .B(n9666), .Z(o[5651]) );
  AND U14498 ( .A(p_input[25651]), .B(p_input[15651]), .Z(n9666) );
  AND U14499 ( .A(p_input[5651]), .B(p_input[35651]), .Z(n9665) );
  AND U14500 ( .A(n9667), .B(n9668), .Z(o[5650]) );
  AND U14501 ( .A(p_input[25650]), .B(p_input[15650]), .Z(n9668) );
  AND U14502 ( .A(p_input[5650]), .B(p_input[35650]), .Z(n9667) );
  AND U14503 ( .A(n9669), .B(n9670), .Z(o[564]) );
  AND U14504 ( .A(p_input[20564]), .B(p_input[10564]), .Z(n9670) );
  AND U14505 ( .A(p_input[564]), .B(p_input[30564]), .Z(n9669) );
  AND U14506 ( .A(n9671), .B(n9672), .Z(o[5649]) );
  AND U14507 ( .A(p_input[25649]), .B(p_input[15649]), .Z(n9672) );
  AND U14508 ( .A(p_input[5649]), .B(p_input[35649]), .Z(n9671) );
  AND U14509 ( .A(n9673), .B(n9674), .Z(o[5648]) );
  AND U14510 ( .A(p_input[25648]), .B(p_input[15648]), .Z(n9674) );
  AND U14511 ( .A(p_input[5648]), .B(p_input[35648]), .Z(n9673) );
  AND U14512 ( .A(n9675), .B(n9676), .Z(o[5647]) );
  AND U14513 ( .A(p_input[25647]), .B(p_input[15647]), .Z(n9676) );
  AND U14514 ( .A(p_input[5647]), .B(p_input[35647]), .Z(n9675) );
  AND U14515 ( .A(n9677), .B(n9678), .Z(o[5646]) );
  AND U14516 ( .A(p_input[25646]), .B(p_input[15646]), .Z(n9678) );
  AND U14517 ( .A(p_input[5646]), .B(p_input[35646]), .Z(n9677) );
  AND U14518 ( .A(n9679), .B(n9680), .Z(o[5645]) );
  AND U14519 ( .A(p_input[25645]), .B(p_input[15645]), .Z(n9680) );
  AND U14520 ( .A(p_input[5645]), .B(p_input[35645]), .Z(n9679) );
  AND U14521 ( .A(n9681), .B(n9682), .Z(o[5644]) );
  AND U14522 ( .A(p_input[25644]), .B(p_input[15644]), .Z(n9682) );
  AND U14523 ( .A(p_input[5644]), .B(p_input[35644]), .Z(n9681) );
  AND U14524 ( .A(n9683), .B(n9684), .Z(o[5643]) );
  AND U14525 ( .A(p_input[25643]), .B(p_input[15643]), .Z(n9684) );
  AND U14526 ( .A(p_input[5643]), .B(p_input[35643]), .Z(n9683) );
  AND U14527 ( .A(n9685), .B(n9686), .Z(o[5642]) );
  AND U14528 ( .A(p_input[25642]), .B(p_input[15642]), .Z(n9686) );
  AND U14529 ( .A(p_input[5642]), .B(p_input[35642]), .Z(n9685) );
  AND U14530 ( .A(n9687), .B(n9688), .Z(o[5641]) );
  AND U14531 ( .A(p_input[25641]), .B(p_input[15641]), .Z(n9688) );
  AND U14532 ( .A(p_input[5641]), .B(p_input[35641]), .Z(n9687) );
  AND U14533 ( .A(n9689), .B(n9690), .Z(o[5640]) );
  AND U14534 ( .A(p_input[25640]), .B(p_input[15640]), .Z(n9690) );
  AND U14535 ( .A(p_input[5640]), .B(p_input[35640]), .Z(n9689) );
  AND U14536 ( .A(n9691), .B(n9692), .Z(o[563]) );
  AND U14537 ( .A(p_input[20563]), .B(p_input[10563]), .Z(n9692) );
  AND U14538 ( .A(p_input[563]), .B(p_input[30563]), .Z(n9691) );
  AND U14539 ( .A(n9693), .B(n9694), .Z(o[5639]) );
  AND U14540 ( .A(p_input[25639]), .B(p_input[15639]), .Z(n9694) );
  AND U14541 ( .A(p_input[5639]), .B(p_input[35639]), .Z(n9693) );
  AND U14542 ( .A(n9695), .B(n9696), .Z(o[5638]) );
  AND U14543 ( .A(p_input[25638]), .B(p_input[15638]), .Z(n9696) );
  AND U14544 ( .A(p_input[5638]), .B(p_input[35638]), .Z(n9695) );
  AND U14545 ( .A(n9697), .B(n9698), .Z(o[5637]) );
  AND U14546 ( .A(p_input[25637]), .B(p_input[15637]), .Z(n9698) );
  AND U14547 ( .A(p_input[5637]), .B(p_input[35637]), .Z(n9697) );
  AND U14548 ( .A(n9699), .B(n9700), .Z(o[5636]) );
  AND U14549 ( .A(p_input[25636]), .B(p_input[15636]), .Z(n9700) );
  AND U14550 ( .A(p_input[5636]), .B(p_input[35636]), .Z(n9699) );
  AND U14551 ( .A(n9701), .B(n9702), .Z(o[5635]) );
  AND U14552 ( .A(p_input[25635]), .B(p_input[15635]), .Z(n9702) );
  AND U14553 ( .A(p_input[5635]), .B(p_input[35635]), .Z(n9701) );
  AND U14554 ( .A(n9703), .B(n9704), .Z(o[5634]) );
  AND U14555 ( .A(p_input[25634]), .B(p_input[15634]), .Z(n9704) );
  AND U14556 ( .A(p_input[5634]), .B(p_input[35634]), .Z(n9703) );
  AND U14557 ( .A(n9705), .B(n9706), .Z(o[5633]) );
  AND U14558 ( .A(p_input[25633]), .B(p_input[15633]), .Z(n9706) );
  AND U14559 ( .A(p_input[5633]), .B(p_input[35633]), .Z(n9705) );
  AND U14560 ( .A(n9707), .B(n9708), .Z(o[5632]) );
  AND U14561 ( .A(p_input[25632]), .B(p_input[15632]), .Z(n9708) );
  AND U14562 ( .A(p_input[5632]), .B(p_input[35632]), .Z(n9707) );
  AND U14563 ( .A(n9709), .B(n9710), .Z(o[5631]) );
  AND U14564 ( .A(p_input[25631]), .B(p_input[15631]), .Z(n9710) );
  AND U14565 ( .A(p_input[5631]), .B(p_input[35631]), .Z(n9709) );
  AND U14566 ( .A(n9711), .B(n9712), .Z(o[5630]) );
  AND U14567 ( .A(p_input[25630]), .B(p_input[15630]), .Z(n9712) );
  AND U14568 ( .A(p_input[5630]), .B(p_input[35630]), .Z(n9711) );
  AND U14569 ( .A(n9713), .B(n9714), .Z(o[562]) );
  AND U14570 ( .A(p_input[20562]), .B(p_input[10562]), .Z(n9714) );
  AND U14571 ( .A(p_input[562]), .B(p_input[30562]), .Z(n9713) );
  AND U14572 ( .A(n9715), .B(n9716), .Z(o[5629]) );
  AND U14573 ( .A(p_input[25629]), .B(p_input[15629]), .Z(n9716) );
  AND U14574 ( .A(p_input[5629]), .B(p_input[35629]), .Z(n9715) );
  AND U14575 ( .A(n9717), .B(n9718), .Z(o[5628]) );
  AND U14576 ( .A(p_input[25628]), .B(p_input[15628]), .Z(n9718) );
  AND U14577 ( .A(p_input[5628]), .B(p_input[35628]), .Z(n9717) );
  AND U14578 ( .A(n9719), .B(n9720), .Z(o[5627]) );
  AND U14579 ( .A(p_input[25627]), .B(p_input[15627]), .Z(n9720) );
  AND U14580 ( .A(p_input[5627]), .B(p_input[35627]), .Z(n9719) );
  AND U14581 ( .A(n9721), .B(n9722), .Z(o[5626]) );
  AND U14582 ( .A(p_input[25626]), .B(p_input[15626]), .Z(n9722) );
  AND U14583 ( .A(p_input[5626]), .B(p_input[35626]), .Z(n9721) );
  AND U14584 ( .A(n9723), .B(n9724), .Z(o[5625]) );
  AND U14585 ( .A(p_input[25625]), .B(p_input[15625]), .Z(n9724) );
  AND U14586 ( .A(p_input[5625]), .B(p_input[35625]), .Z(n9723) );
  AND U14587 ( .A(n9725), .B(n9726), .Z(o[5624]) );
  AND U14588 ( .A(p_input[25624]), .B(p_input[15624]), .Z(n9726) );
  AND U14589 ( .A(p_input[5624]), .B(p_input[35624]), .Z(n9725) );
  AND U14590 ( .A(n9727), .B(n9728), .Z(o[5623]) );
  AND U14591 ( .A(p_input[25623]), .B(p_input[15623]), .Z(n9728) );
  AND U14592 ( .A(p_input[5623]), .B(p_input[35623]), .Z(n9727) );
  AND U14593 ( .A(n9729), .B(n9730), .Z(o[5622]) );
  AND U14594 ( .A(p_input[25622]), .B(p_input[15622]), .Z(n9730) );
  AND U14595 ( .A(p_input[5622]), .B(p_input[35622]), .Z(n9729) );
  AND U14596 ( .A(n9731), .B(n9732), .Z(o[5621]) );
  AND U14597 ( .A(p_input[25621]), .B(p_input[15621]), .Z(n9732) );
  AND U14598 ( .A(p_input[5621]), .B(p_input[35621]), .Z(n9731) );
  AND U14599 ( .A(n9733), .B(n9734), .Z(o[5620]) );
  AND U14600 ( .A(p_input[25620]), .B(p_input[15620]), .Z(n9734) );
  AND U14601 ( .A(p_input[5620]), .B(p_input[35620]), .Z(n9733) );
  AND U14602 ( .A(n9735), .B(n9736), .Z(o[561]) );
  AND U14603 ( .A(p_input[20561]), .B(p_input[10561]), .Z(n9736) );
  AND U14604 ( .A(p_input[561]), .B(p_input[30561]), .Z(n9735) );
  AND U14605 ( .A(n9737), .B(n9738), .Z(o[5619]) );
  AND U14606 ( .A(p_input[25619]), .B(p_input[15619]), .Z(n9738) );
  AND U14607 ( .A(p_input[5619]), .B(p_input[35619]), .Z(n9737) );
  AND U14608 ( .A(n9739), .B(n9740), .Z(o[5618]) );
  AND U14609 ( .A(p_input[25618]), .B(p_input[15618]), .Z(n9740) );
  AND U14610 ( .A(p_input[5618]), .B(p_input[35618]), .Z(n9739) );
  AND U14611 ( .A(n9741), .B(n9742), .Z(o[5617]) );
  AND U14612 ( .A(p_input[25617]), .B(p_input[15617]), .Z(n9742) );
  AND U14613 ( .A(p_input[5617]), .B(p_input[35617]), .Z(n9741) );
  AND U14614 ( .A(n9743), .B(n9744), .Z(o[5616]) );
  AND U14615 ( .A(p_input[25616]), .B(p_input[15616]), .Z(n9744) );
  AND U14616 ( .A(p_input[5616]), .B(p_input[35616]), .Z(n9743) );
  AND U14617 ( .A(n9745), .B(n9746), .Z(o[5615]) );
  AND U14618 ( .A(p_input[25615]), .B(p_input[15615]), .Z(n9746) );
  AND U14619 ( .A(p_input[5615]), .B(p_input[35615]), .Z(n9745) );
  AND U14620 ( .A(n9747), .B(n9748), .Z(o[5614]) );
  AND U14621 ( .A(p_input[25614]), .B(p_input[15614]), .Z(n9748) );
  AND U14622 ( .A(p_input[5614]), .B(p_input[35614]), .Z(n9747) );
  AND U14623 ( .A(n9749), .B(n9750), .Z(o[5613]) );
  AND U14624 ( .A(p_input[25613]), .B(p_input[15613]), .Z(n9750) );
  AND U14625 ( .A(p_input[5613]), .B(p_input[35613]), .Z(n9749) );
  AND U14626 ( .A(n9751), .B(n9752), .Z(o[5612]) );
  AND U14627 ( .A(p_input[25612]), .B(p_input[15612]), .Z(n9752) );
  AND U14628 ( .A(p_input[5612]), .B(p_input[35612]), .Z(n9751) );
  AND U14629 ( .A(n9753), .B(n9754), .Z(o[5611]) );
  AND U14630 ( .A(p_input[25611]), .B(p_input[15611]), .Z(n9754) );
  AND U14631 ( .A(p_input[5611]), .B(p_input[35611]), .Z(n9753) );
  AND U14632 ( .A(n9755), .B(n9756), .Z(o[5610]) );
  AND U14633 ( .A(p_input[25610]), .B(p_input[15610]), .Z(n9756) );
  AND U14634 ( .A(p_input[5610]), .B(p_input[35610]), .Z(n9755) );
  AND U14635 ( .A(n9757), .B(n9758), .Z(o[560]) );
  AND U14636 ( .A(p_input[20560]), .B(p_input[10560]), .Z(n9758) );
  AND U14637 ( .A(p_input[560]), .B(p_input[30560]), .Z(n9757) );
  AND U14638 ( .A(n9759), .B(n9760), .Z(o[5609]) );
  AND U14639 ( .A(p_input[25609]), .B(p_input[15609]), .Z(n9760) );
  AND U14640 ( .A(p_input[5609]), .B(p_input[35609]), .Z(n9759) );
  AND U14641 ( .A(n9761), .B(n9762), .Z(o[5608]) );
  AND U14642 ( .A(p_input[25608]), .B(p_input[15608]), .Z(n9762) );
  AND U14643 ( .A(p_input[5608]), .B(p_input[35608]), .Z(n9761) );
  AND U14644 ( .A(n9763), .B(n9764), .Z(o[5607]) );
  AND U14645 ( .A(p_input[25607]), .B(p_input[15607]), .Z(n9764) );
  AND U14646 ( .A(p_input[5607]), .B(p_input[35607]), .Z(n9763) );
  AND U14647 ( .A(n9765), .B(n9766), .Z(o[5606]) );
  AND U14648 ( .A(p_input[25606]), .B(p_input[15606]), .Z(n9766) );
  AND U14649 ( .A(p_input[5606]), .B(p_input[35606]), .Z(n9765) );
  AND U14650 ( .A(n9767), .B(n9768), .Z(o[5605]) );
  AND U14651 ( .A(p_input[25605]), .B(p_input[15605]), .Z(n9768) );
  AND U14652 ( .A(p_input[5605]), .B(p_input[35605]), .Z(n9767) );
  AND U14653 ( .A(n9769), .B(n9770), .Z(o[5604]) );
  AND U14654 ( .A(p_input[25604]), .B(p_input[15604]), .Z(n9770) );
  AND U14655 ( .A(p_input[5604]), .B(p_input[35604]), .Z(n9769) );
  AND U14656 ( .A(n9771), .B(n9772), .Z(o[5603]) );
  AND U14657 ( .A(p_input[25603]), .B(p_input[15603]), .Z(n9772) );
  AND U14658 ( .A(p_input[5603]), .B(p_input[35603]), .Z(n9771) );
  AND U14659 ( .A(n9773), .B(n9774), .Z(o[5602]) );
  AND U14660 ( .A(p_input[25602]), .B(p_input[15602]), .Z(n9774) );
  AND U14661 ( .A(p_input[5602]), .B(p_input[35602]), .Z(n9773) );
  AND U14662 ( .A(n9775), .B(n9776), .Z(o[5601]) );
  AND U14663 ( .A(p_input[25601]), .B(p_input[15601]), .Z(n9776) );
  AND U14664 ( .A(p_input[5601]), .B(p_input[35601]), .Z(n9775) );
  AND U14665 ( .A(n9777), .B(n9778), .Z(o[5600]) );
  AND U14666 ( .A(p_input[25600]), .B(p_input[15600]), .Z(n9778) );
  AND U14667 ( .A(p_input[5600]), .B(p_input[35600]), .Z(n9777) );
  AND U14668 ( .A(n9779), .B(n9780), .Z(o[55]) );
  AND U14669 ( .A(p_input[20055]), .B(p_input[10055]), .Z(n9780) );
  AND U14670 ( .A(p_input[55]), .B(p_input[30055]), .Z(n9779) );
  AND U14671 ( .A(n9781), .B(n9782), .Z(o[559]) );
  AND U14672 ( .A(p_input[20559]), .B(p_input[10559]), .Z(n9782) );
  AND U14673 ( .A(p_input[559]), .B(p_input[30559]), .Z(n9781) );
  AND U14674 ( .A(n9783), .B(n9784), .Z(o[5599]) );
  AND U14675 ( .A(p_input[25599]), .B(p_input[15599]), .Z(n9784) );
  AND U14676 ( .A(p_input[5599]), .B(p_input[35599]), .Z(n9783) );
  AND U14677 ( .A(n9785), .B(n9786), .Z(o[5598]) );
  AND U14678 ( .A(p_input[25598]), .B(p_input[15598]), .Z(n9786) );
  AND U14679 ( .A(p_input[5598]), .B(p_input[35598]), .Z(n9785) );
  AND U14680 ( .A(n9787), .B(n9788), .Z(o[5597]) );
  AND U14681 ( .A(p_input[25597]), .B(p_input[15597]), .Z(n9788) );
  AND U14682 ( .A(p_input[5597]), .B(p_input[35597]), .Z(n9787) );
  AND U14683 ( .A(n9789), .B(n9790), .Z(o[5596]) );
  AND U14684 ( .A(p_input[25596]), .B(p_input[15596]), .Z(n9790) );
  AND U14685 ( .A(p_input[5596]), .B(p_input[35596]), .Z(n9789) );
  AND U14686 ( .A(n9791), .B(n9792), .Z(o[5595]) );
  AND U14687 ( .A(p_input[25595]), .B(p_input[15595]), .Z(n9792) );
  AND U14688 ( .A(p_input[5595]), .B(p_input[35595]), .Z(n9791) );
  AND U14689 ( .A(n9793), .B(n9794), .Z(o[5594]) );
  AND U14690 ( .A(p_input[25594]), .B(p_input[15594]), .Z(n9794) );
  AND U14691 ( .A(p_input[5594]), .B(p_input[35594]), .Z(n9793) );
  AND U14692 ( .A(n9795), .B(n9796), .Z(o[5593]) );
  AND U14693 ( .A(p_input[25593]), .B(p_input[15593]), .Z(n9796) );
  AND U14694 ( .A(p_input[5593]), .B(p_input[35593]), .Z(n9795) );
  AND U14695 ( .A(n9797), .B(n9798), .Z(o[5592]) );
  AND U14696 ( .A(p_input[25592]), .B(p_input[15592]), .Z(n9798) );
  AND U14697 ( .A(p_input[5592]), .B(p_input[35592]), .Z(n9797) );
  AND U14698 ( .A(n9799), .B(n9800), .Z(o[5591]) );
  AND U14699 ( .A(p_input[25591]), .B(p_input[15591]), .Z(n9800) );
  AND U14700 ( .A(p_input[5591]), .B(p_input[35591]), .Z(n9799) );
  AND U14701 ( .A(n9801), .B(n9802), .Z(o[5590]) );
  AND U14702 ( .A(p_input[25590]), .B(p_input[15590]), .Z(n9802) );
  AND U14703 ( .A(p_input[5590]), .B(p_input[35590]), .Z(n9801) );
  AND U14704 ( .A(n9803), .B(n9804), .Z(o[558]) );
  AND U14705 ( .A(p_input[20558]), .B(p_input[10558]), .Z(n9804) );
  AND U14706 ( .A(p_input[558]), .B(p_input[30558]), .Z(n9803) );
  AND U14707 ( .A(n9805), .B(n9806), .Z(o[5589]) );
  AND U14708 ( .A(p_input[25589]), .B(p_input[15589]), .Z(n9806) );
  AND U14709 ( .A(p_input[5589]), .B(p_input[35589]), .Z(n9805) );
  AND U14710 ( .A(n9807), .B(n9808), .Z(o[5588]) );
  AND U14711 ( .A(p_input[25588]), .B(p_input[15588]), .Z(n9808) );
  AND U14712 ( .A(p_input[5588]), .B(p_input[35588]), .Z(n9807) );
  AND U14713 ( .A(n9809), .B(n9810), .Z(o[5587]) );
  AND U14714 ( .A(p_input[25587]), .B(p_input[15587]), .Z(n9810) );
  AND U14715 ( .A(p_input[5587]), .B(p_input[35587]), .Z(n9809) );
  AND U14716 ( .A(n9811), .B(n9812), .Z(o[5586]) );
  AND U14717 ( .A(p_input[25586]), .B(p_input[15586]), .Z(n9812) );
  AND U14718 ( .A(p_input[5586]), .B(p_input[35586]), .Z(n9811) );
  AND U14719 ( .A(n9813), .B(n9814), .Z(o[5585]) );
  AND U14720 ( .A(p_input[25585]), .B(p_input[15585]), .Z(n9814) );
  AND U14721 ( .A(p_input[5585]), .B(p_input[35585]), .Z(n9813) );
  AND U14722 ( .A(n9815), .B(n9816), .Z(o[5584]) );
  AND U14723 ( .A(p_input[25584]), .B(p_input[15584]), .Z(n9816) );
  AND U14724 ( .A(p_input[5584]), .B(p_input[35584]), .Z(n9815) );
  AND U14725 ( .A(n9817), .B(n9818), .Z(o[5583]) );
  AND U14726 ( .A(p_input[25583]), .B(p_input[15583]), .Z(n9818) );
  AND U14727 ( .A(p_input[5583]), .B(p_input[35583]), .Z(n9817) );
  AND U14728 ( .A(n9819), .B(n9820), .Z(o[5582]) );
  AND U14729 ( .A(p_input[25582]), .B(p_input[15582]), .Z(n9820) );
  AND U14730 ( .A(p_input[5582]), .B(p_input[35582]), .Z(n9819) );
  AND U14731 ( .A(n9821), .B(n9822), .Z(o[5581]) );
  AND U14732 ( .A(p_input[25581]), .B(p_input[15581]), .Z(n9822) );
  AND U14733 ( .A(p_input[5581]), .B(p_input[35581]), .Z(n9821) );
  AND U14734 ( .A(n9823), .B(n9824), .Z(o[5580]) );
  AND U14735 ( .A(p_input[25580]), .B(p_input[15580]), .Z(n9824) );
  AND U14736 ( .A(p_input[5580]), .B(p_input[35580]), .Z(n9823) );
  AND U14737 ( .A(n9825), .B(n9826), .Z(o[557]) );
  AND U14738 ( .A(p_input[20557]), .B(p_input[10557]), .Z(n9826) );
  AND U14739 ( .A(p_input[557]), .B(p_input[30557]), .Z(n9825) );
  AND U14740 ( .A(n9827), .B(n9828), .Z(o[5579]) );
  AND U14741 ( .A(p_input[25579]), .B(p_input[15579]), .Z(n9828) );
  AND U14742 ( .A(p_input[5579]), .B(p_input[35579]), .Z(n9827) );
  AND U14743 ( .A(n9829), .B(n9830), .Z(o[5578]) );
  AND U14744 ( .A(p_input[25578]), .B(p_input[15578]), .Z(n9830) );
  AND U14745 ( .A(p_input[5578]), .B(p_input[35578]), .Z(n9829) );
  AND U14746 ( .A(n9831), .B(n9832), .Z(o[5577]) );
  AND U14747 ( .A(p_input[25577]), .B(p_input[15577]), .Z(n9832) );
  AND U14748 ( .A(p_input[5577]), .B(p_input[35577]), .Z(n9831) );
  AND U14749 ( .A(n9833), .B(n9834), .Z(o[5576]) );
  AND U14750 ( .A(p_input[25576]), .B(p_input[15576]), .Z(n9834) );
  AND U14751 ( .A(p_input[5576]), .B(p_input[35576]), .Z(n9833) );
  AND U14752 ( .A(n9835), .B(n9836), .Z(o[5575]) );
  AND U14753 ( .A(p_input[25575]), .B(p_input[15575]), .Z(n9836) );
  AND U14754 ( .A(p_input[5575]), .B(p_input[35575]), .Z(n9835) );
  AND U14755 ( .A(n9837), .B(n9838), .Z(o[5574]) );
  AND U14756 ( .A(p_input[25574]), .B(p_input[15574]), .Z(n9838) );
  AND U14757 ( .A(p_input[5574]), .B(p_input[35574]), .Z(n9837) );
  AND U14758 ( .A(n9839), .B(n9840), .Z(o[5573]) );
  AND U14759 ( .A(p_input[25573]), .B(p_input[15573]), .Z(n9840) );
  AND U14760 ( .A(p_input[5573]), .B(p_input[35573]), .Z(n9839) );
  AND U14761 ( .A(n9841), .B(n9842), .Z(o[5572]) );
  AND U14762 ( .A(p_input[25572]), .B(p_input[15572]), .Z(n9842) );
  AND U14763 ( .A(p_input[5572]), .B(p_input[35572]), .Z(n9841) );
  AND U14764 ( .A(n9843), .B(n9844), .Z(o[5571]) );
  AND U14765 ( .A(p_input[25571]), .B(p_input[15571]), .Z(n9844) );
  AND U14766 ( .A(p_input[5571]), .B(p_input[35571]), .Z(n9843) );
  AND U14767 ( .A(n9845), .B(n9846), .Z(o[5570]) );
  AND U14768 ( .A(p_input[25570]), .B(p_input[15570]), .Z(n9846) );
  AND U14769 ( .A(p_input[5570]), .B(p_input[35570]), .Z(n9845) );
  AND U14770 ( .A(n9847), .B(n9848), .Z(o[556]) );
  AND U14771 ( .A(p_input[20556]), .B(p_input[10556]), .Z(n9848) );
  AND U14772 ( .A(p_input[556]), .B(p_input[30556]), .Z(n9847) );
  AND U14773 ( .A(n9849), .B(n9850), .Z(o[5569]) );
  AND U14774 ( .A(p_input[25569]), .B(p_input[15569]), .Z(n9850) );
  AND U14775 ( .A(p_input[5569]), .B(p_input[35569]), .Z(n9849) );
  AND U14776 ( .A(n9851), .B(n9852), .Z(o[5568]) );
  AND U14777 ( .A(p_input[25568]), .B(p_input[15568]), .Z(n9852) );
  AND U14778 ( .A(p_input[5568]), .B(p_input[35568]), .Z(n9851) );
  AND U14779 ( .A(n9853), .B(n9854), .Z(o[5567]) );
  AND U14780 ( .A(p_input[25567]), .B(p_input[15567]), .Z(n9854) );
  AND U14781 ( .A(p_input[5567]), .B(p_input[35567]), .Z(n9853) );
  AND U14782 ( .A(n9855), .B(n9856), .Z(o[5566]) );
  AND U14783 ( .A(p_input[25566]), .B(p_input[15566]), .Z(n9856) );
  AND U14784 ( .A(p_input[5566]), .B(p_input[35566]), .Z(n9855) );
  AND U14785 ( .A(n9857), .B(n9858), .Z(o[5565]) );
  AND U14786 ( .A(p_input[25565]), .B(p_input[15565]), .Z(n9858) );
  AND U14787 ( .A(p_input[5565]), .B(p_input[35565]), .Z(n9857) );
  AND U14788 ( .A(n9859), .B(n9860), .Z(o[5564]) );
  AND U14789 ( .A(p_input[25564]), .B(p_input[15564]), .Z(n9860) );
  AND U14790 ( .A(p_input[5564]), .B(p_input[35564]), .Z(n9859) );
  AND U14791 ( .A(n9861), .B(n9862), .Z(o[5563]) );
  AND U14792 ( .A(p_input[25563]), .B(p_input[15563]), .Z(n9862) );
  AND U14793 ( .A(p_input[5563]), .B(p_input[35563]), .Z(n9861) );
  AND U14794 ( .A(n9863), .B(n9864), .Z(o[5562]) );
  AND U14795 ( .A(p_input[25562]), .B(p_input[15562]), .Z(n9864) );
  AND U14796 ( .A(p_input[5562]), .B(p_input[35562]), .Z(n9863) );
  AND U14797 ( .A(n9865), .B(n9866), .Z(o[5561]) );
  AND U14798 ( .A(p_input[25561]), .B(p_input[15561]), .Z(n9866) );
  AND U14799 ( .A(p_input[5561]), .B(p_input[35561]), .Z(n9865) );
  AND U14800 ( .A(n9867), .B(n9868), .Z(o[5560]) );
  AND U14801 ( .A(p_input[25560]), .B(p_input[15560]), .Z(n9868) );
  AND U14802 ( .A(p_input[5560]), .B(p_input[35560]), .Z(n9867) );
  AND U14803 ( .A(n9869), .B(n9870), .Z(o[555]) );
  AND U14804 ( .A(p_input[20555]), .B(p_input[10555]), .Z(n9870) );
  AND U14805 ( .A(p_input[555]), .B(p_input[30555]), .Z(n9869) );
  AND U14806 ( .A(n9871), .B(n9872), .Z(o[5559]) );
  AND U14807 ( .A(p_input[25559]), .B(p_input[15559]), .Z(n9872) );
  AND U14808 ( .A(p_input[5559]), .B(p_input[35559]), .Z(n9871) );
  AND U14809 ( .A(n9873), .B(n9874), .Z(o[5558]) );
  AND U14810 ( .A(p_input[25558]), .B(p_input[15558]), .Z(n9874) );
  AND U14811 ( .A(p_input[5558]), .B(p_input[35558]), .Z(n9873) );
  AND U14812 ( .A(n9875), .B(n9876), .Z(o[5557]) );
  AND U14813 ( .A(p_input[25557]), .B(p_input[15557]), .Z(n9876) );
  AND U14814 ( .A(p_input[5557]), .B(p_input[35557]), .Z(n9875) );
  AND U14815 ( .A(n9877), .B(n9878), .Z(o[5556]) );
  AND U14816 ( .A(p_input[25556]), .B(p_input[15556]), .Z(n9878) );
  AND U14817 ( .A(p_input[5556]), .B(p_input[35556]), .Z(n9877) );
  AND U14818 ( .A(n9879), .B(n9880), .Z(o[5555]) );
  AND U14819 ( .A(p_input[25555]), .B(p_input[15555]), .Z(n9880) );
  AND U14820 ( .A(p_input[5555]), .B(p_input[35555]), .Z(n9879) );
  AND U14821 ( .A(n9881), .B(n9882), .Z(o[5554]) );
  AND U14822 ( .A(p_input[25554]), .B(p_input[15554]), .Z(n9882) );
  AND U14823 ( .A(p_input[5554]), .B(p_input[35554]), .Z(n9881) );
  AND U14824 ( .A(n9883), .B(n9884), .Z(o[5553]) );
  AND U14825 ( .A(p_input[25553]), .B(p_input[15553]), .Z(n9884) );
  AND U14826 ( .A(p_input[5553]), .B(p_input[35553]), .Z(n9883) );
  AND U14827 ( .A(n9885), .B(n9886), .Z(o[5552]) );
  AND U14828 ( .A(p_input[25552]), .B(p_input[15552]), .Z(n9886) );
  AND U14829 ( .A(p_input[5552]), .B(p_input[35552]), .Z(n9885) );
  AND U14830 ( .A(n9887), .B(n9888), .Z(o[5551]) );
  AND U14831 ( .A(p_input[25551]), .B(p_input[15551]), .Z(n9888) );
  AND U14832 ( .A(p_input[5551]), .B(p_input[35551]), .Z(n9887) );
  AND U14833 ( .A(n9889), .B(n9890), .Z(o[5550]) );
  AND U14834 ( .A(p_input[25550]), .B(p_input[15550]), .Z(n9890) );
  AND U14835 ( .A(p_input[5550]), .B(p_input[35550]), .Z(n9889) );
  AND U14836 ( .A(n9891), .B(n9892), .Z(o[554]) );
  AND U14837 ( .A(p_input[20554]), .B(p_input[10554]), .Z(n9892) );
  AND U14838 ( .A(p_input[554]), .B(p_input[30554]), .Z(n9891) );
  AND U14839 ( .A(n9893), .B(n9894), .Z(o[5549]) );
  AND U14840 ( .A(p_input[25549]), .B(p_input[15549]), .Z(n9894) );
  AND U14841 ( .A(p_input[5549]), .B(p_input[35549]), .Z(n9893) );
  AND U14842 ( .A(n9895), .B(n9896), .Z(o[5548]) );
  AND U14843 ( .A(p_input[25548]), .B(p_input[15548]), .Z(n9896) );
  AND U14844 ( .A(p_input[5548]), .B(p_input[35548]), .Z(n9895) );
  AND U14845 ( .A(n9897), .B(n9898), .Z(o[5547]) );
  AND U14846 ( .A(p_input[25547]), .B(p_input[15547]), .Z(n9898) );
  AND U14847 ( .A(p_input[5547]), .B(p_input[35547]), .Z(n9897) );
  AND U14848 ( .A(n9899), .B(n9900), .Z(o[5546]) );
  AND U14849 ( .A(p_input[25546]), .B(p_input[15546]), .Z(n9900) );
  AND U14850 ( .A(p_input[5546]), .B(p_input[35546]), .Z(n9899) );
  AND U14851 ( .A(n9901), .B(n9902), .Z(o[5545]) );
  AND U14852 ( .A(p_input[25545]), .B(p_input[15545]), .Z(n9902) );
  AND U14853 ( .A(p_input[5545]), .B(p_input[35545]), .Z(n9901) );
  AND U14854 ( .A(n9903), .B(n9904), .Z(o[5544]) );
  AND U14855 ( .A(p_input[25544]), .B(p_input[15544]), .Z(n9904) );
  AND U14856 ( .A(p_input[5544]), .B(p_input[35544]), .Z(n9903) );
  AND U14857 ( .A(n9905), .B(n9906), .Z(o[5543]) );
  AND U14858 ( .A(p_input[25543]), .B(p_input[15543]), .Z(n9906) );
  AND U14859 ( .A(p_input[5543]), .B(p_input[35543]), .Z(n9905) );
  AND U14860 ( .A(n9907), .B(n9908), .Z(o[5542]) );
  AND U14861 ( .A(p_input[25542]), .B(p_input[15542]), .Z(n9908) );
  AND U14862 ( .A(p_input[5542]), .B(p_input[35542]), .Z(n9907) );
  AND U14863 ( .A(n9909), .B(n9910), .Z(o[5541]) );
  AND U14864 ( .A(p_input[25541]), .B(p_input[15541]), .Z(n9910) );
  AND U14865 ( .A(p_input[5541]), .B(p_input[35541]), .Z(n9909) );
  AND U14866 ( .A(n9911), .B(n9912), .Z(o[5540]) );
  AND U14867 ( .A(p_input[25540]), .B(p_input[15540]), .Z(n9912) );
  AND U14868 ( .A(p_input[5540]), .B(p_input[35540]), .Z(n9911) );
  AND U14869 ( .A(n9913), .B(n9914), .Z(o[553]) );
  AND U14870 ( .A(p_input[20553]), .B(p_input[10553]), .Z(n9914) );
  AND U14871 ( .A(p_input[553]), .B(p_input[30553]), .Z(n9913) );
  AND U14872 ( .A(n9915), .B(n9916), .Z(o[5539]) );
  AND U14873 ( .A(p_input[25539]), .B(p_input[15539]), .Z(n9916) );
  AND U14874 ( .A(p_input[5539]), .B(p_input[35539]), .Z(n9915) );
  AND U14875 ( .A(n9917), .B(n9918), .Z(o[5538]) );
  AND U14876 ( .A(p_input[25538]), .B(p_input[15538]), .Z(n9918) );
  AND U14877 ( .A(p_input[5538]), .B(p_input[35538]), .Z(n9917) );
  AND U14878 ( .A(n9919), .B(n9920), .Z(o[5537]) );
  AND U14879 ( .A(p_input[25537]), .B(p_input[15537]), .Z(n9920) );
  AND U14880 ( .A(p_input[5537]), .B(p_input[35537]), .Z(n9919) );
  AND U14881 ( .A(n9921), .B(n9922), .Z(o[5536]) );
  AND U14882 ( .A(p_input[25536]), .B(p_input[15536]), .Z(n9922) );
  AND U14883 ( .A(p_input[5536]), .B(p_input[35536]), .Z(n9921) );
  AND U14884 ( .A(n9923), .B(n9924), .Z(o[5535]) );
  AND U14885 ( .A(p_input[25535]), .B(p_input[15535]), .Z(n9924) );
  AND U14886 ( .A(p_input[5535]), .B(p_input[35535]), .Z(n9923) );
  AND U14887 ( .A(n9925), .B(n9926), .Z(o[5534]) );
  AND U14888 ( .A(p_input[25534]), .B(p_input[15534]), .Z(n9926) );
  AND U14889 ( .A(p_input[5534]), .B(p_input[35534]), .Z(n9925) );
  AND U14890 ( .A(n9927), .B(n9928), .Z(o[5533]) );
  AND U14891 ( .A(p_input[25533]), .B(p_input[15533]), .Z(n9928) );
  AND U14892 ( .A(p_input[5533]), .B(p_input[35533]), .Z(n9927) );
  AND U14893 ( .A(n9929), .B(n9930), .Z(o[5532]) );
  AND U14894 ( .A(p_input[25532]), .B(p_input[15532]), .Z(n9930) );
  AND U14895 ( .A(p_input[5532]), .B(p_input[35532]), .Z(n9929) );
  AND U14896 ( .A(n9931), .B(n9932), .Z(o[5531]) );
  AND U14897 ( .A(p_input[25531]), .B(p_input[15531]), .Z(n9932) );
  AND U14898 ( .A(p_input[5531]), .B(p_input[35531]), .Z(n9931) );
  AND U14899 ( .A(n9933), .B(n9934), .Z(o[5530]) );
  AND U14900 ( .A(p_input[25530]), .B(p_input[15530]), .Z(n9934) );
  AND U14901 ( .A(p_input[5530]), .B(p_input[35530]), .Z(n9933) );
  AND U14902 ( .A(n9935), .B(n9936), .Z(o[552]) );
  AND U14903 ( .A(p_input[20552]), .B(p_input[10552]), .Z(n9936) );
  AND U14904 ( .A(p_input[552]), .B(p_input[30552]), .Z(n9935) );
  AND U14905 ( .A(n9937), .B(n9938), .Z(o[5529]) );
  AND U14906 ( .A(p_input[25529]), .B(p_input[15529]), .Z(n9938) );
  AND U14907 ( .A(p_input[5529]), .B(p_input[35529]), .Z(n9937) );
  AND U14908 ( .A(n9939), .B(n9940), .Z(o[5528]) );
  AND U14909 ( .A(p_input[25528]), .B(p_input[15528]), .Z(n9940) );
  AND U14910 ( .A(p_input[5528]), .B(p_input[35528]), .Z(n9939) );
  AND U14911 ( .A(n9941), .B(n9942), .Z(o[5527]) );
  AND U14912 ( .A(p_input[25527]), .B(p_input[15527]), .Z(n9942) );
  AND U14913 ( .A(p_input[5527]), .B(p_input[35527]), .Z(n9941) );
  AND U14914 ( .A(n9943), .B(n9944), .Z(o[5526]) );
  AND U14915 ( .A(p_input[25526]), .B(p_input[15526]), .Z(n9944) );
  AND U14916 ( .A(p_input[5526]), .B(p_input[35526]), .Z(n9943) );
  AND U14917 ( .A(n9945), .B(n9946), .Z(o[5525]) );
  AND U14918 ( .A(p_input[25525]), .B(p_input[15525]), .Z(n9946) );
  AND U14919 ( .A(p_input[5525]), .B(p_input[35525]), .Z(n9945) );
  AND U14920 ( .A(n9947), .B(n9948), .Z(o[5524]) );
  AND U14921 ( .A(p_input[25524]), .B(p_input[15524]), .Z(n9948) );
  AND U14922 ( .A(p_input[5524]), .B(p_input[35524]), .Z(n9947) );
  AND U14923 ( .A(n9949), .B(n9950), .Z(o[5523]) );
  AND U14924 ( .A(p_input[25523]), .B(p_input[15523]), .Z(n9950) );
  AND U14925 ( .A(p_input[5523]), .B(p_input[35523]), .Z(n9949) );
  AND U14926 ( .A(n9951), .B(n9952), .Z(o[5522]) );
  AND U14927 ( .A(p_input[25522]), .B(p_input[15522]), .Z(n9952) );
  AND U14928 ( .A(p_input[5522]), .B(p_input[35522]), .Z(n9951) );
  AND U14929 ( .A(n9953), .B(n9954), .Z(o[5521]) );
  AND U14930 ( .A(p_input[25521]), .B(p_input[15521]), .Z(n9954) );
  AND U14931 ( .A(p_input[5521]), .B(p_input[35521]), .Z(n9953) );
  AND U14932 ( .A(n9955), .B(n9956), .Z(o[5520]) );
  AND U14933 ( .A(p_input[25520]), .B(p_input[15520]), .Z(n9956) );
  AND U14934 ( .A(p_input[5520]), .B(p_input[35520]), .Z(n9955) );
  AND U14935 ( .A(n9957), .B(n9958), .Z(o[551]) );
  AND U14936 ( .A(p_input[20551]), .B(p_input[10551]), .Z(n9958) );
  AND U14937 ( .A(p_input[551]), .B(p_input[30551]), .Z(n9957) );
  AND U14938 ( .A(n9959), .B(n9960), .Z(o[5519]) );
  AND U14939 ( .A(p_input[25519]), .B(p_input[15519]), .Z(n9960) );
  AND U14940 ( .A(p_input[5519]), .B(p_input[35519]), .Z(n9959) );
  AND U14941 ( .A(n9961), .B(n9962), .Z(o[5518]) );
  AND U14942 ( .A(p_input[25518]), .B(p_input[15518]), .Z(n9962) );
  AND U14943 ( .A(p_input[5518]), .B(p_input[35518]), .Z(n9961) );
  AND U14944 ( .A(n9963), .B(n9964), .Z(o[5517]) );
  AND U14945 ( .A(p_input[25517]), .B(p_input[15517]), .Z(n9964) );
  AND U14946 ( .A(p_input[5517]), .B(p_input[35517]), .Z(n9963) );
  AND U14947 ( .A(n9965), .B(n9966), .Z(o[5516]) );
  AND U14948 ( .A(p_input[25516]), .B(p_input[15516]), .Z(n9966) );
  AND U14949 ( .A(p_input[5516]), .B(p_input[35516]), .Z(n9965) );
  AND U14950 ( .A(n9967), .B(n9968), .Z(o[5515]) );
  AND U14951 ( .A(p_input[25515]), .B(p_input[15515]), .Z(n9968) );
  AND U14952 ( .A(p_input[5515]), .B(p_input[35515]), .Z(n9967) );
  AND U14953 ( .A(n9969), .B(n9970), .Z(o[5514]) );
  AND U14954 ( .A(p_input[25514]), .B(p_input[15514]), .Z(n9970) );
  AND U14955 ( .A(p_input[5514]), .B(p_input[35514]), .Z(n9969) );
  AND U14956 ( .A(n9971), .B(n9972), .Z(o[5513]) );
  AND U14957 ( .A(p_input[25513]), .B(p_input[15513]), .Z(n9972) );
  AND U14958 ( .A(p_input[5513]), .B(p_input[35513]), .Z(n9971) );
  AND U14959 ( .A(n9973), .B(n9974), .Z(o[5512]) );
  AND U14960 ( .A(p_input[25512]), .B(p_input[15512]), .Z(n9974) );
  AND U14961 ( .A(p_input[5512]), .B(p_input[35512]), .Z(n9973) );
  AND U14962 ( .A(n9975), .B(n9976), .Z(o[5511]) );
  AND U14963 ( .A(p_input[25511]), .B(p_input[15511]), .Z(n9976) );
  AND U14964 ( .A(p_input[5511]), .B(p_input[35511]), .Z(n9975) );
  AND U14965 ( .A(n9977), .B(n9978), .Z(o[5510]) );
  AND U14966 ( .A(p_input[25510]), .B(p_input[15510]), .Z(n9978) );
  AND U14967 ( .A(p_input[5510]), .B(p_input[35510]), .Z(n9977) );
  AND U14968 ( .A(n9979), .B(n9980), .Z(o[550]) );
  AND U14969 ( .A(p_input[20550]), .B(p_input[10550]), .Z(n9980) );
  AND U14970 ( .A(p_input[550]), .B(p_input[30550]), .Z(n9979) );
  AND U14971 ( .A(n9981), .B(n9982), .Z(o[5509]) );
  AND U14972 ( .A(p_input[25509]), .B(p_input[15509]), .Z(n9982) );
  AND U14973 ( .A(p_input[5509]), .B(p_input[35509]), .Z(n9981) );
  AND U14974 ( .A(n9983), .B(n9984), .Z(o[5508]) );
  AND U14975 ( .A(p_input[25508]), .B(p_input[15508]), .Z(n9984) );
  AND U14976 ( .A(p_input[5508]), .B(p_input[35508]), .Z(n9983) );
  AND U14977 ( .A(n9985), .B(n9986), .Z(o[5507]) );
  AND U14978 ( .A(p_input[25507]), .B(p_input[15507]), .Z(n9986) );
  AND U14979 ( .A(p_input[5507]), .B(p_input[35507]), .Z(n9985) );
  AND U14980 ( .A(n9987), .B(n9988), .Z(o[5506]) );
  AND U14981 ( .A(p_input[25506]), .B(p_input[15506]), .Z(n9988) );
  AND U14982 ( .A(p_input[5506]), .B(p_input[35506]), .Z(n9987) );
  AND U14983 ( .A(n9989), .B(n9990), .Z(o[5505]) );
  AND U14984 ( .A(p_input[25505]), .B(p_input[15505]), .Z(n9990) );
  AND U14985 ( .A(p_input[5505]), .B(p_input[35505]), .Z(n9989) );
  AND U14986 ( .A(n9991), .B(n9992), .Z(o[5504]) );
  AND U14987 ( .A(p_input[25504]), .B(p_input[15504]), .Z(n9992) );
  AND U14988 ( .A(p_input[5504]), .B(p_input[35504]), .Z(n9991) );
  AND U14989 ( .A(n9993), .B(n9994), .Z(o[5503]) );
  AND U14990 ( .A(p_input[25503]), .B(p_input[15503]), .Z(n9994) );
  AND U14991 ( .A(p_input[5503]), .B(p_input[35503]), .Z(n9993) );
  AND U14992 ( .A(n9995), .B(n9996), .Z(o[5502]) );
  AND U14993 ( .A(p_input[25502]), .B(p_input[15502]), .Z(n9996) );
  AND U14994 ( .A(p_input[5502]), .B(p_input[35502]), .Z(n9995) );
  AND U14995 ( .A(n9997), .B(n9998), .Z(o[5501]) );
  AND U14996 ( .A(p_input[25501]), .B(p_input[15501]), .Z(n9998) );
  AND U14997 ( .A(p_input[5501]), .B(p_input[35501]), .Z(n9997) );
  AND U14998 ( .A(n9999), .B(n10000), .Z(o[5500]) );
  AND U14999 ( .A(p_input[25500]), .B(p_input[15500]), .Z(n10000) );
  AND U15000 ( .A(p_input[5500]), .B(p_input[35500]), .Z(n9999) );
  AND U15001 ( .A(n10001), .B(n10002), .Z(o[54]) );
  AND U15002 ( .A(p_input[20054]), .B(p_input[10054]), .Z(n10002) );
  AND U15003 ( .A(p_input[54]), .B(p_input[30054]), .Z(n10001) );
  AND U15004 ( .A(n10003), .B(n10004), .Z(o[549]) );
  AND U15005 ( .A(p_input[20549]), .B(p_input[10549]), .Z(n10004) );
  AND U15006 ( .A(p_input[549]), .B(p_input[30549]), .Z(n10003) );
  AND U15007 ( .A(n10005), .B(n10006), .Z(o[5499]) );
  AND U15008 ( .A(p_input[25499]), .B(p_input[15499]), .Z(n10006) );
  AND U15009 ( .A(p_input[5499]), .B(p_input[35499]), .Z(n10005) );
  AND U15010 ( .A(n10007), .B(n10008), .Z(o[5498]) );
  AND U15011 ( .A(p_input[25498]), .B(p_input[15498]), .Z(n10008) );
  AND U15012 ( .A(p_input[5498]), .B(p_input[35498]), .Z(n10007) );
  AND U15013 ( .A(n10009), .B(n10010), .Z(o[5497]) );
  AND U15014 ( .A(p_input[25497]), .B(p_input[15497]), .Z(n10010) );
  AND U15015 ( .A(p_input[5497]), .B(p_input[35497]), .Z(n10009) );
  AND U15016 ( .A(n10011), .B(n10012), .Z(o[5496]) );
  AND U15017 ( .A(p_input[25496]), .B(p_input[15496]), .Z(n10012) );
  AND U15018 ( .A(p_input[5496]), .B(p_input[35496]), .Z(n10011) );
  AND U15019 ( .A(n10013), .B(n10014), .Z(o[5495]) );
  AND U15020 ( .A(p_input[25495]), .B(p_input[15495]), .Z(n10014) );
  AND U15021 ( .A(p_input[5495]), .B(p_input[35495]), .Z(n10013) );
  AND U15022 ( .A(n10015), .B(n10016), .Z(o[5494]) );
  AND U15023 ( .A(p_input[25494]), .B(p_input[15494]), .Z(n10016) );
  AND U15024 ( .A(p_input[5494]), .B(p_input[35494]), .Z(n10015) );
  AND U15025 ( .A(n10017), .B(n10018), .Z(o[5493]) );
  AND U15026 ( .A(p_input[25493]), .B(p_input[15493]), .Z(n10018) );
  AND U15027 ( .A(p_input[5493]), .B(p_input[35493]), .Z(n10017) );
  AND U15028 ( .A(n10019), .B(n10020), .Z(o[5492]) );
  AND U15029 ( .A(p_input[25492]), .B(p_input[15492]), .Z(n10020) );
  AND U15030 ( .A(p_input[5492]), .B(p_input[35492]), .Z(n10019) );
  AND U15031 ( .A(n10021), .B(n10022), .Z(o[5491]) );
  AND U15032 ( .A(p_input[25491]), .B(p_input[15491]), .Z(n10022) );
  AND U15033 ( .A(p_input[5491]), .B(p_input[35491]), .Z(n10021) );
  AND U15034 ( .A(n10023), .B(n10024), .Z(o[5490]) );
  AND U15035 ( .A(p_input[25490]), .B(p_input[15490]), .Z(n10024) );
  AND U15036 ( .A(p_input[5490]), .B(p_input[35490]), .Z(n10023) );
  AND U15037 ( .A(n10025), .B(n10026), .Z(o[548]) );
  AND U15038 ( .A(p_input[20548]), .B(p_input[10548]), .Z(n10026) );
  AND U15039 ( .A(p_input[548]), .B(p_input[30548]), .Z(n10025) );
  AND U15040 ( .A(n10027), .B(n10028), .Z(o[5489]) );
  AND U15041 ( .A(p_input[25489]), .B(p_input[15489]), .Z(n10028) );
  AND U15042 ( .A(p_input[5489]), .B(p_input[35489]), .Z(n10027) );
  AND U15043 ( .A(n10029), .B(n10030), .Z(o[5488]) );
  AND U15044 ( .A(p_input[25488]), .B(p_input[15488]), .Z(n10030) );
  AND U15045 ( .A(p_input[5488]), .B(p_input[35488]), .Z(n10029) );
  AND U15046 ( .A(n10031), .B(n10032), .Z(o[5487]) );
  AND U15047 ( .A(p_input[25487]), .B(p_input[15487]), .Z(n10032) );
  AND U15048 ( .A(p_input[5487]), .B(p_input[35487]), .Z(n10031) );
  AND U15049 ( .A(n10033), .B(n10034), .Z(o[5486]) );
  AND U15050 ( .A(p_input[25486]), .B(p_input[15486]), .Z(n10034) );
  AND U15051 ( .A(p_input[5486]), .B(p_input[35486]), .Z(n10033) );
  AND U15052 ( .A(n10035), .B(n10036), .Z(o[5485]) );
  AND U15053 ( .A(p_input[25485]), .B(p_input[15485]), .Z(n10036) );
  AND U15054 ( .A(p_input[5485]), .B(p_input[35485]), .Z(n10035) );
  AND U15055 ( .A(n10037), .B(n10038), .Z(o[5484]) );
  AND U15056 ( .A(p_input[25484]), .B(p_input[15484]), .Z(n10038) );
  AND U15057 ( .A(p_input[5484]), .B(p_input[35484]), .Z(n10037) );
  AND U15058 ( .A(n10039), .B(n10040), .Z(o[5483]) );
  AND U15059 ( .A(p_input[25483]), .B(p_input[15483]), .Z(n10040) );
  AND U15060 ( .A(p_input[5483]), .B(p_input[35483]), .Z(n10039) );
  AND U15061 ( .A(n10041), .B(n10042), .Z(o[5482]) );
  AND U15062 ( .A(p_input[25482]), .B(p_input[15482]), .Z(n10042) );
  AND U15063 ( .A(p_input[5482]), .B(p_input[35482]), .Z(n10041) );
  AND U15064 ( .A(n10043), .B(n10044), .Z(o[5481]) );
  AND U15065 ( .A(p_input[25481]), .B(p_input[15481]), .Z(n10044) );
  AND U15066 ( .A(p_input[5481]), .B(p_input[35481]), .Z(n10043) );
  AND U15067 ( .A(n10045), .B(n10046), .Z(o[5480]) );
  AND U15068 ( .A(p_input[25480]), .B(p_input[15480]), .Z(n10046) );
  AND U15069 ( .A(p_input[5480]), .B(p_input[35480]), .Z(n10045) );
  AND U15070 ( .A(n10047), .B(n10048), .Z(o[547]) );
  AND U15071 ( .A(p_input[20547]), .B(p_input[10547]), .Z(n10048) );
  AND U15072 ( .A(p_input[547]), .B(p_input[30547]), .Z(n10047) );
  AND U15073 ( .A(n10049), .B(n10050), .Z(o[5479]) );
  AND U15074 ( .A(p_input[25479]), .B(p_input[15479]), .Z(n10050) );
  AND U15075 ( .A(p_input[5479]), .B(p_input[35479]), .Z(n10049) );
  AND U15076 ( .A(n10051), .B(n10052), .Z(o[5478]) );
  AND U15077 ( .A(p_input[25478]), .B(p_input[15478]), .Z(n10052) );
  AND U15078 ( .A(p_input[5478]), .B(p_input[35478]), .Z(n10051) );
  AND U15079 ( .A(n10053), .B(n10054), .Z(o[5477]) );
  AND U15080 ( .A(p_input[25477]), .B(p_input[15477]), .Z(n10054) );
  AND U15081 ( .A(p_input[5477]), .B(p_input[35477]), .Z(n10053) );
  AND U15082 ( .A(n10055), .B(n10056), .Z(o[5476]) );
  AND U15083 ( .A(p_input[25476]), .B(p_input[15476]), .Z(n10056) );
  AND U15084 ( .A(p_input[5476]), .B(p_input[35476]), .Z(n10055) );
  AND U15085 ( .A(n10057), .B(n10058), .Z(o[5475]) );
  AND U15086 ( .A(p_input[25475]), .B(p_input[15475]), .Z(n10058) );
  AND U15087 ( .A(p_input[5475]), .B(p_input[35475]), .Z(n10057) );
  AND U15088 ( .A(n10059), .B(n10060), .Z(o[5474]) );
  AND U15089 ( .A(p_input[25474]), .B(p_input[15474]), .Z(n10060) );
  AND U15090 ( .A(p_input[5474]), .B(p_input[35474]), .Z(n10059) );
  AND U15091 ( .A(n10061), .B(n10062), .Z(o[5473]) );
  AND U15092 ( .A(p_input[25473]), .B(p_input[15473]), .Z(n10062) );
  AND U15093 ( .A(p_input[5473]), .B(p_input[35473]), .Z(n10061) );
  AND U15094 ( .A(n10063), .B(n10064), .Z(o[5472]) );
  AND U15095 ( .A(p_input[25472]), .B(p_input[15472]), .Z(n10064) );
  AND U15096 ( .A(p_input[5472]), .B(p_input[35472]), .Z(n10063) );
  AND U15097 ( .A(n10065), .B(n10066), .Z(o[5471]) );
  AND U15098 ( .A(p_input[25471]), .B(p_input[15471]), .Z(n10066) );
  AND U15099 ( .A(p_input[5471]), .B(p_input[35471]), .Z(n10065) );
  AND U15100 ( .A(n10067), .B(n10068), .Z(o[5470]) );
  AND U15101 ( .A(p_input[25470]), .B(p_input[15470]), .Z(n10068) );
  AND U15102 ( .A(p_input[5470]), .B(p_input[35470]), .Z(n10067) );
  AND U15103 ( .A(n10069), .B(n10070), .Z(o[546]) );
  AND U15104 ( .A(p_input[20546]), .B(p_input[10546]), .Z(n10070) );
  AND U15105 ( .A(p_input[546]), .B(p_input[30546]), .Z(n10069) );
  AND U15106 ( .A(n10071), .B(n10072), .Z(o[5469]) );
  AND U15107 ( .A(p_input[25469]), .B(p_input[15469]), .Z(n10072) );
  AND U15108 ( .A(p_input[5469]), .B(p_input[35469]), .Z(n10071) );
  AND U15109 ( .A(n10073), .B(n10074), .Z(o[5468]) );
  AND U15110 ( .A(p_input[25468]), .B(p_input[15468]), .Z(n10074) );
  AND U15111 ( .A(p_input[5468]), .B(p_input[35468]), .Z(n10073) );
  AND U15112 ( .A(n10075), .B(n10076), .Z(o[5467]) );
  AND U15113 ( .A(p_input[25467]), .B(p_input[15467]), .Z(n10076) );
  AND U15114 ( .A(p_input[5467]), .B(p_input[35467]), .Z(n10075) );
  AND U15115 ( .A(n10077), .B(n10078), .Z(o[5466]) );
  AND U15116 ( .A(p_input[25466]), .B(p_input[15466]), .Z(n10078) );
  AND U15117 ( .A(p_input[5466]), .B(p_input[35466]), .Z(n10077) );
  AND U15118 ( .A(n10079), .B(n10080), .Z(o[5465]) );
  AND U15119 ( .A(p_input[25465]), .B(p_input[15465]), .Z(n10080) );
  AND U15120 ( .A(p_input[5465]), .B(p_input[35465]), .Z(n10079) );
  AND U15121 ( .A(n10081), .B(n10082), .Z(o[5464]) );
  AND U15122 ( .A(p_input[25464]), .B(p_input[15464]), .Z(n10082) );
  AND U15123 ( .A(p_input[5464]), .B(p_input[35464]), .Z(n10081) );
  AND U15124 ( .A(n10083), .B(n10084), .Z(o[5463]) );
  AND U15125 ( .A(p_input[25463]), .B(p_input[15463]), .Z(n10084) );
  AND U15126 ( .A(p_input[5463]), .B(p_input[35463]), .Z(n10083) );
  AND U15127 ( .A(n10085), .B(n10086), .Z(o[5462]) );
  AND U15128 ( .A(p_input[25462]), .B(p_input[15462]), .Z(n10086) );
  AND U15129 ( .A(p_input[5462]), .B(p_input[35462]), .Z(n10085) );
  AND U15130 ( .A(n10087), .B(n10088), .Z(o[5461]) );
  AND U15131 ( .A(p_input[25461]), .B(p_input[15461]), .Z(n10088) );
  AND U15132 ( .A(p_input[5461]), .B(p_input[35461]), .Z(n10087) );
  AND U15133 ( .A(n10089), .B(n10090), .Z(o[5460]) );
  AND U15134 ( .A(p_input[25460]), .B(p_input[15460]), .Z(n10090) );
  AND U15135 ( .A(p_input[5460]), .B(p_input[35460]), .Z(n10089) );
  AND U15136 ( .A(n10091), .B(n10092), .Z(o[545]) );
  AND U15137 ( .A(p_input[20545]), .B(p_input[10545]), .Z(n10092) );
  AND U15138 ( .A(p_input[545]), .B(p_input[30545]), .Z(n10091) );
  AND U15139 ( .A(n10093), .B(n10094), .Z(o[5459]) );
  AND U15140 ( .A(p_input[25459]), .B(p_input[15459]), .Z(n10094) );
  AND U15141 ( .A(p_input[5459]), .B(p_input[35459]), .Z(n10093) );
  AND U15142 ( .A(n10095), .B(n10096), .Z(o[5458]) );
  AND U15143 ( .A(p_input[25458]), .B(p_input[15458]), .Z(n10096) );
  AND U15144 ( .A(p_input[5458]), .B(p_input[35458]), .Z(n10095) );
  AND U15145 ( .A(n10097), .B(n10098), .Z(o[5457]) );
  AND U15146 ( .A(p_input[25457]), .B(p_input[15457]), .Z(n10098) );
  AND U15147 ( .A(p_input[5457]), .B(p_input[35457]), .Z(n10097) );
  AND U15148 ( .A(n10099), .B(n10100), .Z(o[5456]) );
  AND U15149 ( .A(p_input[25456]), .B(p_input[15456]), .Z(n10100) );
  AND U15150 ( .A(p_input[5456]), .B(p_input[35456]), .Z(n10099) );
  AND U15151 ( .A(n10101), .B(n10102), .Z(o[5455]) );
  AND U15152 ( .A(p_input[25455]), .B(p_input[15455]), .Z(n10102) );
  AND U15153 ( .A(p_input[5455]), .B(p_input[35455]), .Z(n10101) );
  AND U15154 ( .A(n10103), .B(n10104), .Z(o[5454]) );
  AND U15155 ( .A(p_input[25454]), .B(p_input[15454]), .Z(n10104) );
  AND U15156 ( .A(p_input[5454]), .B(p_input[35454]), .Z(n10103) );
  AND U15157 ( .A(n10105), .B(n10106), .Z(o[5453]) );
  AND U15158 ( .A(p_input[25453]), .B(p_input[15453]), .Z(n10106) );
  AND U15159 ( .A(p_input[5453]), .B(p_input[35453]), .Z(n10105) );
  AND U15160 ( .A(n10107), .B(n10108), .Z(o[5452]) );
  AND U15161 ( .A(p_input[25452]), .B(p_input[15452]), .Z(n10108) );
  AND U15162 ( .A(p_input[5452]), .B(p_input[35452]), .Z(n10107) );
  AND U15163 ( .A(n10109), .B(n10110), .Z(o[5451]) );
  AND U15164 ( .A(p_input[25451]), .B(p_input[15451]), .Z(n10110) );
  AND U15165 ( .A(p_input[5451]), .B(p_input[35451]), .Z(n10109) );
  AND U15166 ( .A(n10111), .B(n10112), .Z(o[5450]) );
  AND U15167 ( .A(p_input[25450]), .B(p_input[15450]), .Z(n10112) );
  AND U15168 ( .A(p_input[5450]), .B(p_input[35450]), .Z(n10111) );
  AND U15169 ( .A(n10113), .B(n10114), .Z(o[544]) );
  AND U15170 ( .A(p_input[20544]), .B(p_input[10544]), .Z(n10114) );
  AND U15171 ( .A(p_input[544]), .B(p_input[30544]), .Z(n10113) );
  AND U15172 ( .A(n10115), .B(n10116), .Z(o[5449]) );
  AND U15173 ( .A(p_input[25449]), .B(p_input[15449]), .Z(n10116) );
  AND U15174 ( .A(p_input[5449]), .B(p_input[35449]), .Z(n10115) );
  AND U15175 ( .A(n10117), .B(n10118), .Z(o[5448]) );
  AND U15176 ( .A(p_input[25448]), .B(p_input[15448]), .Z(n10118) );
  AND U15177 ( .A(p_input[5448]), .B(p_input[35448]), .Z(n10117) );
  AND U15178 ( .A(n10119), .B(n10120), .Z(o[5447]) );
  AND U15179 ( .A(p_input[25447]), .B(p_input[15447]), .Z(n10120) );
  AND U15180 ( .A(p_input[5447]), .B(p_input[35447]), .Z(n10119) );
  AND U15181 ( .A(n10121), .B(n10122), .Z(o[5446]) );
  AND U15182 ( .A(p_input[25446]), .B(p_input[15446]), .Z(n10122) );
  AND U15183 ( .A(p_input[5446]), .B(p_input[35446]), .Z(n10121) );
  AND U15184 ( .A(n10123), .B(n10124), .Z(o[5445]) );
  AND U15185 ( .A(p_input[25445]), .B(p_input[15445]), .Z(n10124) );
  AND U15186 ( .A(p_input[5445]), .B(p_input[35445]), .Z(n10123) );
  AND U15187 ( .A(n10125), .B(n10126), .Z(o[5444]) );
  AND U15188 ( .A(p_input[25444]), .B(p_input[15444]), .Z(n10126) );
  AND U15189 ( .A(p_input[5444]), .B(p_input[35444]), .Z(n10125) );
  AND U15190 ( .A(n10127), .B(n10128), .Z(o[5443]) );
  AND U15191 ( .A(p_input[25443]), .B(p_input[15443]), .Z(n10128) );
  AND U15192 ( .A(p_input[5443]), .B(p_input[35443]), .Z(n10127) );
  AND U15193 ( .A(n10129), .B(n10130), .Z(o[5442]) );
  AND U15194 ( .A(p_input[25442]), .B(p_input[15442]), .Z(n10130) );
  AND U15195 ( .A(p_input[5442]), .B(p_input[35442]), .Z(n10129) );
  AND U15196 ( .A(n10131), .B(n10132), .Z(o[5441]) );
  AND U15197 ( .A(p_input[25441]), .B(p_input[15441]), .Z(n10132) );
  AND U15198 ( .A(p_input[5441]), .B(p_input[35441]), .Z(n10131) );
  AND U15199 ( .A(n10133), .B(n10134), .Z(o[5440]) );
  AND U15200 ( .A(p_input[25440]), .B(p_input[15440]), .Z(n10134) );
  AND U15201 ( .A(p_input[5440]), .B(p_input[35440]), .Z(n10133) );
  AND U15202 ( .A(n10135), .B(n10136), .Z(o[543]) );
  AND U15203 ( .A(p_input[20543]), .B(p_input[10543]), .Z(n10136) );
  AND U15204 ( .A(p_input[543]), .B(p_input[30543]), .Z(n10135) );
  AND U15205 ( .A(n10137), .B(n10138), .Z(o[5439]) );
  AND U15206 ( .A(p_input[25439]), .B(p_input[15439]), .Z(n10138) );
  AND U15207 ( .A(p_input[5439]), .B(p_input[35439]), .Z(n10137) );
  AND U15208 ( .A(n10139), .B(n10140), .Z(o[5438]) );
  AND U15209 ( .A(p_input[25438]), .B(p_input[15438]), .Z(n10140) );
  AND U15210 ( .A(p_input[5438]), .B(p_input[35438]), .Z(n10139) );
  AND U15211 ( .A(n10141), .B(n10142), .Z(o[5437]) );
  AND U15212 ( .A(p_input[25437]), .B(p_input[15437]), .Z(n10142) );
  AND U15213 ( .A(p_input[5437]), .B(p_input[35437]), .Z(n10141) );
  AND U15214 ( .A(n10143), .B(n10144), .Z(o[5436]) );
  AND U15215 ( .A(p_input[25436]), .B(p_input[15436]), .Z(n10144) );
  AND U15216 ( .A(p_input[5436]), .B(p_input[35436]), .Z(n10143) );
  AND U15217 ( .A(n10145), .B(n10146), .Z(o[5435]) );
  AND U15218 ( .A(p_input[25435]), .B(p_input[15435]), .Z(n10146) );
  AND U15219 ( .A(p_input[5435]), .B(p_input[35435]), .Z(n10145) );
  AND U15220 ( .A(n10147), .B(n10148), .Z(o[5434]) );
  AND U15221 ( .A(p_input[25434]), .B(p_input[15434]), .Z(n10148) );
  AND U15222 ( .A(p_input[5434]), .B(p_input[35434]), .Z(n10147) );
  AND U15223 ( .A(n10149), .B(n10150), .Z(o[5433]) );
  AND U15224 ( .A(p_input[25433]), .B(p_input[15433]), .Z(n10150) );
  AND U15225 ( .A(p_input[5433]), .B(p_input[35433]), .Z(n10149) );
  AND U15226 ( .A(n10151), .B(n10152), .Z(o[5432]) );
  AND U15227 ( .A(p_input[25432]), .B(p_input[15432]), .Z(n10152) );
  AND U15228 ( .A(p_input[5432]), .B(p_input[35432]), .Z(n10151) );
  AND U15229 ( .A(n10153), .B(n10154), .Z(o[5431]) );
  AND U15230 ( .A(p_input[25431]), .B(p_input[15431]), .Z(n10154) );
  AND U15231 ( .A(p_input[5431]), .B(p_input[35431]), .Z(n10153) );
  AND U15232 ( .A(n10155), .B(n10156), .Z(o[5430]) );
  AND U15233 ( .A(p_input[25430]), .B(p_input[15430]), .Z(n10156) );
  AND U15234 ( .A(p_input[5430]), .B(p_input[35430]), .Z(n10155) );
  AND U15235 ( .A(n10157), .B(n10158), .Z(o[542]) );
  AND U15236 ( .A(p_input[20542]), .B(p_input[10542]), .Z(n10158) );
  AND U15237 ( .A(p_input[542]), .B(p_input[30542]), .Z(n10157) );
  AND U15238 ( .A(n10159), .B(n10160), .Z(o[5429]) );
  AND U15239 ( .A(p_input[25429]), .B(p_input[15429]), .Z(n10160) );
  AND U15240 ( .A(p_input[5429]), .B(p_input[35429]), .Z(n10159) );
  AND U15241 ( .A(n10161), .B(n10162), .Z(o[5428]) );
  AND U15242 ( .A(p_input[25428]), .B(p_input[15428]), .Z(n10162) );
  AND U15243 ( .A(p_input[5428]), .B(p_input[35428]), .Z(n10161) );
  AND U15244 ( .A(n10163), .B(n10164), .Z(o[5427]) );
  AND U15245 ( .A(p_input[25427]), .B(p_input[15427]), .Z(n10164) );
  AND U15246 ( .A(p_input[5427]), .B(p_input[35427]), .Z(n10163) );
  AND U15247 ( .A(n10165), .B(n10166), .Z(o[5426]) );
  AND U15248 ( .A(p_input[25426]), .B(p_input[15426]), .Z(n10166) );
  AND U15249 ( .A(p_input[5426]), .B(p_input[35426]), .Z(n10165) );
  AND U15250 ( .A(n10167), .B(n10168), .Z(o[5425]) );
  AND U15251 ( .A(p_input[25425]), .B(p_input[15425]), .Z(n10168) );
  AND U15252 ( .A(p_input[5425]), .B(p_input[35425]), .Z(n10167) );
  AND U15253 ( .A(n10169), .B(n10170), .Z(o[5424]) );
  AND U15254 ( .A(p_input[25424]), .B(p_input[15424]), .Z(n10170) );
  AND U15255 ( .A(p_input[5424]), .B(p_input[35424]), .Z(n10169) );
  AND U15256 ( .A(n10171), .B(n10172), .Z(o[5423]) );
  AND U15257 ( .A(p_input[25423]), .B(p_input[15423]), .Z(n10172) );
  AND U15258 ( .A(p_input[5423]), .B(p_input[35423]), .Z(n10171) );
  AND U15259 ( .A(n10173), .B(n10174), .Z(o[5422]) );
  AND U15260 ( .A(p_input[25422]), .B(p_input[15422]), .Z(n10174) );
  AND U15261 ( .A(p_input[5422]), .B(p_input[35422]), .Z(n10173) );
  AND U15262 ( .A(n10175), .B(n10176), .Z(o[5421]) );
  AND U15263 ( .A(p_input[25421]), .B(p_input[15421]), .Z(n10176) );
  AND U15264 ( .A(p_input[5421]), .B(p_input[35421]), .Z(n10175) );
  AND U15265 ( .A(n10177), .B(n10178), .Z(o[5420]) );
  AND U15266 ( .A(p_input[25420]), .B(p_input[15420]), .Z(n10178) );
  AND U15267 ( .A(p_input[5420]), .B(p_input[35420]), .Z(n10177) );
  AND U15268 ( .A(n10179), .B(n10180), .Z(o[541]) );
  AND U15269 ( .A(p_input[20541]), .B(p_input[10541]), .Z(n10180) );
  AND U15270 ( .A(p_input[541]), .B(p_input[30541]), .Z(n10179) );
  AND U15271 ( .A(n10181), .B(n10182), .Z(o[5419]) );
  AND U15272 ( .A(p_input[25419]), .B(p_input[15419]), .Z(n10182) );
  AND U15273 ( .A(p_input[5419]), .B(p_input[35419]), .Z(n10181) );
  AND U15274 ( .A(n10183), .B(n10184), .Z(o[5418]) );
  AND U15275 ( .A(p_input[25418]), .B(p_input[15418]), .Z(n10184) );
  AND U15276 ( .A(p_input[5418]), .B(p_input[35418]), .Z(n10183) );
  AND U15277 ( .A(n10185), .B(n10186), .Z(o[5417]) );
  AND U15278 ( .A(p_input[25417]), .B(p_input[15417]), .Z(n10186) );
  AND U15279 ( .A(p_input[5417]), .B(p_input[35417]), .Z(n10185) );
  AND U15280 ( .A(n10187), .B(n10188), .Z(o[5416]) );
  AND U15281 ( .A(p_input[25416]), .B(p_input[15416]), .Z(n10188) );
  AND U15282 ( .A(p_input[5416]), .B(p_input[35416]), .Z(n10187) );
  AND U15283 ( .A(n10189), .B(n10190), .Z(o[5415]) );
  AND U15284 ( .A(p_input[25415]), .B(p_input[15415]), .Z(n10190) );
  AND U15285 ( .A(p_input[5415]), .B(p_input[35415]), .Z(n10189) );
  AND U15286 ( .A(n10191), .B(n10192), .Z(o[5414]) );
  AND U15287 ( .A(p_input[25414]), .B(p_input[15414]), .Z(n10192) );
  AND U15288 ( .A(p_input[5414]), .B(p_input[35414]), .Z(n10191) );
  AND U15289 ( .A(n10193), .B(n10194), .Z(o[5413]) );
  AND U15290 ( .A(p_input[25413]), .B(p_input[15413]), .Z(n10194) );
  AND U15291 ( .A(p_input[5413]), .B(p_input[35413]), .Z(n10193) );
  AND U15292 ( .A(n10195), .B(n10196), .Z(o[5412]) );
  AND U15293 ( .A(p_input[25412]), .B(p_input[15412]), .Z(n10196) );
  AND U15294 ( .A(p_input[5412]), .B(p_input[35412]), .Z(n10195) );
  AND U15295 ( .A(n10197), .B(n10198), .Z(o[5411]) );
  AND U15296 ( .A(p_input[25411]), .B(p_input[15411]), .Z(n10198) );
  AND U15297 ( .A(p_input[5411]), .B(p_input[35411]), .Z(n10197) );
  AND U15298 ( .A(n10199), .B(n10200), .Z(o[5410]) );
  AND U15299 ( .A(p_input[25410]), .B(p_input[15410]), .Z(n10200) );
  AND U15300 ( .A(p_input[5410]), .B(p_input[35410]), .Z(n10199) );
  AND U15301 ( .A(n10201), .B(n10202), .Z(o[540]) );
  AND U15302 ( .A(p_input[20540]), .B(p_input[10540]), .Z(n10202) );
  AND U15303 ( .A(p_input[540]), .B(p_input[30540]), .Z(n10201) );
  AND U15304 ( .A(n10203), .B(n10204), .Z(o[5409]) );
  AND U15305 ( .A(p_input[25409]), .B(p_input[15409]), .Z(n10204) );
  AND U15306 ( .A(p_input[5409]), .B(p_input[35409]), .Z(n10203) );
  AND U15307 ( .A(n10205), .B(n10206), .Z(o[5408]) );
  AND U15308 ( .A(p_input[25408]), .B(p_input[15408]), .Z(n10206) );
  AND U15309 ( .A(p_input[5408]), .B(p_input[35408]), .Z(n10205) );
  AND U15310 ( .A(n10207), .B(n10208), .Z(o[5407]) );
  AND U15311 ( .A(p_input[25407]), .B(p_input[15407]), .Z(n10208) );
  AND U15312 ( .A(p_input[5407]), .B(p_input[35407]), .Z(n10207) );
  AND U15313 ( .A(n10209), .B(n10210), .Z(o[5406]) );
  AND U15314 ( .A(p_input[25406]), .B(p_input[15406]), .Z(n10210) );
  AND U15315 ( .A(p_input[5406]), .B(p_input[35406]), .Z(n10209) );
  AND U15316 ( .A(n10211), .B(n10212), .Z(o[5405]) );
  AND U15317 ( .A(p_input[25405]), .B(p_input[15405]), .Z(n10212) );
  AND U15318 ( .A(p_input[5405]), .B(p_input[35405]), .Z(n10211) );
  AND U15319 ( .A(n10213), .B(n10214), .Z(o[5404]) );
  AND U15320 ( .A(p_input[25404]), .B(p_input[15404]), .Z(n10214) );
  AND U15321 ( .A(p_input[5404]), .B(p_input[35404]), .Z(n10213) );
  AND U15322 ( .A(n10215), .B(n10216), .Z(o[5403]) );
  AND U15323 ( .A(p_input[25403]), .B(p_input[15403]), .Z(n10216) );
  AND U15324 ( .A(p_input[5403]), .B(p_input[35403]), .Z(n10215) );
  AND U15325 ( .A(n10217), .B(n10218), .Z(o[5402]) );
  AND U15326 ( .A(p_input[25402]), .B(p_input[15402]), .Z(n10218) );
  AND U15327 ( .A(p_input[5402]), .B(p_input[35402]), .Z(n10217) );
  AND U15328 ( .A(n10219), .B(n10220), .Z(o[5401]) );
  AND U15329 ( .A(p_input[25401]), .B(p_input[15401]), .Z(n10220) );
  AND U15330 ( .A(p_input[5401]), .B(p_input[35401]), .Z(n10219) );
  AND U15331 ( .A(n10221), .B(n10222), .Z(o[5400]) );
  AND U15332 ( .A(p_input[25400]), .B(p_input[15400]), .Z(n10222) );
  AND U15333 ( .A(p_input[5400]), .B(p_input[35400]), .Z(n10221) );
  AND U15334 ( .A(n10223), .B(n10224), .Z(o[53]) );
  AND U15335 ( .A(p_input[20053]), .B(p_input[10053]), .Z(n10224) );
  AND U15336 ( .A(p_input[53]), .B(p_input[30053]), .Z(n10223) );
  AND U15337 ( .A(n10225), .B(n10226), .Z(o[539]) );
  AND U15338 ( .A(p_input[20539]), .B(p_input[10539]), .Z(n10226) );
  AND U15339 ( .A(p_input[539]), .B(p_input[30539]), .Z(n10225) );
  AND U15340 ( .A(n10227), .B(n10228), .Z(o[5399]) );
  AND U15341 ( .A(p_input[25399]), .B(p_input[15399]), .Z(n10228) );
  AND U15342 ( .A(p_input[5399]), .B(p_input[35399]), .Z(n10227) );
  AND U15343 ( .A(n10229), .B(n10230), .Z(o[5398]) );
  AND U15344 ( .A(p_input[25398]), .B(p_input[15398]), .Z(n10230) );
  AND U15345 ( .A(p_input[5398]), .B(p_input[35398]), .Z(n10229) );
  AND U15346 ( .A(n10231), .B(n10232), .Z(o[5397]) );
  AND U15347 ( .A(p_input[25397]), .B(p_input[15397]), .Z(n10232) );
  AND U15348 ( .A(p_input[5397]), .B(p_input[35397]), .Z(n10231) );
  AND U15349 ( .A(n10233), .B(n10234), .Z(o[5396]) );
  AND U15350 ( .A(p_input[25396]), .B(p_input[15396]), .Z(n10234) );
  AND U15351 ( .A(p_input[5396]), .B(p_input[35396]), .Z(n10233) );
  AND U15352 ( .A(n10235), .B(n10236), .Z(o[5395]) );
  AND U15353 ( .A(p_input[25395]), .B(p_input[15395]), .Z(n10236) );
  AND U15354 ( .A(p_input[5395]), .B(p_input[35395]), .Z(n10235) );
  AND U15355 ( .A(n10237), .B(n10238), .Z(o[5394]) );
  AND U15356 ( .A(p_input[25394]), .B(p_input[15394]), .Z(n10238) );
  AND U15357 ( .A(p_input[5394]), .B(p_input[35394]), .Z(n10237) );
  AND U15358 ( .A(n10239), .B(n10240), .Z(o[5393]) );
  AND U15359 ( .A(p_input[25393]), .B(p_input[15393]), .Z(n10240) );
  AND U15360 ( .A(p_input[5393]), .B(p_input[35393]), .Z(n10239) );
  AND U15361 ( .A(n10241), .B(n10242), .Z(o[5392]) );
  AND U15362 ( .A(p_input[25392]), .B(p_input[15392]), .Z(n10242) );
  AND U15363 ( .A(p_input[5392]), .B(p_input[35392]), .Z(n10241) );
  AND U15364 ( .A(n10243), .B(n10244), .Z(o[5391]) );
  AND U15365 ( .A(p_input[25391]), .B(p_input[15391]), .Z(n10244) );
  AND U15366 ( .A(p_input[5391]), .B(p_input[35391]), .Z(n10243) );
  AND U15367 ( .A(n10245), .B(n10246), .Z(o[5390]) );
  AND U15368 ( .A(p_input[25390]), .B(p_input[15390]), .Z(n10246) );
  AND U15369 ( .A(p_input[5390]), .B(p_input[35390]), .Z(n10245) );
  AND U15370 ( .A(n10247), .B(n10248), .Z(o[538]) );
  AND U15371 ( .A(p_input[20538]), .B(p_input[10538]), .Z(n10248) );
  AND U15372 ( .A(p_input[538]), .B(p_input[30538]), .Z(n10247) );
  AND U15373 ( .A(n10249), .B(n10250), .Z(o[5389]) );
  AND U15374 ( .A(p_input[25389]), .B(p_input[15389]), .Z(n10250) );
  AND U15375 ( .A(p_input[5389]), .B(p_input[35389]), .Z(n10249) );
  AND U15376 ( .A(n10251), .B(n10252), .Z(o[5388]) );
  AND U15377 ( .A(p_input[25388]), .B(p_input[15388]), .Z(n10252) );
  AND U15378 ( .A(p_input[5388]), .B(p_input[35388]), .Z(n10251) );
  AND U15379 ( .A(n10253), .B(n10254), .Z(o[5387]) );
  AND U15380 ( .A(p_input[25387]), .B(p_input[15387]), .Z(n10254) );
  AND U15381 ( .A(p_input[5387]), .B(p_input[35387]), .Z(n10253) );
  AND U15382 ( .A(n10255), .B(n10256), .Z(o[5386]) );
  AND U15383 ( .A(p_input[25386]), .B(p_input[15386]), .Z(n10256) );
  AND U15384 ( .A(p_input[5386]), .B(p_input[35386]), .Z(n10255) );
  AND U15385 ( .A(n10257), .B(n10258), .Z(o[5385]) );
  AND U15386 ( .A(p_input[25385]), .B(p_input[15385]), .Z(n10258) );
  AND U15387 ( .A(p_input[5385]), .B(p_input[35385]), .Z(n10257) );
  AND U15388 ( .A(n10259), .B(n10260), .Z(o[5384]) );
  AND U15389 ( .A(p_input[25384]), .B(p_input[15384]), .Z(n10260) );
  AND U15390 ( .A(p_input[5384]), .B(p_input[35384]), .Z(n10259) );
  AND U15391 ( .A(n10261), .B(n10262), .Z(o[5383]) );
  AND U15392 ( .A(p_input[25383]), .B(p_input[15383]), .Z(n10262) );
  AND U15393 ( .A(p_input[5383]), .B(p_input[35383]), .Z(n10261) );
  AND U15394 ( .A(n10263), .B(n10264), .Z(o[5382]) );
  AND U15395 ( .A(p_input[25382]), .B(p_input[15382]), .Z(n10264) );
  AND U15396 ( .A(p_input[5382]), .B(p_input[35382]), .Z(n10263) );
  AND U15397 ( .A(n10265), .B(n10266), .Z(o[5381]) );
  AND U15398 ( .A(p_input[25381]), .B(p_input[15381]), .Z(n10266) );
  AND U15399 ( .A(p_input[5381]), .B(p_input[35381]), .Z(n10265) );
  AND U15400 ( .A(n10267), .B(n10268), .Z(o[5380]) );
  AND U15401 ( .A(p_input[25380]), .B(p_input[15380]), .Z(n10268) );
  AND U15402 ( .A(p_input[5380]), .B(p_input[35380]), .Z(n10267) );
  AND U15403 ( .A(n10269), .B(n10270), .Z(o[537]) );
  AND U15404 ( .A(p_input[20537]), .B(p_input[10537]), .Z(n10270) );
  AND U15405 ( .A(p_input[537]), .B(p_input[30537]), .Z(n10269) );
  AND U15406 ( .A(n10271), .B(n10272), .Z(o[5379]) );
  AND U15407 ( .A(p_input[25379]), .B(p_input[15379]), .Z(n10272) );
  AND U15408 ( .A(p_input[5379]), .B(p_input[35379]), .Z(n10271) );
  AND U15409 ( .A(n10273), .B(n10274), .Z(o[5378]) );
  AND U15410 ( .A(p_input[25378]), .B(p_input[15378]), .Z(n10274) );
  AND U15411 ( .A(p_input[5378]), .B(p_input[35378]), .Z(n10273) );
  AND U15412 ( .A(n10275), .B(n10276), .Z(o[5377]) );
  AND U15413 ( .A(p_input[25377]), .B(p_input[15377]), .Z(n10276) );
  AND U15414 ( .A(p_input[5377]), .B(p_input[35377]), .Z(n10275) );
  AND U15415 ( .A(n10277), .B(n10278), .Z(o[5376]) );
  AND U15416 ( .A(p_input[25376]), .B(p_input[15376]), .Z(n10278) );
  AND U15417 ( .A(p_input[5376]), .B(p_input[35376]), .Z(n10277) );
  AND U15418 ( .A(n10279), .B(n10280), .Z(o[5375]) );
  AND U15419 ( .A(p_input[25375]), .B(p_input[15375]), .Z(n10280) );
  AND U15420 ( .A(p_input[5375]), .B(p_input[35375]), .Z(n10279) );
  AND U15421 ( .A(n10281), .B(n10282), .Z(o[5374]) );
  AND U15422 ( .A(p_input[25374]), .B(p_input[15374]), .Z(n10282) );
  AND U15423 ( .A(p_input[5374]), .B(p_input[35374]), .Z(n10281) );
  AND U15424 ( .A(n10283), .B(n10284), .Z(o[5373]) );
  AND U15425 ( .A(p_input[25373]), .B(p_input[15373]), .Z(n10284) );
  AND U15426 ( .A(p_input[5373]), .B(p_input[35373]), .Z(n10283) );
  AND U15427 ( .A(n10285), .B(n10286), .Z(o[5372]) );
  AND U15428 ( .A(p_input[25372]), .B(p_input[15372]), .Z(n10286) );
  AND U15429 ( .A(p_input[5372]), .B(p_input[35372]), .Z(n10285) );
  AND U15430 ( .A(n10287), .B(n10288), .Z(o[5371]) );
  AND U15431 ( .A(p_input[25371]), .B(p_input[15371]), .Z(n10288) );
  AND U15432 ( .A(p_input[5371]), .B(p_input[35371]), .Z(n10287) );
  AND U15433 ( .A(n10289), .B(n10290), .Z(o[5370]) );
  AND U15434 ( .A(p_input[25370]), .B(p_input[15370]), .Z(n10290) );
  AND U15435 ( .A(p_input[5370]), .B(p_input[35370]), .Z(n10289) );
  AND U15436 ( .A(n10291), .B(n10292), .Z(o[536]) );
  AND U15437 ( .A(p_input[20536]), .B(p_input[10536]), .Z(n10292) );
  AND U15438 ( .A(p_input[536]), .B(p_input[30536]), .Z(n10291) );
  AND U15439 ( .A(n10293), .B(n10294), .Z(o[5369]) );
  AND U15440 ( .A(p_input[25369]), .B(p_input[15369]), .Z(n10294) );
  AND U15441 ( .A(p_input[5369]), .B(p_input[35369]), .Z(n10293) );
  AND U15442 ( .A(n10295), .B(n10296), .Z(o[5368]) );
  AND U15443 ( .A(p_input[25368]), .B(p_input[15368]), .Z(n10296) );
  AND U15444 ( .A(p_input[5368]), .B(p_input[35368]), .Z(n10295) );
  AND U15445 ( .A(n10297), .B(n10298), .Z(o[5367]) );
  AND U15446 ( .A(p_input[25367]), .B(p_input[15367]), .Z(n10298) );
  AND U15447 ( .A(p_input[5367]), .B(p_input[35367]), .Z(n10297) );
  AND U15448 ( .A(n10299), .B(n10300), .Z(o[5366]) );
  AND U15449 ( .A(p_input[25366]), .B(p_input[15366]), .Z(n10300) );
  AND U15450 ( .A(p_input[5366]), .B(p_input[35366]), .Z(n10299) );
  AND U15451 ( .A(n10301), .B(n10302), .Z(o[5365]) );
  AND U15452 ( .A(p_input[25365]), .B(p_input[15365]), .Z(n10302) );
  AND U15453 ( .A(p_input[5365]), .B(p_input[35365]), .Z(n10301) );
  AND U15454 ( .A(n10303), .B(n10304), .Z(o[5364]) );
  AND U15455 ( .A(p_input[25364]), .B(p_input[15364]), .Z(n10304) );
  AND U15456 ( .A(p_input[5364]), .B(p_input[35364]), .Z(n10303) );
  AND U15457 ( .A(n10305), .B(n10306), .Z(o[5363]) );
  AND U15458 ( .A(p_input[25363]), .B(p_input[15363]), .Z(n10306) );
  AND U15459 ( .A(p_input[5363]), .B(p_input[35363]), .Z(n10305) );
  AND U15460 ( .A(n10307), .B(n10308), .Z(o[5362]) );
  AND U15461 ( .A(p_input[25362]), .B(p_input[15362]), .Z(n10308) );
  AND U15462 ( .A(p_input[5362]), .B(p_input[35362]), .Z(n10307) );
  AND U15463 ( .A(n10309), .B(n10310), .Z(o[5361]) );
  AND U15464 ( .A(p_input[25361]), .B(p_input[15361]), .Z(n10310) );
  AND U15465 ( .A(p_input[5361]), .B(p_input[35361]), .Z(n10309) );
  AND U15466 ( .A(n10311), .B(n10312), .Z(o[5360]) );
  AND U15467 ( .A(p_input[25360]), .B(p_input[15360]), .Z(n10312) );
  AND U15468 ( .A(p_input[5360]), .B(p_input[35360]), .Z(n10311) );
  AND U15469 ( .A(n10313), .B(n10314), .Z(o[535]) );
  AND U15470 ( .A(p_input[20535]), .B(p_input[10535]), .Z(n10314) );
  AND U15471 ( .A(p_input[535]), .B(p_input[30535]), .Z(n10313) );
  AND U15472 ( .A(n10315), .B(n10316), .Z(o[5359]) );
  AND U15473 ( .A(p_input[25359]), .B(p_input[15359]), .Z(n10316) );
  AND U15474 ( .A(p_input[5359]), .B(p_input[35359]), .Z(n10315) );
  AND U15475 ( .A(n10317), .B(n10318), .Z(o[5358]) );
  AND U15476 ( .A(p_input[25358]), .B(p_input[15358]), .Z(n10318) );
  AND U15477 ( .A(p_input[5358]), .B(p_input[35358]), .Z(n10317) );
  AND U15478 ( .A(n10319), .B(n10320), .Z(o[5357]) );
  AND U15479 ( .A(p_input[25357]), .B(p_input[15357]), .Z(n10320) );
  AND U15480 ( .A(p_input[5357]), .B(p_input[35357]), .Z(n10319) );
  AND U15481 ( .A(n10321), .B(n10322), .Z(o[5356]) );
  AND U15482 ( .A(p_input[25356]), .B(p_input[15356]), .Z(n10322) );
  AND U15483 ( .A(p_input[5356]), .B(p_input[35356]), .Z(n10321) );
  AND U15484 ( .A(n10323), .B(n10324), .Z(o[5355]) );
  AND U15485 ( .A(p_input[25355]), .B(p_input[15355]), .Z(n10324) );
  AND U15486 ( .A(p_input[5355]), .B(p_input[35355]), .Z(n10323) );
  AND U15487 ( .A(n10325), .B(n10326), .Z(o[5354]) );
  AND U15488 ( .A(p_input[25354]), .B(p_input[15354]), .Z(n10326) );
  AND U15489 ( .A(p_input[5354]), .B(p_input[35354]), .Z(n10325) );
  AND U15490 ( .A(n10327), .B(n10328), .Z(o[5353]) );
  AND U15491 ( .A(p_input[25353]), .B(p_input[15353]), .Z(n10328) );
  AND U15492 ( .A(p_input[5353]), .B(p_input[35353]), .Z(n10327) );
  AND U15493 ( .A(n10329), .B(n10330), .Z(o[5352]) );
  AND U15494 ( .A(p_input[25352]), .B(p_input[15352]), .Z(n10330) );
  AND U15495 ( .A(p_input[5352]), .B(p_input[35352]), .Z(n10329) );
  AND U15496 ( .A(n10331), .B(n10332), .Z(o[5351]) );
  AND U15497 ( .A(p_input[25351]), .B(p_input[15351]), .Z(n10332) );
  AND U15498 ( .A(p_input[5351]), .B(p_input[35351]), .Z(n10331) );
  AND U15499 ( .A(n10333), .B(n10334), .Z(o[5350]) );
  AND U15500 ( .A(p_input[25350]), .B(p_input[15350]), .Z(n10334) );
  AND U15501 ( .A(p_input[5350]), .B(p_input[35350]), .Z(n10333) );
  AND U15502 ( .A(n10335), .B(n10336), .Z(o[534]) );
  AND U15503 ( .A(p_input[20534]), .B(p_input[10534]), .Z(n10336) );
  AND U15504 ( .A(p_input[534]), .B(p_input[30534]), .Z(n10335) );
  AND U15505 ( .A(n10337), .B(n10338), .Z(o[5349]) );
  AND U15506 ( .A(p_input[25349]), .B(p_input[15349]), .Z(n10338) );
  AND U15507 ( .A(p_input[5349]), .B(p_input[35349]), .Z(n10337) );
  AND U15508 ( .A(n10339), .B(n10340), .Z(o[5348]) );
  AND U15509 ( .A(p_input[25348]), .B(p_input[15348]), .Z(n10340) );
  AND U15510 ( .A(p_input[5348]), .B(p_input[35348]), .Z(n10339) );
  AND U15511 ( .A(n10341), .B(n10342), .Z(o[5347]) );
  AND U15512 ( .A(p_input[25347]), .B(p_input[15347]), .Z(n10342) );
  AND U15513 ( .A(p_input[5347]), .B(p_input[35347]), .Z(n10341) );
  AND U15514 ( .A(n10343), .B(n10344), .Z(o[5346]) );
  AND U15515 ( .A(p_input[25346]), .B(p_input[15346]), .Z(n10344) );
  AND U15516 ( .A(p_input[5346]), .B(p_input[35346]), .Z(n10343) );
  AND U15517 ( .A(n10345), .B(n10346), .Z(o[5345]) );
  AND U15518 ( .A(p_input[25345]), .B(p_input[15345]), .Z(n10346) );
  AND U15519 ( .A(p_input[5345]), .B(p_input[35345]), .Z(n10345) );
  AND U15520 ( .A(n10347), .B(n10348), .Z(o[5344]) );
  AND U15521 ( .A(p_input[25344]), .B(p_input[15344]), .Z(n10348) );
  AND U15522 ( .A(p_input[5344]), .B(p_input[35344]), .Z(n10347) );
  AND U15523 ( .A(n10349), .B(n10350), .Z(o[5343]) );
  AND U15524 ( .A(p_input[25343]), .B(p_input[15343]), .Z(n10350) );
  AND U15525 ( .A(p_input[5343]), .B(p_input[35343]), .Z(n10349) );
  AND U15526 ( .A(n10351), .B(n10352), .Z(o[5342]) );
  AND U15527 ( .A(p_input[25342]), .B(p_input[15342]), .Z(n10352) );
  AND U15528 ( .A(p_input[5342]), .B(p_input[35342]), .Z(n10351) );
  AND U15529 ( .A(n10353), .B(n10354), .Z(o[5341]) );
  AND U15530 ( .A(p_input[25341]), .B(p_input[15341]), .Z(n10354) );
  AND U15531 ( .A(p_input[5341]), .B(p_input[35341]), .Z(n10353) );
  AND U15532 ( .A(n10355), .B(n10356), .Z(o[5340]) );
  AND U15533 ( .A(p_input[25340]), .B(p_input[15340]), .Z(n10356) );
  AND U15534 ( .A(p_input[5340]), .B(p_input[35340]), .Z(n10355) );
  AND U15535 ( .A(n10357), .B(n10358), .Z(o[533]) );
  AND U15536 ( .A(p_input[20533]), .B(p_input[10533]), .Z(n10358) );
  AND U15537 ( .A(p_input[533]), .B(p_input[30533]), .Z(n10357) );
  AND U15538 ( .A(n10359), .B(n10360), .Z(o[5339]) );
  AND U15539 ( .A(p_input[25339]), .B(p_input[15339]), .Z(n10360) );
  AND U15540 ( .A(p_input[5339]), .B(p_input[35339]), .Z(n10359) );
  AND U15541 ( .A(n10361), .B(n10362), .Z(o[5338]) );
  AND U15542 ( .A(p_input[25338]), .B(p_input[15338]), .Z(n10362) );
  AND U15543 ( .A(p_input[5338]), .B(p_input[35338]), .Z(n10361) );
  AND U15544 ( .A(n10363), .B(n10364), .Z(o[5337]) );
  AND U15545 ( .A(p_input[25337]), .B(p_input[15337]), .Z(n10364) );
  AND U15546 ( .A(p_input[5337]), .B(p_input[35337]), .Z(n10363) );
  AND U15547 ( .A(n10365), .B(n10366), .Z(o[5336]) );
  AND U15548 ( .A(p_input[25336]), .B(p_input[15336]), .Z(n10366) );
  AND U15549 ( .A(p_input[5336]), .B(p_input[35336]), .Z(n10365) );
  AND U15550 ( .A(n10367), .B(n10368), .Z(o[5335]) );
  AND U15551 ( .A(p_input[25335]), .B(p_input[15335]), .Z(n10368) );
  AND U15552 ( .A(p_input[5335]), .B(p_input[35335]), .Z(n10367) );
  AND U15553 ( .A(n10369), .B(n10370), .Z(o[5334]) );
  AND U15554 ( .A(p_input[25334]), .B(p_input[15334]), .Z(n10370) );
  AND U15555 ( .A(p_input[5334]), .B(p_input[35334]), .Z(n10369) );
  AND U15556 ( .A(n10371), .B(n10372), .Z(o[5333]) );
  AND U15557 ( .A(p_input[25333]), .B(p_input[15333]), .Z(n10372) );
  AND U15558 ( .A(p_input[5333]), .B(p_input[35333]), .Z(n10371) );
  AND U15559 ( .A(n10373), .B(n10374), .Z(o[5332]) );
  AND U15560 ( .A(p_input[25332]), .B(p_input[15332]), .Z(n10374) );
  AND U15561 ( .A(p_input[5332]), .B(p_input[35332]), .Z(n10373) );
  AND U15562 ( .A(n10375), .B(n10376), .Z(o[5331]) );
  AND U15563 ( .A(p_input[25331]), .B(p_input[15331]), .Z(n10376) );
  AND U15564 ( .A(p_input[5331]), .B(p_input[35331]), .Z(n10375) );
  AND U15565 ( .A(n10377), .B(n10378), .Z(o[5330]) );
  AND U15566 ( .A(p_input[25330]), .B(p_input[15330]), .Z(n10378) );
  AND U15567 ( .A(p_input[5330]), .B(p_input[35330]), .Z(n10377) );
  AND U15568 ( .A(n10379), .B(n10380), .Z(o[532]) );
  AND U15569 ( .A(p_input[20532]), .B(p_input[10532]), .Z(n10380) );
  AND U15570 ( .A(p_input[532]), .B(p_input[30532]), .Z(n10379) );
  AND U15571 ( .A(n10381), .B(n10382), .Z(o[5329]) );
  AND U15572 ( .A(p_input[25329]), .B(p_input[15329]), .Z(n10382) );
  AND U15573 ( .A(p_input[5329]), .B(p_input[35329]), .Z(n10381) );
  AND U15574 ( .A(n10383), .B(n10384), .Z(o[5328]) );
  AND U15575 ( .A(p_input[25328]), .B(p_input[15328]), .Z(n10384) );
  AND U15576 ( .A(p_input[5328]), .B(p_input[35328]), .Z(n10383) );
  AND U15577 ( .A(n10385), .B(n10386), .Z(o[5327]) );
  AND U15578 ( .A(p_input[25327]), .B(p_input[15327]), .Z(n10386) );
  AND U15579 ( .A(p_input[5327]), .B(p_input[35327]), .Z(n10385) );
  AND U15580 ( .A(n10387), .B(n10388), .Z(o[5326]) );
  AND U15581 ( .A(p_input[25326]), .B(p_input[15326]), .Z(n10388) );
  AND U15582 ( .A(p_input[5326]), .B(p_input[35326]), .Z(n10387) );
  AND U15583 ( .A(n10389), .B(n10390), .Z(o[5325]) );
  AND U15584 ( .A(p_input[25325]), .B(p_input[15325]), .Z(n10390) );
  AND U15585 ( .A(p_input[5325]), .B(p_input[35325]), .Z(n10389) );
  AND U15586 ( .A(n10391), .B(n10392), .Z(o[5324]) );
  AND U15587 ( .A(p_input[25324]), .B(p_input[15324]), .Z(n10392) );
  AND U15588 ( .A(p_input[5324]), .B(p_input[35324]), .Z(n10391) );
  AND U15589 ( .A(n10393), .B(n10394), .Z(o[5323]) );
  AND U15590 ( .A(p_input[25323]), .B(p_input[15323]), .Z(n10394) );
  AND U15591 ( .A(p_input[5323]), .B(p_input[35323]), .Z(n10393) );
  AND U15592 ( .A(n10395), .B(n10396), .Z(o[5322]) );
  AND U15593 ( .A(p_input[25322]), .B(p_input[15322]), .Z(n10396) );
  AND U15594 ( .A(p_input[5322]), .B(p_input[35322]), .Z(n10395) );
  AND U15595 ( .A(n10397), .B(n10398), .Z(o[5321]) );
  AND U15596 ( .A(p_input[25321]), .B(p_input[15321]), .Z(n10398) );
  AND U15597 ( .A(p_input[5321]), .B(p_input[35321]), .Z(n10397) );
  AND U15598 ( .A(n10399), .B(n10400), .Z(o[5320]) );
  AND U15599 ( .A(p_input[25320]), .B(p_input[15320]), .Z(n10400) );
  AND U15600 ( .A(p_input[5320]), .B(p_input[35320]), .Z(n10399) );
  AND U15601 ( .A(n10401), .B(n10402), .Z(o[531]) );
  AND U15602 ( .A(p_input[20531]), .B(p_input[10531]), .Z(n10402) );
  AND U15603 ( .A(p_input[531]), .B(p_input[30531]), .Z(n10401) );
  AND U15604 ( .A(n10403), .B(n10404), .Z(o[5319]) );
  AND U15605 ( .A(p_input[25319]), .B(p_input[15319]), .Z(n10404) );
  AND U15606 ( .A(p_input[5319]), .B(p_input[35319]), .Z(n10403) );
  AND U15607 ( .A(n10405), .B(n10406), .Z(o[5318]) );
  AND U15608 ( .A(p_input[25318]), .B(p_input[15318]), .Z(n10406) );
  AND U15609 ( .A(p_input[5318]), .B(p_input[35318]), .Z(n10405) );
  AND U15610 ( .A(n10407), .B(n10408), .Z(o[5317]) );
  AND U15611 ( .A(p_input[25317]), .B(p_input[15317]), .Z(n10408) );
  AND U15612 ( .A(p_input[5317]), .B(p_input[35317]), .Z(n10407) );
  AND U15613 ( .A(n10409), .B(n10410), .Z(o[5316]) );
  AND U15614 ( .A(p_input[25316]), .B(p_input[15316]), .Z(n10410) );
  AND U15615 ( .A(p_input[5316]), .B(p_input[35316]), .Z(n10409) );
  AND U15616 ( .A(n10411), .B(n10412), .Z(o[5315]) );
  AND U15617 ( .A(p_input[25315]), .B(p_input[15315]), .Z(n10412) );
  AND U15618 ( .A(p_input[5315]), .B(p_input[35315]), .Z(n10411) );
  AND U15619 ( .A(n10413), .B(n10414), .Z(o[5314]) );
  AND U15620 ( .A(p_input[25314]), .B(p_input[15314]), .Z(n10414) );
  AND U15621 ( .A(p_input[5314]), .B(p_input[35314]), .Z(n10413) );
  AND U15622 ( .A(n10415), .B(n10416), .Z(o[5313]) );
  AND U15623 ( .A(p_input[25313]), .B(p_input[15313]), .Z(n10416) );
  AND U15624 ( .A(p_input[5313]), .B(p_input[35313]), .Z(n10415) );
  AND U15625 ( .A(n10417), .B(n10418), .Z(o[5312]) );
  AND U15626 ( .A(p_input[25312]), .B(p_input[15312]), .Z(n10418) );
  AND U15627 ( .A(p_input[5312]), .B(p_input[35312]), .Z(n10417) );
  AND U15628 ( .A(n10419), .B(n10420), .Z(o[5311]) );
  AND U15629 ( .A(p_input[25311]), .B(p_input[15311]), .Z(n10420) );
  AND U15630 ( .A(p_input[5311]), .B(p_input[35311]), .Z(n10419) );
  AND U15631 ( .A(n10421), .B(n10422), .Z(o[5310]) );
  AND U15632 ( .A(p_input[25310]), .B(p_input[15310]), .Z(n10422) );
  AND U15633 ( .A(p_input[5310]), .B(p_input[35310]), .Z(n10421) );
  AND U15634 ( .A(n10423), .B(n10424), .Z(o[530]) );
  AND U15635 ( .A(p_input[20530]), .B(p_input[10530]), .Z(n10424) );
  AND U15636 ( .A(p_input[530]), .B(p_input[30530]), .Z(n10423) );
  AND U15637 ( .A(n10425), .B(n10426), .Z(o[5309]) );
  AND U15638 ( .A(p_input[25309]), .B(p_input[15309]), .Z(n10426) );
  AND U15639 ( .A(p_input[5309]), .B(p_input[35309]), .Z(n10425) );
  AND U15640 ( .A(n10427), .B(n10428), .Z(o[5308]) );
  AND U15641 ( .A(p_input[25308]), .B(p_input[15308]), .Z(n10428) );
  AND U15642 ( .A(p_input[5308]), .B(p_input[35308]), .Z(n10427) );
  AND U15643 ( .A(n10429), .B(n10430), .Z(o[5307]) );
  AND U15644 ( .A(p_input[25307]), .B(p_input[15307]), .Z(n10430) );
  AND U15645 ( .A(p_input[5307]), .B(p_input[35307]), .Z(n10429) );
  AND U15646 ( .A(n10431), .B(n10432), .Z(o[5306]) );
  AND U15647 ( .A(p_input[25306]), .B(p_input[15306]), .Z(n10432) );
  AND U15648 ( .A(p_input[5306]), .B(p_input[35306]), .Z(n10431) );
  AND U15649 ( .A(n10433), .B(n10434), .Z(o[5305]) );
  AND U15650 ( .A(p_input[25305]), .B(p_input[15305]), .Z(n10434) );
  AND U15651 ( .A(p_input[5305]), .B(p_input[35305]), .Z(n10433) );
  AND U15652 ( .A(n10435), .B(n10436), .Z(o[5304]) );
  AND U15653 ( .A(p_input[25304]), .B(p_input[15304]), .Z(n10436) );
  AND U15654 ( .A(p_input[5304]), .B(p_input[35304]), .Z(n10435) );
  AND U15655 ( .A(n10437), .B(n10438), .Z(o[5303]) );
  AND U15656 ( .A(p_input[25303]), .B(p_input[15303]), .Z(n10438) );
  AND U15657 ( .A(p_input[5303]), .B(p_input[35303]), .Z(n10437) );
  AND U15658 ( .A(n10439), .B(n10440), .Z(o[5302]) );
  AND U15659 ( .A(p_input[25302]), .B(p_input[15302]), .Z(n10440) );
  AND U15660 ( .A(p_input[5302]), .B(p_input[35302]), .Z(n10439) );
  AND U15661 ( .A(n10441), .B(n10442), .Z(o[5301]) );
  AND U15662 ( .A(p_input[25301]), .B(p_input[15301]), .Z(n10442) );
  AND U15663 ( .A(p_input[5301]), .B(p_input[35301]), .Z(n10441) );
  AND U15664 ( .A(n10443), .B(n10444), .Z(o[5300]) );
  AND U15665 ( .A(p_input[25300]), .B(p_input[15300]), .Z(n10444) );
  AND U15666 ( .A(p_input[5300]), .B(p_input[35300]), .Z(n10443) );
  AND U15667 ( .A(n10445), .B(n10446), .Z(o[52]) );
  AND U15668 ( .A(p_input[20052]), .B(p_input[10052]), .Z(n10446) );
  AND U15669 ( .A(p_input[52]), .B(p_input[30052]), .Z(n10445) );
  AND U15670 ( .A(n10447), .B(n10448), .Z(o[529]) );
  AND U15671 ( .A(p_input[20529]), .B(p_input[10529]), .Z(n10448) );
  AND U15672 ( .A(p_input[529]), .B(p_input[30529]), .Z(n10447) );
  AND U15673 ( .A(n10449), .B(n10450), .Z(o[5299]) );
  AND U15674 ( .A(p_input[25299]), .B(p_input[15299]), .Z(n10450) );
  AND U15675 ( .A(p_input[5299]), .B(p_input[35299]), .Z(n10449) );
  AND U15676 ( .A(n10451), .B(n10452), .Z(o[5298]) );
  AND U15677 ( .A(p_input[25298]), .B(p_input[15298]), .Z(n10452) );
  AND U15678 ( .A(p_input[5298]), .B(p_input[35298]), .Z(n10451) );
  AND U15679 ( .A(n10453), .B(n10454), .Z(o[5297]) );
  AND U15680 ( .A(p_input[25297]), .B(p_input[15297]), .Z(n10454) );
  AND U15681 ( .A(p_input[5297]), .B(p_input[35297]), .Z(n10453) );
  AND U15682 ( .A(n10455), .B(n10456), .Z(o[5296]) );
  AND U15683 ( .A(p_input[25296]), .B(p_input[15296]), .Z(n10456) );
  AND U15684 ( .A(p_input[5296]), .B(p_input[35296]), .Z(n10455) );
  AND U15685 ( .A(n10457), .B(n10458), .Z(o[5295]) );
  AND U15686 ( .A(p_input[25295]), .B(p_input[15295]), .Z(n10458) );
  AND U15687 ( .A(p_input[5295]), .B(p_input[35295]), .Z(n10457) );
  AND U15688 ( .A(n10459), .B(n10460), .Z(o[5294]) );
  AND U15689 ( .A(p_input[25294]), .B(p_input[15294]), .Z(n10460) );
  AND U15690 ( .A(p_input[5294]), .B(p_input[35294]), .Z(n10459) );
  AND U15691 ( .A(n10461), .B(n10462), .Z(o[5293]) );
  AND U15692 ( .A(p_input[25293]), .B(p_input[15293]), .Z(n10462) );
  AND U15693 ( .A(p_input[5293]), .B(p_input[35293]), .Z(n10461) );
  AND U15694 ( .A(n10463), .B(n10464), .Z(o[5292]) );
  AND U15695 ( .A(p_input[25292]), .B(p_input[15292]), .Z(n10464) );
  AND U15696 ( .A(p_input[5292]), .B(p_input[35292]), .Z(n10463) );
  AND U15697 ( .A(n10465), .B(n10466), .Z(o[5291]) );
  AND U15698 ( .A(p_input[25291]), .B(p_input[15291]), .Z(n10466) );
  AND U15699 ( .A(p_input[5291]), .B(p_input[35291]), .Z(n10465) );
  AND U15700 ( .A(n10467), .B(n10468), .Z(o[5290]) );
  AND U15701 ( .A(p_input[25290]), .B(p_input[15290]), .Z(n10468) );
  AND U15702 ( .A(p_input[5290]), .B(p_input[35290]), .Z(n10467) );
  AND U15703 ( .A(n10469), .B(n10470), .Z(o[528]) );
  AND U15704 ( .A(p_input[20528]), .B(p_input[10528]), .Z(n10470) );
  AND U15705 ( .A(p_input[528]), .B(p_input[30528]), .Z(n10469) );
  AND U15706 ( .A(n10471), .B(n10472), .Z(o[5289]) );
  AND U15707 ( .A(p_input[25289]), .B(p_input[15289]), .Z(n10472) );
  AND U15708 ( .A(p_input[5289]), .B(p_input[35289]), .Z(n10471) );
  AND U15709 ( .A(n10473), .B(n10474), .Z(o[5288]) );
  AND U15710 ( .A(p_input[25288]), .B(p_input[15288]), .Z(n10474) );
  AND U15711 ( .A(p_input[5288]), .B(p_input[35288]), .Z(n10473) );
  AND U15712 ( .A(n10475), .B(n10476), .Z(o[5287]) );
  AND U15713 ( .A(p_input[25287]), .B(p_input[15287]), .Z(n10476) );
  AND U15714 ( .A(p_input[5287]), .B(p_input[35287]), .Z(n10475) );
  AND U15715 ( .A(n10477), .B(n10478), .Z(o[5286]) );
  AND U15716 ( .A(p_input[25286]), .B(p_input[15286]), .Z(n10478) );
  AND U15717 ( .A(p_input[5286]), .B(p_input[35286]), .Z(n10477) );
  AND U15718 ( .A(n10479), .B(n10480), .Z(o[5285]) );
  AND U15719 ( .A(p_input[25285]), .B(p_input[15285]), .Z(n10480) );
  AND U15720 ( .A(p_input[5285]), .B(p_input[35285]), .Z(n10479) );
  AND U15721 ( .A(n10481), .B(n10482), .Z(o[5284]) );
  AND U15722 ( .A(p_input[25284]), .B(p_input[15284]), .Z(n10482) );
  AND U15723 ( .A(p_input[5284]), .B(p_input[35284]), .Z(n10481) );
  AND U15724 ( .A(n10483), .B(n10484), .Z(o[5283]) );
  AND U15725 ( .A(p_input[25283]), .B(p_input[15283]), .Z(n10484) );
  AND U15726 ( .A(p_input[5283]), .B(p_input[35283]), .Z(n10483) );
  AND U15727 ( .A(n10485), .B(n10486), .Z(o[5282]) );
  AND U15728 ( .A(p_input[25282]), .B(p_input[15282]), .Z(n10486) );
  AND U15729 ( .A(p_input[5282]), .B(p_input[35282]), .Z(n10485) );
  AND U15730 ( .A(n10487), .B(n10488), .Z(o[5281]) );
  AND U15731 ( .A(p_input[25281]), .B(p_input[15281]), .Z(n10488) );
  AND U15732 ( .A(p_input[5281]), .B(p_input[35281]), .Z(n10487) );
  AND U15733 ( .A(n10489), .B(n10490), .Z(o[5280]) );
  AND U15734 ( .A(p_input[25280]), .B(p_input[15280]), .Z(n10490) );
  AND U15735 ( .A(p_input[5280]), .B(p_input[35280]), .Z(n10489) );
  AND U15736 ( .A(n10491), .B(n10492), .Z(o[527]) );
  AND U15737 ( .A(p_input[20527]), .B(p_input[10527]), .Z(n10492) );
  AND U15738 ( .A(p_input[527]), .B(p_input[30527]), .Z(n10491) );
  AND U15739 ( .A(n10493), .B(n10494), .Z(o[5279]) );
  AND U15740 ( .A(p_input[25279]), .B(p_input[15279]), .Z(n10494) );
  AND U15741 ( .A(p_input[5279]), .B(p_input[35279]), .Z(n10493) );
  AND U15742 ( .A(n10495), .B(n10496), .Z(o[5278]) );
  AND U15743 ( .A(p_input[25278]), .B(p_input[15278]), .Z(n10496) );
  AND U15744 ( .A(p_input[5278]), .B(p_input[35278]), .Z(n10495) );
  AND U15745 ( .A(n10497), .B(n10498), .Z(o[5277]) );
  AND U15746 ( .A(p_input[25277]), .B(p_input[15277]), .Z(n10498) );
  AND U15747 ( .A(p_input[5277]), .B(p_input[35277]), .Z(n10497) );
  AND U15748 ( .A(n10499), .B(n10500), .Z(o[5276]) );
  AND U15749 ( .A(p_input[25276]), .B(p_input[15276]), .Z(n10500) );
  AND U15750 ( .A(p_input[5276]), .B(p_input[35276]), .Z(n10499) );
  AND U15751 ( .A(n10501), .B(n10502), .Z(o[5275]) );
  AND U15752 ( .A(p_input[25275]), .B(p_input[15275]), .Z(n10502) );
  AND U15753 ( .A(p_input[5275]), .B(p_input[35275]), .Z(n10501) );
  AND U15754 ( .A(n10503), .B(n10504), .Z(o[5274]) );
  AND U15755 ( .A(p_input[25274]), .B(p_input[15274]), .Z(n10504) );
  AND U15756 ( .A(p_input[5274]), .B(p_input[35274]), .Z(n10503) );
  AND U15757 ( .A(n10505), .B(n10506), .Z(o[5273]) );
  AND U15758 ( .A(p_input[25273]), .B(p_input[15273]), .Z(n10506) );
  AND U15759 ( .A(p_input[5273]), .B(p_input[35273]), .Z(n10505) );
  AND U15760 ( .A(n10507), .B(n10508), .Z(o[5272]) );
  AND U15761 ( .A(p_input[25272]), .B(p_input[15272]), .Z(n10508) );
  AND U15762 ( .A(p_input[5272]), .B(p_input[35272]), .Z(n10507) );
  AND U15763 ( .A(n10509), .B(n10510), .Z(o[5271]) );
  AND U15764 ( .A(p_input[25271]), .B(p_input[15271]), .Z(n10510) );
  AND U15765 ( .A(p_input[5271]), .B(p_input[35271]), .Z(n10509) );
  AND U15766 ( .A(n10511), .B(n10512), .Z(o[5270]) );
  AND U15767 ( .A(p_input[25270]), .B(p_input[15270]), .Z(n10512) );
  AND U15768 ( .A(p_input[5270]), .B(p_input[35270]), .Z(n10511) );
  AND U15769 ( .A(n10513), .B(n10514), .Z(o[526]) );
  AND U15770 ( .A(p_input[20526]), .B(p_input[10526]), .Z(n10514) );
  AND U15771 ( .A(p_input[526]), .B(p_input[30526]), .Z(n10513) );
  AND U15772 ( .A(n10515), .B(n10516), .Z(o[5269]) );
  AND U15773 ( .A(p_input[25269]), .B(p_input[15269]), .Z(n10516) );
  AND U15774 ( .A(p_input[5269]), .B(p_input[35269]), .Z(n10515) );
  AND U15775 ( .A(n10517), .B(n10518), .Z(o[5268]) );
  AND U15776 ( .A(p_input[25268]), .B(p_input[15268]), .Z(n10518) );
  AND U15777 ( .A(p_input[5268]), .B(p_input[35268]), .Z(n10517) );
  AND U15778 ( .A(n10519), .B(n10520), .Z(o[5267]) );
  AND U15779 ( .A(p_input[25267]), .B(p_input[15267]), .Z(n10520) );
  AND U15780 ( .A(p_input[5267]), .B(p_input[35267]), .Z(n10519) );
  AND U15781 ( .A(n10521), .B(n10522), .Z(o[5266]) );
  AND U15782 ( .A(p_input[25266]), .B(p_input[15266]), .Z(n10522) );
  AND U15783 ( .A(p_input[5266]), .B(p_input[35266]), .Z(n10521) );
  AND U15784 ( .A(n10523), .B(n10524), .Z(o[5265]) );
  AND U15785 ( .A(p_input[25265]), .B(p_input[15265]), .Z(n10524) );
  AND U15786 ( .A(p_input[5265]), .B(p_input[35265]), .Z(n10523) );
  AND U15787 ( .A(n10525), .B(n10526), .Z(o[5264]) );
  AND U15788 ( .A(p_input[25264]), .B(p_input[15264]), .Z(n10526) );
  AND U15789 ( .A(p_input[5264]), .B(p_input[35264]), .Z(n10525) );
  AND U15790 ( .A(n10527), .B(n10528), .Z(o[5263]) );
  AND U15791 ( .A(p_input[25263]), .B(p_input[15263]), .Z(n10528) );
  AND U15792 ( .A(p_input[5263]), .B(p_input[35263]), .Z(n10527) );
  AND U15793 ( .A(n10529), .B(n10530), .Z(o[5262]) );
  AND U15794 ( .A(p_input[25262]), .B(p_input[15262]), .Z(n10530) );
  AND U15795 ( .A(p_input[5262]), .B(p_input[35262]), .Z(n10529) );
  AND U15796 ( .A(n10531), .B(n10532), .Z(o[5261]) );
  AND U15797 ( .A(p_input[25261]), .B(p_input[15261]), .Z(n10532) );
  AND U15798 ( .A(p_input[5261]), .B(p_input[35261]), .Z(n10531) );
  AND U15799 ( .A(n10533), .B(n10534), .Z(o[5260]) );
  AND U15800 ( .A(p_input[25260]), .B(p_input[15260]), .Z(n10534) );
  AND U15801 ( .A(p_input[5260]), .B(p_input[35260]), .Z(n10533) );
  AND U15802 ( .A(n10535), .B(n10536), .Z(o[525]) );
  AND U15803 ( .A(p_input[20525]), .B(p_input[10525]), .Z(n10536) );
  AND U15804 ( .A(p_input[525]), .B(p_input[30525]), .Z(n10535) );
  AND U15805 ( .A(n10537), .B(n10538), .Z(o[5259]) );
  AND U15806 ( .A(p_input[25259]), .B(p_input[15259]), .Z(n10538) );
  AND U15807 ( .A(p_input[5259]), .B(p_input[35259]), .Z(n10537) );
  AND U15808 ( .A(n10539), .B(n10540), .Z(o[5258]) );
  AND U15809 ( .A(p_input[25258]), .B(p_input[15258]), .Z(n10540) );
  AND U15810 ( .A(p_input[5258]), .B(p_input[35258]), .Z(n10539) );
  AND U15811 ( .A(n10541), .B(n10542), .Z(o[5257]) );
  AND U15812 ( .A(p_input[25257]), .B(p_input[15257]), .Z(n10542) );
  AND U15813 ( .A(p_input[5257]), .B(p_input[35257]), .Z(n10541) );
  AND U15814 ( .A(n10543), .B(n10544), .Z(o[5256]) );
  AND U15815 ( .A(p_input[25256]), .B(p_input[15256]), .Z(n10544) );
  AND U15816 ( .A(p_input[5256]), .B(p_input[35256]), .Z(n10543) );
  AND U15817 ( .A(n10545), .B(n10546), .Z(o[5255]) );
  AND U15818 ( .A(p_input[25255]), .B(p_input[15255]), .Z(n10546) );
  AND U15819 ( .A(p_input[5255]), .B(p_input[35255]), .Z(n10545) );
  AND U15820 ( .A(n10547), .B(n10548), .Z(o[5254]) );
  AND U15821 ( .A(p_input[25254]), .B(p_input[15254]), .Z(n10548) );
  AND U15822 ( .A(p_input[5254]), .B(p_input[35254]), .Z(n10547) );
  AND U15823 ( .A(n10549), .B(n10550), .Z(o[5253]) );
  AND U15824 ( .A(p_input[25253]), .B(p_input[15253]), .Z(n10550) );
  AND U15825 ( .A(p_input[5253]), .B(p_input[35253]), .Z(n10549) );
  AND U15826 ( .A(n10551), .B(n10552), .Z(o[5252]) );
  AND U15827 ( .A(p_input[25252]), .B(p_input[15252]), .Z(n10552) );
  AND U15828 ( .A(p_input[5252]), .B(p_input[35252]), .Z(n10551) );
  AND U15829 ( .A(n10553), .B(n10554), .Z(o[5251]) );
  AND U15830 ( .A(p_input[25251]), .B(p_input[15251]), .Z(n10554) );
  AND U15831 ( .A(p_input[5251]), .B(p_input[35251]), .Z(n10553) );
  AND U15832 ( .A(n10555), .B(n10556), .Z(o[5250]) );
  AND U15833 ( .A(p_input[25250]), .B(p_input[15250]), .Z(n10556) );
  AND U15834 ( .A(p_input[5250]), .B(p_input[35250]), .Z(n10555) );
  AND U15835 ( .A(n10557), .B(n10558), .Z(o[524]) );
  AND U15836 ( .A(p_input[20524]), .B(p_input[10524]), .Z(n10558) );
  AND U15837 ( .A(p_input[524]), .B(p_input[30524]), .Z(n10557) );
  AND U15838 ( .A(n10559), .B(n10560), .Z(o[5249]) );
  AND U15839 ( .A(p_input[25249]), .B(p_input[15249]), .Z(n10560) );
  AND U15840 ( .A(p_input[5249]), .B(p_input[35249]), .Z(n10559) );
  AND U15841 ( .A(n10561), .B(n10562), .Z(o[5248]) );
  AND U15842 ( .A(p_input[25248]), .B(p_input[15248]), .Z(n10562) );
  AND U15843 ( .A(p_input[5248]), .B(p_input[35248]), .Z(n10561) );
  AND U15844 ( .A(n10563), .B(n10564), .Z(o[5247]) );
  AND U15845 ( .A(p_input[25247]), .B(p_input[15247]), .Z(n10564) );
  AND U15846 ( .A(p_input[5247]), .B(p_input[35247]), .Z(n10563) );
  AND U15847 ( .A(n10565), .B(n10566), .Z(o[5246]) );
  AND U15848 ( .A(p_input[25246]), .B(p_input[15246]), .Z(n10566) );
  AND U15849 ( .A(p_input[5246]), .B(p_input[35246]), .Z(n10565) );
  AND U15850 ( .A(n10567), .B(n10568), .Z(o[5245]) );
  AND U15851 ( .A(p_input[25245]), .B(p_input[15245]), .Z(n10568) );
  AND U15852 ( .A(p_input[5245]), .B(p_input[35245]), .Z(n10567) );
  AND U15853 ( .A(n10569), .B(n10570), .Z(o[5244]) );
  AND U15854 ( .A(p_input[25244]), .B(p_input[15244]), .Z(n10570) );
  AND U15855 ( .A(p_input[5244]), .B(p_input[35244]), .Z(n10569) );
  AND U15856 ( .A(n10571), .B(n10572), .Z(o[5243]) );
  AND U15857 ( .A(p_input[25243]), .B(p_input[15243]), .Z(n10572) );
  AND U15858 ( .A(p_input[5243]), .B(p_input[35243]), .Z(n10571) );
  AND U15859 ( .A(n10573), .B(n10574), .Z(o[5242]) );
  AND U15860 ( .A(p_input[25242]), .B(p_input[15242]), .Z(n10574) );
  AND U15861 ( .A(p_input[5242]), .B(p_input[35242]), .Z(n10573) );
  AND U15862 ( .A(n10575), .B(n10576), .Z(o[5241]) );
  AND U15863 ( .A(p_input[25241]), .B(p_input[15241]), .Z(n10576) );
  AND U15864 ( .A(p_input[5241]), .B(p_input[35241]), .Z(n10575) );
  AND U15865 ( .A(n10577), .B(n10578), .Z(o[5240]) );
  AND U15866 ( .A(p_input[25240]), .B(p_input[15240]), .Z(n10578) );
  AND U15867 ( .A(p_input[5240]), .B(p_input[35240]), .Z(n10577) );
  AND U15868 ( .A(n10579), .B(n10580), .Z(o[523]) );
  AND U15869 ( .A(p_input[20523]), .B(p_input[10523]), .Z(n10580) );
  AND U15870 ( .A(p_input[523]), .B(p_input[30523]), .Z(n10579) );
  AND U15871 ( .A(n10581), .B(n10582), .Z(o[5239]) );
  AND U15872 ( .A(p_input[25239]), .B(p_input[15239]), .Z(n10582) );
  AND U15873 ( .A(p_input[5239]), .B(p_input[35239]), .Z(n10581) );
  AND U15874 ( .A(n10583), .B(n10584), .Z(o[5238]) );
  AND U15875 ( .A(p_input[25238]), .B(p_input[15238]), .Z(n10584) );
  AND U15876 ( .A(p_input[5238]), .B(p_input[35238]), .Z(n10583) );
  AND U15877 ( .A(n10585), .B(n10586), .Z(o[5237]) );
  AND U15878 ( .A(p_input[25237]), .B(p_input[15237]), .Z(n10586) );
  AND U15879 ( .A(p_input[5237]), .B(p_input[35237]), .Z(n10585) );
  AND U15880 ( .A(n10587), .B(n10588), .Z(o[5236]) );
  AND U15881 ( .A(p_input[25236]), .B(p_input[15236]), .Z(n10588) );
  AND U15882 ( .A(p_input[5236]), .B(p_input[35236]), .Z(n10587) );
  AND U15883 ( .A(n10589), .B(n10590), .Z(o[5235]) );
  AND U15884 ( .A(p_input[25235]), .B(p_input[15235]), .Z(n10590) );
  AND U15885 ( .A(p_input[5235]), .B(p_input[35235]), .Z(n10589) );
  AND U15886 ( .A(n10591), .B(n10592), .Z(o[5234]) );
  AND U15887 ( .A(p_input[25234]), .B(p_input[15234]), .Z(n10592) );
  AND U15888 ( .A(p_input[5234]), .B(p_input[35234]), .Z(n10591) );
  AND U15889 ( .A(n10593), .B(n10594), .Z(o[5233]) );
  AND U15890 ( .A(p_input[25233]), .B(p_input[15233]), .Z(n10594) );
  AND U15891 ( .A(p_input[5233]), .B(p_input[35233]), .Z(n10593) );
  AND U15892 ( .A(n10595), .B(n10596), .Z(o[5232]) );
  AND U15893 ( .A(p_input[25232]), .B(p_input[15232]), .Z(n10596) );
  AND U15894 ( .A(p_input[5232]), .B(p_input[35232]), .Z(n10595) );
  AND U15895 ( .A(n10597), .B(n10598), .Z(o[5231]) );
  AND U15896 ( .A(p_input[25231]), .B(p_input[15231]), .Z(n10598) );
  AND U15897 ( .A(p_input[5231]), .B(p_input[35231]), .Z(n10597) );
  AND U15898 ( .A(n10599), .B(n10600), .Z(o[5230]) );
  AND U15899 ( .A(p_input[25230]), .B(p_input[15230]), .Z(n10600) );
  AND U15900 ( .A(p_input[5230]), .B(p_input[35230]), .Z(n10599) );
  AND U15901 ( .A(n10601), .B(n10602), .Z(o[522]) );
  AND U15902 ( .A(p_input[20522]), .B(p_input[10522]), .Z(n10602) );
  AND U15903 ( .A(p_input[522]), .B(p_input[30522]), .Z(n10601) );
  AND U15904 ( .A(n10603), .B(n10604), .Z(o[5229]) );
  AND U15905 ( .A(p_input[25229]), .B(p_input[15229]), .Z(n10604) );
  AND U15906 ( .A(p_input[5229]), .B(p_input[35229]), .Z(n10603) );
  AND U15907 ( .A(n10605), .B(n10606), .Z(o[5228]) );
  AND U15908 ( .A(p_input[25228]), .B(p_input[15228]), .Z(n10606) );
  AND U15909 ( .A(p_input[5228]), .B(p_input[35228]), .Z(n10605) );
  AND U15910 ( .A(n10607), .B(n10608), .Z(o[5227]) );
  AND U15911 ( .A(p_input[25227]), .B(p_input[15227]), .Z(n10608) );
  AND U15912 ( .A(p_input[5227]), .B(p_input[35227]), .Z(n10607) );
  AND U15913 ( .A(n10609), .B(n10610), .Z(o[5226]) );
  AND U15914 ( .A(p_input[25226]), .B(p_input[15226]), .Z(n10610) );
  AND U15915 ( .A(p_input[5226]), .B(p_input[35226]), .Z(n10609) );
  AND U15916 ( .A(n10611), .B(n10612), .Z(o[5225]) );
  AND U15917 ( .A(p_input[25225]), .B(p_input[15225]), .Z(n10612) );
  AND U15918 ( .A(p_input[5225]), .B(p_input[35225]), .Z(n10611) );
  AND U15919 ( .A(n10613), .B(n10614), .Z(o[5224]) );
  AND U15920 ( .A(p_input[25224]), .B(p_input[15224]), .Z(n10614) );
  AND U15921 ( .A(p_input[5224]), .B(p_input[35224]), .Z(n10613) );
  AND U15922 ( .A(n10615), .B(n10616), .Z(o[5223]) );
  AND U15923 ( .A(p_input[25223]), .B(p_input[15223]), .Z(n10616) );
  AND U15924 ( .A(p_input[5223]), .B(p_input[35223]), .Z(n10615) );
  AND U15925 ( .A(n10617), .B(n10618), .Z(o[5222]) );
  AND U15926 ( .A(p_input[25222]), .B(p_input[15222]), .Z(n10618) );
  AND U15927 ( .A(p_input[5222]), .B(p_input[35222]), .Z(n10617) );
  AND U15928 ( .A(n10619), .B(n10620), .Z(o[5221]) );
  AND U15929 ( .A(p_input[25221]), .B(p_input[15221]), .Z(n10620) );
  AND U15930 ( .A(p_input[5221]), .B(p_input[35221]), .Z(n10619) );
  AND U15931 ( .A(n10621), .B(n10622), .Z(o[5220]) );
  AND U15932 ( .A(p_input[25220]), .B(p_input[15220]), .Z(n10622) );
  AND U15933 ( .A(p_input[5220]), .B(p_input[35220]), .Z(n10621) );
  AND U15934 ( .A(n10623), .B(n10624), .Z(o[521]) );
  AND U15935 ( .A(p_input[20521]), .B(p_input[10521]), .Z(n10624) );
  AND U15936 ( .A(p_input[521]), .B(p_input[30521]), .Z(n10623) );
  AND U15937 ( .A(n10625), .B(n10626), .Z(o[5219]) );
  AND U15938 ( .A(p_input[25219]), .B(p_input[15219]), .Z(n10626) );
  AND U15939 ( .A(p_input[5219]), .B(p_input[35219]), .Z(n10625) );
  AND U15940 ( .A(n10627), .B(n10628), .Z(o[5218]) );
  AND U15941 ( .A(p_input[25218]), .B(p_input[15218]), .Z(n10628) );
  AND U15942 ( .A(p_input[5218]), .B(p_input[35218]), .Z(n10627) );
  AND U15943 ( .A(n10629), .B(n10630), .Z(o[5217]) );
  AND U15944 ( .A(p_input[25217]), .B(p_input[15217]), .Z(n10630) );
  AND U15945 ( .A(p_input[5217]), .B(p_input[35217]), .Z(n10629) );
  AND U15946 ( .A(n10631), .B(n10632), .Z(o[5216]) );
  AND U15947 ( .A(p_input[25216]), .B(p_input[15216]), .Z(n10632) );
  AND U15948 ( .A(p_input[5216]), .B(p_input[35216]), .Z(n10631) );
  AND U15949 ( .A(n10633), .B(n10634), .Z(o[5215]) );
  AND U15950 ( .A(p_input[25215]), .B(p_input[15215]), .Z(n10634) );
  AND U15951 ( .A(p_input[5215]), .B(p_input[35215]), .Z(n10633) );
  AND U15952 ( .A(n10635), .B(n10636), .Z(o[5214]) );
  AND U15953 ( .A(p_input[25214]), .B(p_input[15214]), .Z(n10636) );
  AND U15954 ( .A(p_input[5214]), .B(p_input[35214]), .Z(n10635) );
  AND U15955 ( .A(n10637), .B(n10638), .Z(o[5213]) );
  AND U15956 ( .A(p_input[25213]), .B(p_input[15213]), .Z(n10638) );
  AND U15957 ( .A(p_input[5213]), .B(p_input[35213]), .Z(n10637) );
  AND U15958 ( .A(n10639), .B(n10640), .Z(o[5212]) );
  AND U15959 ( .A(p_input[25212]), .B(p_input[15212]), .Z(n10640) );
  AND U15960 ( .A(p_input[5212]), .B(p_input[35212]), .Z(n10639) );
  AND U15961 ( .A(n10641), .B(n10642), .Z(o[5211]) );
  AND U15962 ( .A(p_input[25211]), .B(p_input[15211]), .Z(n10642) );
  AND U15963 ( .A(p_input[5211]), .B(p_input[35211]), .Z(n10641) );
  AND U15964 ( .A(n10643), .B(n10644), .Z(o[5210]) );
  AND U15965 ( .A(p_input[25210]), .B(p_input[15210]), .Z(n10644) );
  AND U15966 ( .A(p_input[5210]), .B(p_input[35210]), .Z(n10643) );
  AND U15967 ( .A(n10645), .B(n10646), .Z(o[520]) );
  AND U15968 ( .A(p_input[20520]), .B(p_input[10520]), .Z(n10646) );
  AND U15969 ( .A(p_input[520]), .B(p_input[30520]), .Z(n10645) );
  AND U15970 ( .A(n10647), .B(n10648), .Z(o[5209]) );
  AND U15971 ( .A(p_input[25209]), .B(p_input[15209]), .Z(n10648) );
  AND U15972 ( .A(p_input[5209]), .B(p_input[35209]), .Z(n10647) );
  AND U15973 ( .A(n10649), .B(n10650), .Z(o[5208]) );
  AND U15974 ( .A(p_input[25208]), .B(p_input[15208]), .Z(n10650) );
  AND U15975 ( .A(p_input[5208]), .B(p_input[35208]), .Z(n10649) );
  AND U15976 ( .A(n10651), .B(n10652), .Z(o[5207]) );
  AND U15977 ( .A(p_input[25207]), .B(p_input[15207]), .Z(n10652) );
  AND U15978 ( .A(p_input[5207]), .B(p_input[35207]), .Z(n10651) );
  AND U15979 ( .A(n10653), .B(n10654), .Z(o[5206]) );
  AND U15980 ( .A(p_input[25206]), .B(p_input[15206]), .Z(n10654) );
  AND U15981 ( .A(p_input[5206]), .B(p_input[35206]), .Z(n10653) );
  AND U15982 ( .A(n10655), .B(n10656), .Z(o[5205]) );
  AND U15983 ( .A(p_input[25205]), .B(p_input[15205]), .Z(n10656) );
  AND U15984 ( .A(p_input[5205]), .B(p_input[35205]), .Z(n10655) );
  AND U15985 ( .A(n10657), .B(n10658), .Z(o[5204]) );
  AND U15986 ( .A(p_input[25204]), .B(p_input[15204]), .Z(n10658) );
  AND U15987 ( .A(p_input[5204]), .B(p_input[35204]), .Z(n10657) );
  AND U15988 ( .A(n10659), .B(n10660), .Z(o[5203]) );
  AND U15989 ( .A(p_input[25203]), .B(p_input[15203]), .Z(n10660) );
  AND U15990 ( .A(p_input[5203]), .B(p_input[35203]), .Z(n10659) );
  AND U15991 ( .A(n10661), .B(n10662), .Z(o[5202]) );
  AND U15992 ( .A(p_input[25202]), .B(p_input[15202]), .Z(n10662) );
  AND U15993 ( .A(p_input[5202]), .B(p_input[35202]), .Z(n10661) );
  AND U15994 ( .A(n10663), .B(n10664), .Z(o[5201]) );
  AND U15995 ( .A(p_input[25201]), .B(p_input[15201]), .Z(n10664) );
  AND U15996 ( .A(p_input[5201]), .B(p_input[35201]), .Z(n10663) );
  AND U15997 ( .A(n10665), .B(n10666), .Z(o[5200]) );
  AND U15998 ( .A(p_input[25200]), .B(p_input[15200]), .Z(n10666) );
  AND U15999 ( .A(p_input[5200]), .B(p_input[35200]), .Z(n10665) );
  AND U16000 ( .A(n10667), .B(n10668), .Z(o[51]) );
  AND U16001 ( .A(p_input[20051]), .B(p_input[10051]), .Z(n10668) );
  AND U16002 ( .A(p_input[51]), .B(p_input[30051]), .Z(n10667) );
  AND U16003 ( .A(n10669), .B(n10670), .Z(o[519]) );
  AND U16004 ( .A(p_input[20519]), .B(p_input[10519]), .Z(n10670) );
  AND U16005 ( .A(p_input[519]), .B(p_input[30519]), .Z(n10669) );
  AND U16006 ( .A(n10671), .B(n10672), .Z(o[5199]) );
  AND U16007 ( .A(p_input[25199]), .B(p_input[15199]), .Z(n10672) );
  AND U16008 ( .A(p_input[5199]), .B(p_input[35199]), .Z(n10671) );
  AND U16009 ( .A(n10673), .B(n10674), .Z(o[5198]) );
  AND U16010 ( .A(p_input[25198]), .B(p_input[15198]), .Z(n10674) );
  AND U16011 ( .A(p_input[5198]), .B(p_input[35198]), .Z(n10673) );
  AND U16012 ( .A(n10675), .B(n10676), .Z(o[5197]) );
  AND U16013 ( .A(p_input[25197]), .B(p_input[15197]), .Z(n10676) );
  AND U16014 ( .A(p_input[5197]), .B(p_input[35197]), .Z(n10675) );
  AND U16015 ( .A(n10677), .B(n10678), .Z(o[5196]) );
  AND U16016 ( .A(p_input[25196]), .B(p_input[15196]), .Z(n10678) );
  AND U16017 ( .A(p_input[5196]), .B(p_input[35196]), .Z(n10677) );
  AND U16018 ( .A(n10679), .B(n10680), .Z(o[5195]) );
  AND U16019 ( .A(p_input[25195]), .B(p_input[15195]), .Z(n10680) );
  AND U16020 ( .A(p_input[5195]), .B(p_input[35195]), .Z(n10679) );
  AND U16021 ( .A(n10681), .B(n10682), .Z(o[5194]) );
  AND U16022 ( .A(p_input[25194]), .B(p_input[15194]), .Z(n10682) );
  AND U16023 ( .A(p_input[5194]), .B(p_input[35194]), .Z(n10681) );
  AND U16024 ( .A(n10683), .B(n10684), .Z(o[5193]) );
  AND U16025 ( .A(p_input[25193]), .B(p_input[15193]), .Z(n10684) );
  AND U16026 ( .A(p_input[5193]), .B(p_input[35193]), .Z(n10683) );
  AND U16027 ( .A(n10685), .B(n10686), .Z(o[5192]) );
  AND U16028 ( .A(p_input[25192]), .B(p_input[15192]), .Z(n10686) );
  AND U16029 ( .A(p_input[5192]), .B(p_input[35192]), .Z(n10685) );
  AND U16030 ( .A(n10687), .B(n10688), .Z(o[5191]) );
  AND U16031 ( .A(p_input[25191]), .B(p_input[15191]), .Z(n10688) );
  AND U16032 ( .A(p_input[5191]), .B(p_input[35191]), .Z(n10687) );
  AND U16033 ( .A(n10689), .B(n10690), .Z(o[5190]) );
  AND U16034 ( .A(p_input[25190]), .B(p_input[15190]), .Z(n10690) );
  AND U16035 ( .A(p_input[5190]), .B(p_input[35190]), .Z(n10689) );
  AND U16036 ( .A(n10691), .B(n10692), .Z(o[518]) );
  AND U16037 ( .A(p_input[20518]), .B(p_input[10518]), .Z(n10692) );
  AND U16038 ( .A(p_input[518]), .B(p_input[30518]), .Z(n10691) );
  AND U16039 ( .A(n10693), .B(n10694), .Z(o[5189]) );
  AND U16040 ( .A(p_input[25189]), .B(p_input[15189]), .Z(n10694) );
  AND U16041 ( .A(p_input[5189]), .B(p_input[35189]), .Z(n10693) );
  AND U16042 ( .A(n10695), .B(n10696), .Z(o[5188]) );
  AND U16043 ( .A(p_input[25188]), .B(p_input[15188]), .Z(n10696) );
  AND U16044 ( .A(p_input[5188]), .B(p_input[35188]), .Z(n10695) );
  AND U16045 ( .A(n10697), .B(n10698), .Z(o[5187]) );
  AND U16046 ( .A(p_input[25187]), .B(p_input[15187]), .Z(n10698) );
  AND U16047 ( .A(p_input[5187]), .B(p_input[35187]), .Z(n10697) );
  AND U16048 ( .A(n10699), .B(n10700), .Z(o[5186]) );
  AND U16049 ( .A(p_input[25186]), .B(p_input[15186]), .Z(n10700) );
  AND U16050 ( .A(p_input[5186]), .B(p_input[35186]), .Z(n10699) );
  AND U16051 ( .A(n10701), .B(n10702), .Z(o[5185]) );
  AND U16052 ( .A(p_input[25185]), .B(p_input[15185]), .Z(n10702) );
  AND U16053 ( .A(p_input[5185]), .B(p_input[35185]), .Z(n10701) );
  AND U16054 ( .A(n10703), .B(n10704), .Z(o[5184]) );
  AND U16055 ( .A(p_input[25184]), .B(p_input[15184]), .Z(n10704) );
  AND U16056 ( .A(p_input[5184]), .B(p_input[35184]), .Z(n10703) );
  AND U16057 ( .A(n10705), .B(n10706), .Z(o[5183]) );
  AND U16058 ( .A(p_input[25183]), .B(p_input[15183]), .Z(n10706) );
  AND U16059 ( .A(p_input[5183]), .B(p_input[35183]), .Z(n10705) );
  AND U16060 ( .A(n10707), .B(n10708), .Z(o[5182]) );
  AND U16061 ( .A(p_input[25182]), .B(p_input[15182]), .Z(n10708) );
  AND U16062 ( .A(p_input[5182]), .B(p_input[35182]), .Z(n10707) );
  AND U16063 ( .A(n10709), .B(n10710), .Z(o[5181]) );
  AND U16064 ( .A(p_input[25181]), .B(p_input[15181]), .Z(n10710) );
  AND U16065 ( .A(p_input[5181]), .B(p_input[35181]), .Z(n10709) );
  AND U16066 ( .A(n10711), .B(n10712), .Z(o[5180]) );
  AND U16067 ( .A(p_input[25180]), .B(p_input[15180]), .Z(n10712) );
  AND U16068 ( .A(p_input[5180]), .B(p_input[35180]), .Z(n10711) );
  AND U16069 ( .A(n10713), .B(n10714), .Z(o[517]) );
  AND U16070 ( .A(p_input[20517]), .B(p_input[10517]), .Z(n10714) );
  AND U16071 ( .A(p_input[517]), .B(p_input[30517]), .Z(n10713) );
  AND U16072 ( .A(n10715), .B(n10716), .Z(o[5179]) );
  AND U16073 ( .A(p_input[25179]), .B(p_input[15179]), .Z(n10716) );
  AND U16074 ( .A(p_input[5179]), .B(p_input[35179]), .Z(n10715) );
  AND U16075 ( .A(n10717), .B(n10718), .Z(o[5178]) );
  AND U16076 ( .A(p_input[25178]), .B(p_input[15178]), .Z(n10718) );
  AND U16077 ( .A(p_input[5178]), .B(p_input[35178]), .Z(n10717) );
  AND U16078 ( .A(n10719), .B(n10720), .Z(o[5177]) );
  AND U16079 ( .A(p_input[25177]), .B(p_input[15177]), .Z(n10720) );
  AND U16080 ( .A(p_input[5177]), .B(p_input[35177]), .Z(n10719) );
  AND U16081 ( .A(n10721), .B(n10722), .Z(o[5176]) );
  AND U16082 ( .A(p_input[25176]), .B(p_input[15176]), .Z(n10722) );
  AND U16083 ( .A(p_input[5176]), .B(p_input[35176]), .Z(n10721) );
  AND U16084 ( .A(n10723), .B(n10724), .Z(o[5175]) );
  AND U16085 ( .A(p_input[25175]), .B(p_input[15175]), .Z(n10724) );
  AND U16086 ( .A(p_input[5175]), .B(p_input[35175]), .Z(n10723) );
  AND U16087 ( .A(n10725), .B(n10726), .Z(o[5174]) );
  AND U16088 ( .A(p_input[25174]), .B(p_input[15174]), .Z(n10726) );
  AND U16089 ( .A(p_input[5174]), .B(p_input[35174]), .Z(n10725) );
  AND U16090 ( .A(n10727), .B(n10728), .Z(o[5173]) );
  AND U16091 ( .A(p_input[25173]), .B(p_input[15173]), .Z(n10728) );
  AND U16092 ( .A(p_input[5173]), .B(p_input[35173]), .Z(n10727) );
  AND U16093 ( .A(n10729), .B(n10730), .Z(o[5172]) );
  AND U16094 ( .A(p_input[25172]), .B(p_input[15172]), .Z(n10730) );
  AND U16095 ( .A(p_input[5172]), .B(p_input[35172]), .Z(n10729) );
  AND U16096 ( .A(n10731), .B(n10732), .Z(o[5171]) );
  AND U16097 ( .A(p_input[25171]), .B(p_input[15171]), .Z(n10732) );
  AND U16098 ( .A(p_input[5171]), .B(p_input[35171]), .Z(n10731) );
  AND U16099 ( .A(n10733), .B(n10734), .Z(o[5170]) );
  AND U16100 ( .A(p_input[25170]), .B(p_input[15170]), .Z(n10734) );
  AND U16101 ( .A(p_input[5170]), .B(p_input[35170]), .Z(n10733) );
  AND U16102 ( .A(n10735), .B(n10736), .Z(o[516]) );
  AND U16103 ( .A(p_input[20516]), .B(p_input[10516]), .Z(n10736) );
  AND U16104 ( .A(p_input[516]), .B(p_input[30516]), .Z(n10735) );
  AND U16105 ( .A(n10737), .B(n10738), .Z(o[5169]) );
  AND U16106 ( .A(p_input[25169]), .B(p_input[15169]), .Z(n10738) );
  AND U16107 ( .A(p_input[5169]), .B(p_input[35169]), .Z(n10737) );
  AND U16108 ( .A(n10739), .B(n10740), .Z(o[5168]) );
  AND U16109 ( .A(p_input[25168]), .B(p_input[15168]), .Z(n10740) );
  AND U16110 ( .A(p_input[5168]), .B(p_input[35168]), .Z(n10739) );
  AND U16111 ( .A(n10741), .B(n10742), .Z(o[5167]) );
  AND U16112 ( .A(p_input[25167]), .B(p_input[15167]), .Z(n10742) );
  AND U16113 ( .A(p_input[5167]), .B(p_input[35167]), .Z(n10741) );
  AND U16114 ( .A(n10743), .B(n10744), .Z(o[5166]) );
  AND U16115 ( .A(p_input[25166]), .B(p_input[15166]), .Z(n10744) );
  AND U16116 ( .A(p_input[5166]), .B(p_input[35166]), .Z(n10743) );
  AND U16117 ( .A(n10745), .B(n10746), .Z(o[5165]) );
  AND U16118 ( .A(p_input[25165]), .B(p_input[15165]), .Z(n10746) );
  AND U16119 ( .A(p_input[5165]), .B(p_input[35165]), .Z(n10745) );
  AND U16120 ( .A(n10747), .B(n10748), .Z(o[5164]) );
  AND U16121 ( .A(p_input[25164]), .B(p_input[15164]), .Z(n10748) );
  AND U16122 ( .A(p_input[5164]), .B(p_input[35164]), .Z(n10747) );
  AND U16123 ( .A(n10749), .B(n10750), .Z(o[5163]) );
  AND U16124 ( .A(p_input[25163]), .B(p_input[15163]), .Z(n10750) );
  AND U16125 ( .A(p_input[5163]), .B(p_input[35163]), .Z(n10749) );
  AND U16126 ( .A(n10751), .B(n10752), .Z(o[5162]) );
  AND U16127 ( .A(p_input[25162]), .B(p_input[15162]), .Z(n10752) );
  AND U16128 ( .A(p_input[5162]), .B(p_input[35162]), .Z(n10751) );
  AND U16129 ( .A(n10753), .B(n10754), .Z(o[5161]) );
  AND U16130 ( .A(p_input[25161]), .B(p_input[15161]), .Z(n10754) );
  AND U16131 ( .A(p_input[5161]), .B(p_input[35161]), .Z(n10753) );
  AND U16132 ( .A(n10755), .B(n10756), .Z(o[5160]) );
  AND U16133 ( .A(p_input[25160]), .B(p_input[15160]), .Z(n10756) );
  AND U16134 ( .A(p_input[5160]), .B(p_input[35160]), .Z(n10755) );
  AND U16135 ( .A(n10757), .B(n10758), .Z(o[515]) );
  AND U16136 ( .A(p_input[20515]), .B(p_input[10515]), .Z(n10758) );
  AND U16137 ( .A(p_input[515]), .B(p_input[30515]), .Z(n10757) );
  AND U16138 ( .A(n10759), .B(n10760), .Z(o[5159]) );
  AND U16139 ( .A(p_input[25159]), .B(p_input[15159]), .Z(n10760) );
  AND U16140 ( .A(p_input[5159]), .B(p_input[35159]), .Z(n10759) );
  AND U16141 ( .A(n10761), .B(n10762), .Z(o[5158]) );
  AND U16142 ( .A(p_input[25158]), .B(p_input[15158]), .Z(n10762) );
  AND U16143 ( .A(p_input[5158]), .B(p_input[35158]), .Z(n10761) );
  AND U16144 ( .A(n10763), .B(n10764), .Z(o[5157]) );
  AND U16145 ( .A(p_input[25157]), .B(p_input[15157]), .Z(n10764) );
  AND U16146 ( .A(p_input[5157]), .B(p_input[35157]), .Z(n10763) );
  AND U16147 ( .A(n10765), .B(n10766), .Z(o[5156]) );
  AND U16148 ( .A(p_input[25156]), .B(p_input[15156]), .Z(n10766) );
  AND U16149 ( .A(p_input[5156]), .B(p_input[35156]), .Z(n10765) );
  AND U16150 ( .A(n10767), .B(n10768), .Z(o[5155]) );
  AND U16151 ( .A(p_input[25155]), .B(p_input[15155]), .Z(n10768) );
  AND U16152 ( .A(p_input[5155]), .B(p_input[35155]), .Z(n10767) );
  AND U16153 ( .A(n10769), .B(n10770), .Z(o[5154]) );
  AND U16154 ( .A(p_input[25154]), .B(p_input[15154]), .Z(n10770) );
  AND U16155 ( .A(p_input[5154]), .B(p_input[35154]), .Z(n10769) );
  AND U16156 ( .A(n10771), .B(n10772), .Z(o[5153]) );
  AND U16157 ( .A(p_input[25153]), .B(p_input[15153]), .Z(n10772) );
  AND U16158 ( .A(p_input[5153]), .B(p_input[35153]), .Z(n10771) );
  AND U16159 ( .A(n10773), .B(n10774), .Z(o[5152]) );
  AND U16160 ( .A(p_input[25152]), .B(p_input[15152]), .Z(n10774) );
  AND U16161 ( .A(p_input[5152]), .B(p_input[35152]), .Z(n10773) );
  AND U16162 ( .A(n10775), .B(n10776), .Z(o[5151]) );
  AND U16163 ( .A(p_input[25151]), .B(p_input[15151]), .Z(n10776) );
  AND U16164 ( .A(p_input[5151]), .B(p_input[35151]), .Z(n10775) );
  AND U16165 ( .A(n10777), .B(n10778), .Z(o[5150]) );
  AND U16166 ( .A(p_input[25150]), .B(p_input[15150]), .Z(n10778) );
  AND U16167 ( .A(p_input[5150]), .B(p_input[35150]), .Z(n10777) );
  AND U16168 ( .A(n10779), .B(n10780), .Z(o[514]) );
  AND U16169 ( .A(p_input[20514]), .B(p_input[10514]), .Z(n10780) );
  AND U16170 ( .A(p_input[514]), .B(p_input[30514]), .Z(n10779) );
  AND U16171 ( .A(n10781), .B(n10782), .Z(o[5149]) );
  AND U16172 ( .A(p_input[25149]), .B(p_input[15149]), .Z(n10782) );
  AND U16173 ( .A(p_input[5149]), .B(p_input[35149]), .Z(n10781) );
  AND U16174 ( .A(n10783), .B(n10784), .Z(o[5148]) );
  AND U16175 ( .A(p_input[25148]), .B(p_input[15148]), .Z(n10784) );
  AND U16176 ( .A(p_input[5148]), .B(p_input[35148]), .Z(n10783) );
  AND U16177 ( .A(n10785), .B(n10786), .Z(o[5147]) );
  AND U16178 ( .A(p_input[25147]), .B(p_input[15147]), .Z(n10786) );
  AND U16179 ( .A(p_input[5147]), .B(p_input[35147]), .Z(n10785) );
  AND U16180 ( .A(n10787), .B(n10788), .Z(o[5146]) );
  AND U16181 ( .A(p_input[25146]), .B(p_input[15146]), .Z(n10788) );
  AND U16182 ( .A(p_input[5146]), .B(p_input[35146]), .Z(n10787) );
  AND U16183 ( .A(n10789), .B(n10790), .Z(o[5145]) );
  AND U16184 ( .A(p_input[25145]), .B(p_input[15145]), .Z(n10790) );
  AND U16185 ( .A(p_input[5145]), .B(p_input[35145]), .Z(n10789) );
  AND U16186 ( .A(n10791), .B(n10792), .Z(o[5144]) );
  AND U16187 ( .A(p_input[25144]), .B(p_input[15144]), .Z(n10792) );
  AND U16188 ( .A(p_input[5144]), .B(p_input[35144]), .Z(n10791) );
  AND U16189 ( .A(n10793), .B(n10794), .Z(o[5143]) );
  AND U16190 ( .A(p_input[25143]), .B(p_input[15143]), .Z(n10794) );
  AND U16191 ( .A(p_input[5143]), .B(p_input[35143]), .Z(n10793) );
  AND U16192 ( .A(n10795), .B(n10796), .Z(o[5142]) );
  AND U16193 ( .A(p_input[25142]), .B(p_input[15142]), .Z(n10796) );
  AND U16194 ( .A(p_input[5142]), .B(p_input[35142]), .Z(n10795) );
  AND U16195 ( .A(n10797), .B(n10798), .Z(o[5141]) );
  AND U16196 ( .A(p_input[25141]), .B(p_input[15141]), .Z(n10798) );
  AND U16197 ( .A(p_input[5141]), .B(p_input[35141]), .Z(n10797) );
  AND U16198 ( .A(n10799), .B(n10800), .Z(o[5140]) );
  AND U16199 ( .A(p_input[25140]), .B(p_input[15140]), .Z(n10800) );
  AND U16200 ( .A(p_input[5140]), .B(p_input[35140]), .Z(n10799) );
  AND U16201 ( .A(n10801), .B(n10802), .Z(o[513]) );
  AND U16202 ( .A(p_input[20513]), .B(p_input[10513]), .Z(n10802) );
  AND U16203 ( .A(p_input[513]), .B(p_input[30513]), .Z(n10801) );
  AND U16204 ( .A(n10803), .B(n10804), .Z(o[5139]) );
  AND U16205 ( .A(p_input[25139]), .B(p_input[15139]), .Z(n10804) );
  AND U16206 ( .A(p_input[5139]), .B(p_input[35139]), .Z(n10803) );
  AND U16207 ( .A(n10805), .B(n10806), .Z(o[5138]) );
  AND U16208 ( .A(p_input[25138]), .B(p_input[15138]), .Z(n10806) );
  AND U16209 ( .A(p_input[5138]), .B(p_input[35138]), .Z(n10805) );
  AND U16210 ( .A(n10807), .B(n10808), .Z(o[5137]) );
  AND U16211 ( .A(p_input[25137]), .B(p_input[15137]), .Z(n10808) );
  AND U16212 ( .A(p_input[5137]), .B(p_input[35137]), .Z(n10807) );
  AND U16213 ( .A(n10809), .B(n10810), .Z(o[5136]) );
  AND U16214 ( .A(p_input[25136]), .B(p_input[15136]), .Z(n10810) );
  AND U16215 ( .A(p_input[5136]), .B(p_input[35136]), .Z(n10809) );
  AND U16216 ( .A(n10811), .B(n10812), .Z(o[5135]) );
  AND U16217 ( .A(p_input[25135]), .B(p_input[15135]), .Z(n10812) );
  AND U16218 ( .A(p_input[5135]), .B(p_input[35135]), .Z(n10811) );
  AND U16219 ( .A(n10813), .B(n10814), .Z(o[5134]) );
  AND U16220 ( .A(p_input[25134]), .B(p_input[15134]), .Z(n10814) );
  AND U16221 ( .A(p_input[5134]), .B(p_input[35134]), .Z(n10813) );
  AND U16222 ( .A(n10815), .B(n10816), .Z(o[5133]) );
  AND U16223 ( .A(p_input[25133]), .B(p_input[15133]), .Z(n10816) );
  AND U16224 ( .A(p_input[5133]), .B(p_input[35133]), .Z(n10815) );
  AND U16225 ( .A(n10817), .B(n10818), .Z(o[5132]) );
  AND U16226 ( .A(p_input[25132]), .B(p_input[15132]), .Z(n10818) );
  AND U16227 ( .A(p_input[5132]), .B(p_input[35132]), .Z(n10817) );
  AND U16228 ( .A(n10819), .B(n10820), .Z(o[5131]) );
  AND U16229 ( .A(p_input[25131]), .B(p_input[15131]), .Z(n10820) );
  AND U16230 ( .A(p_input[5131]), .B(p_input[35131]), .Z(n10819) );
  AND U16231 ( .A(n10821), .B(n10822), .Z(o[5130]) );
  AND U16232 ( .A(p_input[25130]), .B(p_input[15130]), .Z(n10822) );
  AND U16233 ( .A(p_input[5130]), .B(p_input[35130]), .Z(n10821) );
  AND U16234 ( .A(n10823), .B(n10824), .Z(o[512]) );
  AND U16235 ( .A(p_input[20512]), .B(p_input[10512]), .Z(n10824) );
  AND U16236 ( .A(p_input[512]), .B(p_input[30512]), .Z(n10823) );
  AND U16237 ( .A(n10825), .B(n10826), .Z(o[5129]) );
  AND U16238 ( .A(p_input[25129]), .B(p_input[15129]), .Z(n10826) );
  AND U16239 ( .A(p_input[5129]), .B(p_input[35129]), .Z(n10825) );
  AND U16240 ( .A(n10827), .B(n10828), .Z(o[5128]) );
  AND U16241 ( .A(p_input[25128]), .B(p_input[15128]), .Z(n10828) );
  AND U16242 ( .A(p_input[5128]), .B(p_input[35128]), .Z(n10827) );
  AND U16243 ( .A(n10829), .B(n10830), .Z(o[5127]) );
  AND U16244 ( .A(p_input[25127]), .B(p_input[15127]), .Z(n10830) );
  AND U16245 ( .A(p_input[5127]), .B(p_input[35127]), .Z(n10829) );
  AND U16246 ( .A(n10831), .B(n10832), .Z(o[5126]) );
  AND U16247 ( .A(p_input[25126]), .B(p_input[15126]), .Z(n10832) );
  AND U16248 ( .A(p_input[5126]), .B(p_input[35126]), .Z(n10831) );
  AND U16249 ( .A(n10833), .B(n10834), .Z(o[5125]) );
  AND U16250 ( .A(p_input[25125]), .B(p_input[15125]), .Z(n10834) );
  AND U16251 ( .A(p_input[5125]), .B(p_input[35125]), .Z(n10833) );
  AND U16252 ( .A(n10835), .B(n10836), .Z(o[5124]) );
  AND U16253 ( .A(p_input[25124]), .B(p_input[15124]), .Z(n10836) );
  AND U16254 ( .A(p_input[5124]), .B(p_input[35124]), .Z(n10835) );
  AND U16255 ( .A(n10837), .B(n10838), .Z(o[5123]) );
  AND U16256 ( .A(p_input[25123]), .B(p_input[15123]), .Z(n10838) );
  AND U16257 ( .A(p_input[5123]), .B(p_input[35123]), .Z(n10837) );
  AND U16258 ( .A(n10839), .B(n10840), .Z(o[5122]) );
  AND U16259 ( .A(p_input[25122]), .B(p_input[15122]), .Z(n10840) );
  AND U16260 ( .A(p_input[5122]), .B(p_input[35122]), .Z(n10839) );
  AND U16261 ( .A(n10841), .B(n10842), .Z(o[5121]) );
  AND U16262 ( .A(p_input[25121]), .B(p_input[15121]), .Z(n10842) );
  AND U16263 ( .A(p_input[5121]), .B(p_input[35121]), .Z(n10841) );
  AND U16264 ( .A(n10843), .B(n10844), .Z(o[5120]) );
  AND U16265 ( .A(p_input[25120]), .B(p_input[15120]), .Z(n10844) );
  AND U16266 ( .A(p_input[5120]), .B(p_input[35120]), .Z(n10843) );
  AND U16267 ( .A(n10845), .B(n10846), .Z(o[511]) );
  AND U16268 ( .A(p_input[20511]), .B(p_input[10511]), .Z(n10846) );
  AND U16269 ( .A(p_input[511]), .B(p_input[30511]), .Z(n10845) );
  AND U16270 ( .A(n10847), .B(n10848), .Z(o[5119]) );
  AND U16271 ( .A(p_input[25119]), .B(p_input[15119]), .Z(n10848) );
  AND U16272 ( .A(p_input[5119]), .B(p_input[35119]), .Z(n10847) );
  AND U16273 ( .A(n10849), .B(n10850), .Z(o[5118]) );
  AND U16274 ( .A(p_input[25118]), .B(p_input[15118]), .Z(n10850) );
  AND U16275 ( .A(p_input[5118]), .B(p_input[35118]), .Z(n10849) );
  AND U16276 ( .A(n10851), .B(n10852), .Z(o[5117]) );
  AND U16277 ( .A(p_input[25117]), .B(p_input[15117]), .Z(n10852) );
  AND U16278 ( .A(p_input[5117]), .B(p_input[35117]), .Z(n10851) );
  AND U16279 ( .A(n10853), .B(n10854), .Z(o[5116]) );
  AND U16280 ( .A(p_input[25116]), .B(p_input[15116]), .Z(n10854) );
  AND U16281 ( .A(p_input[5116]), .B(p_input[35116]), .Z(n10853) );
  AND U16282 ( .A(n10855), .B(n10856), .Z(o[5115]) );
  AND U16283 ( .A(p_input[25115]), .B(p_input[15115]), .Z(n10856) );
  AND U16284 ( .A(p_input[5115]), .B(p_input[35115]), .Z(n10855) );
  AND U16285 ( .A(n10857), .B(n10858), .Z(o[5114]) );
  AND U16286 ( .A(p_input[25114]), .B(p_input[15114]), .Z(n10858) );
  AND U16287 ( .A(p_input[5114]), .B(p_input[35114]), .Z(n10857) );
  AND U16288 ( .A(n10859), .B(n10860), .Z(o[5113]) );
  AND U16289 ( .A(p_input[25113]), .B(p_input[15113]), .Z(n10860) );
  AND U16290 ( .A(p_input[5113]), .B(p_input[35113]), .Z(n10859) );
  AND U16291 ( .A(n10861), .B(n10862), .Z(o[5112]) );
  AND U16292 ( .A(p_input[25112]), .B(p_input[15112]), .Z(n10862) );
  AND U16293 ( .A(p_input[5112]), .B(p_input[35112]), .Z(n10861) );
  AND U16294 ( .A(n10863), .B(n10864), .Z(o[5111]) );
  AND U16295 ( .A(p_input[25111]), .B(p_input[15111]), .Z(n10864) );
  AND U16296 ( .A(p_input[5111]), .B(p_input[35111]), .Z(n10863) );
  AND U16297 ( .A(n10865), .B(n10866), .Z(o[5110]) );
  AND U16298 ( .A(p_input[25110]), .B(p_input[15110]), .Z(n10866) );
  AND U16299 ( .A(p_input[5110]), .B(p_input[35110]), .Z(n10865) );
  AND U16300 ( .A(n10867), .B(n10868), .Z(o[510]) );
  AND U16301 ( .A(p_input[20510]), .B(p_input[10510]), .Z(n10868) );
  AND U16302 ( .A(p_input[510]), .B(p_input[30510]), .Z(n10867) );
  AND U16303 ( .A(n10869), .B(n10870), .Z(o[5109]) );
  AND U16304 ( .A(p_input[25109]), .B(p_input[15109]), .Z(n10870) );
  AND U16305 ( .A(p_input[5109]), .B(p_input[35109]), .Z(n10869) );
  AND U16306 ( .A(n10871), .B(n10872), .Z(o[5108]) );
  AND U16307 ( .A(p_input[25108]), .B(p_input[15108]), .Z(n10872) );
  AND U16308 ( .A(p_input[5108]), .B(p_input[35108]), .Z(n10871) );
  AND U16309 ( .A(n10873), .B(n10874), .Z(o[5107]) );
  AND U16310 ( .A(p_input[25107]), .B(p_input[15107]), .Z(n10874) );
  AND U16311 ( .A(p_input[5107]), .B(p_input[35107]), .Z(n10873) );
  AND U16312 ( .A(n10875), .B(n10876), .Z(o[5106]) );
  AND U16313 ( .A(p_input[25106]), .B(p_input[15106]), .Z(n10876) );
  AND U16314 ( .A(p_input[5106]), .B(p_input[35106]), .Z(n10875) );
  AND U16315 ( .A(n10877), .B(n10878), .Z(o[5105]) );
  AND U16316 ( .A(p_input[25105]), .B(p_input[15105]), .Z(n10878) );
  AND U16317 ( .A(p_input[5105]), .B(p_input[35105]), .Z(n10877) );
  AND U16318 ( .A(n10879), .B(n10880), .Z(o[5104]) );
  AND U16319 ( .A(p_input[25104]), .B(p_input[15104]), .Z(n10880) );
  AND U16320 ( .A(p_input[5104]), .B(p_input[35104]), .Z(n10879) );
  AND U16321 ( .A(n10881), .B(n10882), .Z(o[5103]) );
  AND U16322 ( .A(p_input[25103]), .B(p_input[15103]), .Z(n10882) );
  AND U16323 ( .A(p_input[5103]), .B(p_input[35103]), .Z(n10881) );
  AND U16324 ( .A(n10883), .B(n10884), .Z(o[5102]) );
  AND U16325 ( .A(p_input[25102]), .B(p_input[15102]), .Z(n10884) );
  AND U16326 ( .A(p_input[5102]), .B(p_input[35102]), .Z(n10883) );
  AND U16327 ( .A(n10885), .B(n10886), .Z(o[5101]) );
  AND U16328 ( .A(p_input[25101]), .B(p_input[15101]), .Z(n10886) );
  AND U16329 ( .A(p_input[5101]), .B(p_input[35101]), .Z(n10885) );
  AND U16330 ( .A(n10887), .B(n10888), .Z(o[5100]) );
  AND U16331 ( .A(p_input[25100]), .B(p_input[15100]), .Z(n10888) );
  AND U16332 ( .A(p_input[5100]), .B(p_input[35100]), .Z(n10887) );
  AND U16333 ( .A(n10889), .B(n10890), .Z(o[50]) );
  AND U16334 ( .A(p_input[20050]), .B(p_input[10050]), .Z(n10890) );
  AND U16335 ( .A(p_input[50]), .B(p_input[30050]), .Z(n10889) );
  AND U16336 ( .A(n10891), .B(n10892), .Z(o[509]) );
  AND U16337 ( .A(p_input[20509]), .B(p_input[10509]), .Z(n10892) );
  AND U16338 ( .A(p_input[509]), .B(p_input[30509]), .Z(n10891) );
  AND U16339 ( .A(n10893), .B(n10894), .Z(o[5099]) );
  AND U16340 ( .A(p_input[25099]), .B(p_input[15099]), .Z(n10894) );
  AND U16341 ( .A(p_input[5099]), .B(p_input[35099]), .Z(n10893) );
  AND U16342 ( .A(n10895), .B(n10896), .Z(o[5098]) );
  AND U16343 ( .A(p_input[25098]), .B(p_input[15098]), .Z(n10896) );
  AND U16344 ( .A(p_input[5098]), .B(p_input[35098]), .Z(n10895) );
  AND U16345 ( .A(n10897), .B(n10898), .Z(o[5097]) );
  AND U16346 ( .A(p_input[25097]), .B(p_input[15097]), .Z(n10898) );
  AND U16347 ( .A(p_input[5097]), .B(p_input[35097]), .Z(n10897) );
  AND U16348 ( .A(n10899), .B(n10900), .Z(o[5096]) );
  AND U16349 ( .A(p_input[25096]), .B(p_input[15096]), .Z(n10900) );
  AND U16350 ( .A(p_input[5096]), .B(p_input[35096]), .Z(n10899) );
  AND U16351 ( .A(n10901), .B(n10902), .Z(o[5095]) );
  AND U16352 ( .A(p_input[25095]), .B(p_input[15095]), .Z(n10902) );
  AND U16353 ( .A(p_input[5095]), .B(p_input[35095]), .Z(n10901) );
  AND U16354 ( .A(n10903), .B(n10904), .Z(o[5094]) );
  AND U16355 ( .A(p_input[25094]), .B(p_input[15094]), .Z(n10904) );
  AND U16356 ( .A(p_input[5094]), .B(p_input[35094]), .Z(n10903) );
  AND U16357 ( .A(n10905), .B(n10906), .Z(o[5093]) );
  AND U16358 ( .A(p_input[25093]), .B(p_input[15093]), .Z(n10906) );
  AND U16359 ( .A(p_input[5093]), .B(p_input[35093]), .Z(n10905) );
  AND U16360 ( .A(n10907), .B(n10908), .Z(o[5092]) );
  AND U16361 ( .A(p_input[25092]), .B(p_input[15092]), .Z(n10908) );
  AND U16362 ( .A(p_input[5092]), .B(p_input[35092]), .Z(n10907) );
  AND U16363 ( .A(n10909), .B(n10910), .Z(o[5091]) );
  AND U16364 ( .A(p_input[25091]), .B(p_input[15091]), .Z(n10910) );
  AND U16365 ( .A(p_input[5091]), .B(p_input[35091]), .Z(n10909) );
  AND U16366 ( .A(n10911), .B(n10912), .Z(o[5090]) );
  AND U16367 ( .A(p_input[25090]), .B(p_input[15090]), .Z(n10912) );
  AND U16368 ( .A(p_input[5090]), .B(p_input[35090]), .Z(n10911) );
  AND U16369 ( .A(n10913), .B(n10914), .Z(o[508]) );
  AND U16370 ( .A(p_input[20508]), .B(p_input[10508]), .Z(n10914) );
  AND U16371 ( .A(p_input[508]), .B(p_input[30508]), .Z(n10913) );
  AND U16372 ( .A(n10915), .B(n10916), .Z(o[5089]) );
  AND U16373 ( .A(p_input[25089]), .B(p_input[15089]), .Z(n10916) );
  AND U16374 ( .A(p_input[5089]), .B(p_input[35089]), .Z(n10915) );
  AND U16375 ( .A(n10917), .B(n10918), .Z(o[5088]) );
  AND U16376 ( .A(p_input[25088]), .B(p_input[15088]), .Z(n10918) );
  AND U16377 ( .A(p_input[5088]), .B(p_input[35088]), .Z(n10917) );
  AND U16378 ( .A(n10919), .B(n10920), .Z(o[5087]) );
  AND U16379 ( .A(p_input[25087]), .B(p_input[15087]), .Z(n10920) );
  AND U16380 ( .A(p_input[5087]), .B(p_input[35087]), .Z(n10919) );
  AND U16381 ( .A(n10921), .B(n10922), .Z(o[5086]) );
  AND U16382 ( .A(p_input[25086]), .B(p_input[15086]), .Z(n10922) );
  AND U16383 ( .A(p_input[5086]), .B(p_input[35086]), .Z(n10921) );
  AND U16384 ( .A(n10923), .B(n10924), .Z(o[5085]) );
  AND U16385 ( .A(p_input[25085]), .B(p_input[15085]), .Z(n10924) );
  AND U16386 ( .A(p_input[5085]), .B(p_input[35085]), .Z(n10923) );
  AND U16387 ( .A(n10925), .B(n10926), .Z(o[5084]) );
  AND U16388 ( .A(p_input[25084]), .B(p_input[15084]), .Z(n10926) );
  AND U16389 ( .A(p_input[5084]), .B(p_input[35084]), .Z(n10925) );
  AND U16390 ( .A(n10927), .B(n10928), .Z(o[5083]) );
  AND U16391 ( .A(p_input[25083]), .B(p_input[15083]), .Z(n10928) );
  AND U16392 ( .A(p_input[5083]), .B(p_input[35083]), .Z(n10927) );
  AND U16393 ( .A(n10929), .B(n10930), .Z(o[5082]) );
  AND U16394 ( .A(p_input[25082]), .B(p_input[15082]), .Z(n10930) );
  AND U16395 ( .A(p_input[5082]), .B(p_input[35082]), .Z(n10929) );
  AND U16396 ( .A(n10931), .B(n10932), .Z(o[5081]) );
  AND U16397 ( .A(p_input[25081]), .B(p_input[15081]), .Z(n10932) );
  AND U16398 ( .A(p_input[5081]), .B(p_input[35081]), .Z(n10931) );
  AND U16399 ( .A(n10933), .B(n10934), .Z(o[5080]) );
  AND U16400 ( .A(p_input[25080]), .B(p_input[15080]), .Z(n10934) );
  AND U16401 ( .A(p_input[5080]), .B(p_input[35080]), .Z(n10933) );
  AND U16402 ( .A(n10935), .B(n10936), .Z(o[507]) );
  AND U16403 ( .A(p_input[20507]), .B(p_input[10507]), .Z(n10936) );
  AND U16404 ( .A(p_input[507]), .B(p_input[30507]), .Z(n10935) );
  AND U16405 ( .A(n10937), .B(n10938), .Z(o[5079]) );
  AND U16406 ( .A(p_input[25079]), .B(p_input[15079]), .Z(n10938) );
  AND U16407 ( .A(p_input[5079]), .B(p_input[35079]), .Z(n10937) );
  AND U16408 ( .A(n10939), .B(n10940), .Z(o[5078]) );
  AND U16409 ( .A(p_input[25078]), .B(p_input[15078]), .Z(n10940) );
  AND U16410 ( .A(p_input[5078]), .B(p_input[35078]), .Z(n10939) );
  AND U16411 ( .A(n10941), .B(n10942), .Z(o[5077]) );
  AND U16412 ( .A(p_input[25077]), .B(p_input[15077]), .Z(n10942) );
  AND U16413 ( .A(p_input[5077]), .B(p_input[35077]), .Z(n10941) );
  AND U16414 ( .A(n10943), .B(n10944), .Z(o[5076]) );
  AND U16415 ( .A(p_input[25076]), .B(p_input[15076]), .Z(n10944) );
  AND U16416 ( .A(p_input[5076]), .B(p_input[35076]), .Z(n10943) );
  AND U16417 ( .A(n10945), .B(n10946), .Z(o[5075]) );
  AND U16418 ( .A(p_input[25075]), .B(p_input[15075]), .Z(n10946) );
  AND U16419 ( .A(p_input[5075]), .B(p_input[35075]), .Z(n10945) );
  AND U16420 ( .A(n10947), .B(n10948), .Z(o[5074]) );
  AND U16421 ( .A(p_input[25074]), .B(p_input[15074]), .Z(n10948) );
  AND U16422 ( .A(p_input[5074]), .B(p_input[35074]), .Z(n10947) );
  AND U16423 ( .A(n10949), .B(n10950), .Z(o[5073]) );
  AND U16424 ( .A(p_input[25073]), .B(p_input[15073]), .Z(n10950) );
  AND U16425 ( .A(p_input[5073]), .B(p_input[35073]), .Z(n10949) );
  AND U16426 ( .A(n10951), .B(n10952), .Z(o[5072]) );
  AND U16427 ( .A(p_input[25072]), .B(p_input[15072]), .Z(n10952) );
  AND U16428 ( .A(p_input[5072]), .B(p_input[35072]), .Z(n10951) );
  AND U16429 ( .A(n10953), .B(n10954), .Z(o[5071]) );
  AND U16430 ( .A(p_input[25071]), .B(p_input[15071]), .Z(n10954) );
  AND U16431 ( .A(p_input[5071]), .B(p_input[35071]), .Z(n10953) );
  AND U16432 ( .A(n10955), .B(n10956), .Z(o[5070]) );
  AND U16433 ( .A(p_input[25070]), .B(p_input[15070]), .Z(n10956) );
  AND U16434 ( .A(p_input[5070]), .B(p_input[35070]), .Z(n10955) );
  AND U16435 ( .A(n10957), .B(n10958), .Z(o[506]) );
  AND U16436 ( .A(p_input[20506]), .B(p_input[10506]), .Z(n10958) );
  AND U16437 ( .A(p_input[506]), .B(p_input[30506]), .Z(n10957) );
  AND U16438 ( .A(n10959), .B(n10960), .Z(o[5069]) );
  AND U16439 ( .A(p_input[25069]), .B(p_input[15069]), .Z(n10960) );
  AND U16440 ( .A(p_input[5069]), .B(p_input[35069]), .Z(n10959) );
  AND U16441 ( .A(n10961), .B(n10962), .Z(o[5068]) );
  AND U16442 ( .A(p_input[25068]), .B(p_input[15068]), .Z(n10962) );
  AND U16443 ( .A(p_input[5068]), .B(p_input[35068]), .Z(n10961) );
  AND U16444 ( .A(n10963), .B(n10964), .Z(o[5067]) );
  AND U16445 ( .A(p_input[25067]), .B(p_input[15067]), .Z(n10964) );
  AND U16446 ( .A(p_input[5067]), .B(p_input[35067]), .Z(n10963) );
  AND U16447 ( .A(n10965), .B(n10966), .Z(o[5066]) );
  AND U16448 ( .A(p_input[25066]), .B(p_input[15066]), .Z(n10966) );
  AND U16449 ( .A(p_input[5066]), .B(p_input[35066]), .Z(n10965) );
  AND U16450 ( .A(n10967), .B(n10968), .Z(o[5065]) );
  AND U16451 ( .A(p_input[25065]), .B(p_input[15065]), .Z(n10968) );
  AND U16452 ( .A(p_input[5065]), .B(p_input[35065]), .Z(n10967) );
  AND U16453 ( .A(n10969), .B(n10970), .Z(o[5064]) );
  AND U16454 ( .A(p_input[25064]), .B(p_input[15064]), .Z(n10970) );
  AND U16455 ( .A(p_input[5064]), .B(p_input[35064]), .Z(n10969) );
  AND U16456 ( .A(n10971), .B(n10972), .Z(o[5063]) );
  AND U16457 ( .A(p_input[25063]), .B(p_input[15063]), .Z(n10972) );
  AND U16458 ( .A(p_input[5063]), .B(p_input[35063]), .Z(n10971) );
  AND U16459 ( .A(n10973), .B(n10974), .Z(o[5062]) );
  AND U16460 ( .A(p_input[25062]), .B(p_input[15062]), .Z(n10974) );
  AND U16461 ( .A(p_input[5062]), .B(p_input[35062]), .Z(n10973) );
  AND U16462 ( .A(n10975), .B(n10976), .Z(o[5061]) );
  AND U16463 ( .A(p_input[25061]), .B(p_input[15061]), .Z(n10976) );
  AND U16464 ( .A(p_input[5061]), .B(p_input[35061]), .Z(n10975) );
  AND U16465 ( .A(n10977), .B(n10978), .Z(o[5060]) );
  AND U16466 ( .A(p_input[25060]), .B(p_input[15060]), .Z(n10978) );
  AND U16467 ( .A(p_input[5060]), .B(p_input[35060]), .Z(n10977) );
  AND U16468 ( .A(n10979), .B(n10980), .Z(o[505]) );
  AND U16469 ( .A(p_input[20505]), .B(p_input[10505]), .Z(n10980) );
  AND U16470 ( .A(p_input[505]), .B(p_input[30505]), .Z(n10979) );
  AND U16471 ( .A(n10981), .B(n10982), .Z(o[5059]) );
  AND U16472 ( .A(p_input[25059]), .B(p_input[15059]), .Z(n10982) );
  AND U16473 ( .A(p_input[5059]), .B(p_input[35059]), .Z(n10981) );
  AND U16474 ( .A(n10983), .B(n10984), .Z(o[5058]) );
  AND U16475 ( .A(p_input[25058]), .B(p_input[15058]), .Z(n10984) );
  AND U16476 ( .A(p_input[5058]), .B(p_input[35058]), .Z(n10983) );
  AND U16477 ( .A(n10985), .B(n10986), .Z(o[5057]) );
  AND U16478 ( .A(p_input[25057]), .B(p_input[15057]), .Z(n10986) );
  AND U16479 ( .A(p_input[5057]), .B(p_input[35057]), .Z(n10985) );
  AND U16480 ( .A(n10987), .B(n10988), .Z(o[5056]) );
  AND U16481 ( .A(p_input[25056]), .B(p_input[15056]), .Z(n10988) );
  AND U16482 ( .A(p_input[5056]), .B(p_input[35056]), .Z(n10987) );
  AND U16483 ( .A(n10989), .B(n10990), .Z(o[5055]) );
  AND U16484 ( .A(p_input[25055]), .B(p_input[15055]), .Z(n10990) );
  AND U16485 ( .A(p_input[5055]), .B(p_input[35055]), .Z(n10989) );
  AND U16486 ( .A(n10991), .B(n10992), .Z(o[5054]) );
  AND U16487 ( .A(p_input[25054]), .B(p_input[15054]), .Z(n10992) );
  AND U16488 ( .A(p_input[5054]), .B(p_input[35054]), .Z(n10991) );
  AND U16489 ( .A(n10993), .B(n10994), .Z(o[5053]) );
  AND U16490 ( .A(p_input[25053]), .B(p_input[15053]), .Z(n10994) );
  AND U16491 ( .A(p_input[5053]), .B(p_input[35053]), .Z(n10993) );
  AND U16492 ( .A(n10995), .B(n10996), .Z(o[5052]) );
  AND U16493 ( .A(p_input[25052]), .B(p_input[15052]), .Z(n10996) );
  AND U16494 ( .A(p_input[5052]), .B(p_input[35052]), .Z(n10995) );
  AND U16495 ( .A(n10997), .B(n10998), .Z(o[5051]) );
  AND U16496 ( .A(p_input[25051]), .B(p_input[15051]), .Z(n10998) );
  AND U16497 ( .A(p_input[5051]), .B(p_input[35051]), .Z(n10997) );
  AND U16498 ( .A(n10999), .B(n11000), .Z(o[5050]) );
  AND U16499 ( .A(p_input[25050]), .B(p_input[15050]), .Z(n11000) );
  AND U16500 ( .A(p_input[5050]), .B(p_input[35050]), .Z(n10999) );
  AND U16501 ( .A(n11001), .B(n11002), .Z(o[504]) );
  AND U16502 ( .A(p_input[20504]), .B(p_input[10504]), .Z(n11002) );
  AND U16503 ( .A(p_input[504]), .B(p_input[30504]), .Z(n11001) );
  AND U16504 ( .A(n11003), .B(n11004), .Z(o[5049]) );
  AND U16505 ( .A(p_input[25049]), .B(p_input[15049]), .Z(n11004) );
  AND U16506 ( .A(p_input[5049]), .B(p_input[35049]), .Z(n11003) );
  AND U16507 ( .A(n11005), .B(n11006), .Z(o[5048]) );
  AND U16508 ( .A(p_input[25048]), .B(p_input[15048]), .Z(n11006) );
  AND U16509 ( .A(p_input[5048]), .B(p_input[35048]), .Z(n11005) );
  AND U16510 ( .A(n11007), .B(n11008), .Z(o[5047]) );
  AND U16511 ( .A(p_input[25047]), .B(p_input[15047]), .Z(n11008) );
  AND U16512 ( .A(p_input[5047]), .B(p_input[35047]), .Z(n11007) );
  AND U16513 ( .A(n11009), .B(n11010), .Z(o[5046]) );
  AND U16514 ( .A(p_input[25046]), .B(p_input[15046]), .Z(n11010) );
  AND U16515 ( .A(p_input[5046]), .B(p_input[35046]), .Z(n11009) );
  AND U16516 ( .A(n11011), .B(n11012), .Z(o[5045]) );
  AND U16517 ( .A(p_input[25045]), .B(p_input[15045]), .Z(n11012) );
  AND U16518 ( .A(p_input[5045]), .B(p_input[35045]), .Z(n11011) );
  AND U16519 ( .A(n11013), .B(n11014), .Z(o[5044]) );
  AND U16520 ( .A(p_input[25044]), .B(p_input[15044]), .Z(n11014) );
  AND U16521 ( .A(p_input[5044]), .B(p_input[35044]), .Z(n11013) );
  AND U16522 ( .A(n11015), .B(n11016), .Z(o[5043]) );
  AND U16523 ( .A(p_input[25043]), .B(p_input[15043]), .Z(n11016) );
  AND U16524 ( .A(p_input[5043]), .B(p_input[35043]), .Z(n11015) );
  AND U16525 ( .A(n11017), .B(n11018), .Z(o[5042]) );
  AND U16526 ( .A(p_input[25042]), .B(p_input[15042]), .Z(n11018) );
  AND U16527 ( .A(p_input[5042]), .B(p_input[35042]), .Z(n11017) );
  AND U16528 ( .A(n11019), .B(n11020), .Z(o[5041]) );
  AND U16529 ( .A(p_input[25041]), .B(p_input[15041]), .Z(n11020) );
  AND U16530 ( .A(p_input[5041]), .B(p_input[35041]), .Z(n11019) );
  AND U16531 ( .A(n11021), .B(n11022), .Z(o[5040]) );
  AND U16532 ( .A(p_input[25040]), .B(p_input[15040]), .Z(n11022) );
  AND U16533 ( .A(p_input[5040]), .B(p_input[35040]), .Z(n11021) );
  AND U16534 ( .A(n11023), .B(n11024), .Z(o[503]) );
  AND U16535 ( .A(p_input[20503]), .B(p_input[10503]), .Z(n11024) );
  AND U16536 ( .A(p_input[503]), .B(p_input[30503]), .Z(n11023) );
  AND U16537 ( .A(n11025), .B(n11026), .Z(o[5039]) );
  AND U16538 ( .A(p_input[25039]), .B(p_input[15039]), .Z(n11026) );
  AND U16539 ( .A(p_input[5039]), .B(p_input[35039]), .Z(n11025) );
  AND U16540 ( .A(n11027), .B(n11028), .Z(o[5038]) );
  AND U16541 ( .A(p_input[25038]), .B(p_input[15038]), .Z(n11028) );
  AND U16542 ( .A(p_input[5038]), .B(p_input[35038]), .Z(n11027) );
  AND U16543 ( .A(n11029), .B(n11030), .Z(o[5037]) );
  AND U16544 ( .A(p_input[25037]), .B(p_input[15037]), .Z(n11030) );
  AND U16545 ( .A(p_input[5037]), .B(p_input[35037]), .Z(n11029) );
  AND U16546 ( .A(n11031), .B(n11032), .Z(o[5036]) );
  AND U16547 ( .A(p_input[25036]), .B(p_input[15036]), .Z(n11032) );
  AND U16548 ( .A(p_input[5036]), .B(p_input[35036]), .Z(n11031) );
  AND U16549 ( .A(n11033), .B(n11034), .Z(o[5035]) );
  AND U16550 ( .A(p_input[25035]), .B(p_input[15035]), .Z(n11034) );
  AND U16551 ( .A(p_input[5035]), .B(p_input[35035]), .Z(n11033) );
  AND U16552 ( .A(n11035), .B(n11036), .Z(o[5034]) );
  AND U16553 ( .A(p_input[25034]), .B(p_input[15034]), .Z(n11036) );
  AND U16554 ( .A(p_input[5034]), .B(p_input[35034]), .Z(n11035) );
  AND U16555 ( .A(n11037), .B(n11038), .Z(o[5033]) );
  AND U16556 ( .A(p_input[25033]), .B(p_input[15033]), .Z(n11038) );
  AND U16557 ( .A(p_input[5033]), .B(p_input[35033]), .Z(n11037) );
  AND U16558 ( .A(n11039), .B(n11040), .Z(o[5032]) );
  AND U16559 ( .A(p_input[25032]), .B(p_input[15032]), .Z(n11040) );
  AND U16560 ( .A(p_input[5032]), .B(p_input[35032]), .Z(n11039) );
  AND U16561 ( .A(n11041), .B(n11042), .Z(o[5031]) );
  AND U16562 ( .A(p_input[25031]), .B(p_input[15031]), .Z(n11042) );
  AND U16563 ( .A(p_input[5031]), .B(p_input[35031]), .Z(n11041) );
  AND U16564 ( .A(n11043), .B(n11044), .Z(o[5030]) );
  AND U16565 ( .A(p_input[25030]), .B(p_input[15030]), .Z(n11044) );
  AND U16566 ( .A(p_input[5030]), .B(p_input[35030]), .Z(n11043) );
  AND U16567 ( .A(n11045), .B(n11046), .Z(o[502]) );
  AND U16568 ( .A(p_input[20502]), .B(p_input[10502]), .Z(n11046) );
  AND U16569 ( .A(p_input[502]), .B(p_input[30502]), .Z(n11045) );
  AND U16570 ( .A(n11047), .B(n11048), .Z(o[5029]) );
  AND U16571 ( .A(p_input[25029]), .B(p_input[15029]), .Z(n11048) );
  AND U16572 ( .A(p_input[5029]), .B(p_input[35029]), .Z(n11047) );
  AND U16573 ( .A(n11049), .B(n11050), .Z(o[5028]) );
  AND U16574 ( .A(p_input[25028]), .B(p_input[15028]), .Z(n11050) );
  AND U16575 ( .A(p_input[5028]), .B(p_input[35028]), .Z(n11049) );
  AND U16576 ( .A(n11051), .B(n11052), .Z(o[5027]) );
  AND U16577 ( .A(p_input[25027]), .B(p_input[15027]), .Z(n11052) );
  AND U16578 ( .A(p_input[5027]), .B(p_input[35027]), .Z(n11051) );
  AND U16579 ( .A(n11053), .B(n11054), .Z(o[5026]) );
  AND U16580 ( .A(p_input[25026]), .B(p_input[15026]), .Z(n11054) );
  AND U16581 ( .A(p_input[5026]), .B(p_input[35026]), .Z(n11053) );
  AND U16582 ( .A(n11055), .B(n11056), .Z(o[5025]) );
  AND U16583 ( .A(p_input[25025]), .B(p_input[15025]), .Z(n11056) );
  AND U16584 ( .A(p_input[5025]), .B(p_input[35025]), .Z(n11055) );
  AND U16585 ( .A(n11057), .B(n11058), .Z(o[5024]) );
  AND U16586 ( .A(p_input[25024]), .B(p_input[15024]), .Z(n11058) );
  AND U16587 ( .A(p_input[5024]), .B(p_input[35024]), .Z(n11057) );
  AND U16588 ( .A(n11059), .B(n11060), .Z(o[5023]) );
  AND U16589 ( .A(p_input[25023]), .B(p_input[15023]), .Z(n11060) );
  AND U16590 ( .A(p_input[5023]), .B(p_input[35023]), .Z(n11059) );
  AND U16591 ( .A(n11061), .B(n11062), .Z(o[5022]) );
  AND U16592 ( .A(p_input[25022]), .B(p_input[15022]), .Z(n11062) );
  AND U16593 ( .A(p_input[5022]), .B(p_input[35022]), .Z(n11061) );
  AND U16594 ( .A(n11063), .B(n11064), .Z(o[5021]) );
  AND U16595 ( .A(p_input[25021]), .B(p_input[15021]), .Z(n11064) );
  AND U16596 ( .A(p_input[5021]), .B(p_input[35021]), .Z(n11063) );
  AND U16597 ( .A(n11065), .B(n11066), .Z(o[5020]) );
  AND U16598 ( .A(p_input[25020]), .B(p_input[15020]), .Z(n11066) );
  AND U16599 ( .A(p_input[5020]), .B(p_input[35020]), .Z(n11065) );
  AND U16600 ( .A(n11067), .B(n11068), .Z(o[501]) );
  AND U16601 ( .A(p_input[20501]), .B(p_input[10501]), .Z(n11068) );
  AND U16602 ( .A(p_input[501]), .B(p_input[30501]), .Z(n11067) );
  AND U16603 ( .A(n11069), .B(n11070), .Z(o[5019]) );
  AND U16604 ( .A(p_input[25019]), .B(p_input[15019]), .Z(n11070) );
  AND U16605 ( .A(p_input[5019]), .B(p_input[35019]), .Z(n11069) );
  AND U16606 ( .A(n11071), .B(n11072), .Z(o[5018]) );
  AND U16607 ( .A(p_input[25018]), .B(p_input[15018]), .Z(n11072) );
  AND U16608 ( .A(p_input[5018]), .B(p_input[35018]), .Z(n11071) );
  AND U16609 ( .A(n11073), .B(n11074), .Z(o[5017]) );
  AND U16610 ( .A(p_input[25017]), .B(p_input[15017]), .Z(n11074) );
  AND U16611 ( .A(p_input[5017]), .B(p_input[35017]), .Z(n11073) );
  AND U16612 ( .A(n11075), .B(n11076), .Z(o[5016]) );
  AND U16613 ( .A(p_input[25016]), .B(p_input[15016]), .Z(n11076) );
  AND U16614 ( .A(p_input[5016]), .B(p_input[35016]), .Z(n11075) );
  AND U16615 ( .A(n11077), .B(n11078), .Z(o[5015]) );
  AND U16616 ( .A(p_input[25015]), .B(p_input[15015]), .Z(n11078) );
  AND U16617 ( .A(p_input[5015]), .B(p_input[35015]), .Z(n11077) );
  AND U16618 ( .A(n11079), .B(n11080), .Z(o[5014]) );
  AND U16619 ( .A(p_input[25014]), .B(p_input[15014]), .Z(n11080) );
  AND U16620 ( .A(p_input[5014]), .B(p_input[35014]), .Z(n11079) );
  AND U16621 ( .A(n11081), .B(n11082), .Z(o[5013]) );
  AND U16622 ( .A(p_input[25013]), .B(p_input[15013]), .Z(n11082) );
  AND U16623 ( .A(p_input[5013]), .B(p_input[35013]), .Z(n11081) );
  AND U16624 ( .A(n11083), .B(n11084), .Z(o[5012]) );
  AND U16625 ( .A(p_input[25012]), .B(p_input[15012]), .Z(n11084) );
  AND U16626 ( .A(p_input[5012]), .B(p_input[35012]), .Z(n11083) );
  AND U16627 ( .A(n11085), .B(n11086), .Z(o[5011]) );
  AND U16628 ( .A(p_input[25011]), .B(p_input[15011]), .Z(n11086) );
  AND U16629 ( .A(p_input[5011]), .B(p_input[35011]), .Z(n11085) );
  AND U16630 ( .A(n11087), .B(n11088), .Z(o[5010]) );
  AND U16631 ( .A(p_input[25010]), .B(p_input[15010]), .Z(n11088) );
  AND U16632 ( .A(p_input[5010]), .B(p_input[35010]), .Z(n11087) );
  AND U16633 ( .A(n11089), .B(n11090), .Z(o[500]) );
  AND U16634 ( .A(p_input[20500]), .B(p_input[10500]), .Z(n11090) );
  AND U16635 ( .A(p_input[500]), .B(p_input[30500]), .Z(n11089) );
  AND U16636 ( .A(n11091), .B(n11092), .Z(o[5009]) );
  AND U16637 ( .A(p_input[25009]), .B(p_input[15009]), .Z(n11092) );
  AND U16638 ( .A(p_input[5009]), .B(p_input[35009]), .Z(n11091) );
  AND U16639 ( .A(n11093), .B(n11094), .Z(o[5008]) );
  AND U16640 ( .A(p_input[25008]), .B(p_input[15008]), .Z(n11094) );
  AND U16641 ( .A(p_input[5008]), .B(p_input[35008]), .Z(n11093) );
  AND U16642 ( .A(n11095), .B(n11096), .Z(o[5007]) );
  AND U16643 ( .A(p_input[25007]), .B(p_input[15007]), .Z(n11096) );
  AND U16644 ( .A(p_input[5007]), .B(p_input[35007]), .Z(n11095) );
  AND U16645 ( .A(n11097), .B(n11098), .Z(o[5006]) );
  AND U16646 ( .A(p_input[25006]), .B(p_input[15006]), .Z(n11098) );
  AND U16647 ( .A(p_input[5006]), .B(p_input[35006]), .Z(n11097) );
  AND U16648 ( .A(n11099), .B(n11100), .Z(o[5005]) );
  AND U16649 ( .A(p_input[25005]), .B(p_input[15005]), .Z(n11100) );
  AND U16650 ( .A(p_input[5005]), .B(p_input[35005]), .Z(n11099) );
  AND U16651 ( .A(n11101), .B(n11102), .Z(o[5004]) );
  AND U16652 ( .A(p_input[25004]), .B(p_input[15004]), .Z(n11102) );
  AND U16653 ( .A(p_input[5004]), .B(p_input[35004]), .Z(n11101) );
  AND U16654 ( .A(n11103), .B(n11104), .Z(o[5003]) );
  AND U16655 ( .A(p_input[25003]), .B(p_input[15003]), .Z(n11104) );
  AND U16656 ( .A(p_input[5003]), .B(p_input[35003]), .Z(n11103) );
  AND U16657 ( .A(n11105), .B(n11106), .Z(o[5002]) );
  AND U16658 ( .A(p_input[25002]), .B(p_input[15002]), .Z(n11106) );
  AND U16659 ( .A(p_input[5002]), .B(p_input[35002]), .Z(n11105) );
  AND U16660 ( .A(n11107), .B(n11108), .Z(o[5001]) );
  AND U16661 ( .A(p_input[25001]), .B(p_input[15001]), .Z(n11108) );
  AND U16662 ( .A(p_input[5001]), .B(p_input[35001]), .Z(n11107) );
  AND U16663 ( .A(n11109), .B(n11110), .Z(o[5000]) );
  AND U16664 ( .A(p_input[25000]), .B(p_input[15000]), .Z(n11110) );
  AND U16665 ( .A(p_input[5000]), .B(p_input[35000]), .Z(n11109) );
  AND U16666 ( .A(n11111), .B(n11112), .Z(o[4]) );
  AND U16667 ( .A(p_input[20004]), .B(p_input[10004]), .Z(n11112) );
  AND U16668 ( .A(p_input[4]), .B(p_input[30004]), .Z(n11111) );
  AND U16669 ( .A(n11113), .B(n11114), .Z(o[49]) );
  AND U16670 ( .A(p_input[20049]), .B(p_input[10049]), .Z(n11114) );
  AND U16671 ( .A(p_input[49]), .B(p_input[30049]), .Z(n11113) );
  AND U16672 ( .A(n11115), .B(n11116), .Z(o[499]) );
  AND U16673 ( .A(p_input[20499]), .B(p_input[10499]), .Z(n11116) );
  AND U16674 ( .A(p_input[499]), .B(p_input[30499]), .Z(n11115) );
  AND U16675 ( .A(n11117), .B(n11118), .Z(o[4999]) );
  AND U16676 ( .A(p_input[24999]), .B(p_input[14999]), .Z(n11118) );
  AND U16677 ( .A(p_input[4999]), .B(p_input[34999]), .Z(n11117) );
  AND U16678 ( .A(n11119), .B(n11120), .Z(o[4998]) );
  AND U16679 ( .A(p_input[24998]), .B(p_input[14998]), .Z(n11120) );
  AND U16680 ( .A(p_input[4998]), .B(p_input[34998]), .Z(n11119) );
  AND U16681 ( .A(n11121), .B(n11122), .Z(o[4997]) );
  AND U16682 ( .A(p_input[24997]), .B(p_input[14997]), .Z(n11122) );
  AND U16683 ( .A(p_input[4997]), .B(p_input[34997]), .Z(n11121) );
  AND U16684 ( .A(n11123), .B(n11124), .Z(o[4996]) );
  AND U16685 ( .A(p_input[24996]), .B(p_input[14996]), .Z(n11124) );
  AND U16686 ( .A(p_input[4996]), .B(p_input[34996]), .Z(n11123) );
  AND U16687 ( .A(n11125), .B(n11126), .Z(o[4995]) );
  AND U16688 ( .A(p_input[24995]), .B(p_input[14995]), .Z(n11126) );
  AND U16689 ( .A(p_input[4995]), .B(p_input[34995]), .Z(n11125) );
  AND U16690 ( .A(n11127), .B(n11128), .Z(o[4994]) );
  AND U16691 ( .A(p_input[24994]), .B(p_input[14994]), .Z(n11128) );
  AND U16692 ( .A(p_input[4994]), .B(p_input[34994]), .Z(n11127) );
  AND U16693 ( .A(n11129), .B(n11130), .Z(o[4993]) );
  AND U16694 ( .A(p_input[24993]), .B(p_input[14993]), .Z(n11130) );
  AND U16695 ( .A(p_input[4993]), .B(p_input[34993]), .Z(n11129) );
  AND U16696 ( .A(n11131), .B(n11132), .Z(o[4992]) );
  AND U16697 ( .A(p_input[24992]), .B(p_input[14992]), .Z(n11132) );
  AND U16698 ( .A(p_input[4992]), .B(p_input[34992]), .Z(n11131) );
  AND U16699 ( .A(n11133), .B(n11134), .Z(o[4991]) );
  AND U16700 ( .A(p_input[24991]), .B(p_input[14991]), .Z(n11134) );
  AND U16701 ( .A(p_input[4991]), .B(p_input[34991]), .Z(n11133) );
  AND U16702 ( .A(n11135), .B(n11136), .Z(o[4990]) );
  AND U16703 ( .A(p_input[24990]), .B(p_input[14990]), .Z(n11136) );
  AND U16704 ( .A(p_input[4990]), .B(p_input[34990]), .Z(n11135) );
  AND U16705 ( .A(n11137), .B(n11138), .Z(o[498]) );
  AND U16706 ( .A(p_input[20498]), .B(p_input[10498]), .Z(n11138) );
  AND U16707 ( .A(p_input[498]), .B(p_input[30498]), .Z(n11137) );
  AND U16708 ( .A(n11139), .B(n11140), .Z(o[4989]) );
  AND U16709 ( .A(p_input[24989]), .B(p_input[14989]), .Z(n11140) );
  AND U16710 ( .A(p_input[4989]), .B(p_input[34989]), .Z(n11139) );
  AND U16711 ( .A(n11141), .B(n11142), .Z(o[4988]) );
  AND U16712 ( .A(p_input[24988]), .B(p_input[14988]), .Z(n11142) );
  AND U16713 ( .A(p_input[4988]), .B(p_input[34988]), .Z(n11141) );
  AND U16714 ( .A(n11143), .B(n11144), .Z(o[4987]) );
  AND U16715 ( .A(p_input[24987]), .B(p_input[14987]), .Z(n11144) );
  AND U16716 ( .A(p_input[4987]), .B(p_input[34987]), .Z(n11143) );
  AND U16717 ( .A(n11145), .B(n11146), .Z(o[4986]) );
  AND U16718 ( .A(p_input[24986]), .B(p_input[14986]), .Z(n11146) );
  AND U16719 ( .A(p_input[4986]), .B(p_input[34986]), .Z(n11145) );
  AND U16720 ( .A(n11147), .B(n11148), .Z(o[4985]) );
  AND U16721 ( .A(p_input[24985]), .B(p_input[14985]), .Z(n11148) );
  AND U16722 ( .A(p_input[4985]), .B(p_input[34985]), .Z(n11147) );
  AND U16723 ( .A(n11149), .B(n11150), .Z(o[4984]) );
  AND U16724 ( .A(p_input[24984]), .B(p_input[14984]), .Z(n11150) );
  AND U16725 ( .A(p_input[4984]), .B(p_input[34984]), .Z(n11149) );
  AND U16726 ( .A(n11151), .B(n11152), .Z(o[4983]) );
  AND U16727 ( .A(p_input[24983]), .B(p_input[14983]), .Z(n11152) );
  AND U16728 ( .A(p_input[4983]), .B(p_input[34983]), .Z(n11151) );
  AND U16729 ( .A(n11153), .B(n11154), .Z(o[4982]) );
  AND U16730 ( .A(p_input[24982]), .B(p_input[14982]), .Z(n11154) );
  AND U16731 ( .A(p_input[4982]), .B(p_input[34982]), .Z(n11153) );
  AND U16732 ( .A(n11155), .B(n11156), .Z(o[4981]) );
  AND U16733 ( .A(p_input[24981]), .B(p_input[14981]), .Z(n11156) );
  AND U16734 ( .A(p_input[4981]), .B(p_input[34981]), .Z(n11155) );
  AND U16735 ( .A(n11157), .B(n11158), .Z(o[4980]) );
  AND U16736 ( .A(p_input[24980]), .B(p_input[14980]), .Z(n11158) );
  AND U16737 ( .A(p_input[4980]), .B(p_input[34980]), .Z(n11157) );
  AND U16738 ( .A(n11159), .B(n11160), .Z(o[497]) );
  AND U16739 ( .A(p_input[20497]), .B(p_input[10497]), .Z(n11160) );
  AND U16740 ( .A(p_input[497]), .B(p_input[30497]), .Z(n11159) );
  AND U16741 ( .A(n11161), .B(n11162), .Z(o[4979]) );
  AND U16742 ( .A(p_input[24979]), .B(p_input[14979]), .Z(n11162) );
  AND U16743 ( .A(p_input[4979]), .B(p_input[34979]), .Z(n11161) );
  AND U16744 ( .A(n11163), .B(n11164), .Z(o[4978]) );
  AND U16745 ( .A(p_input[24978]), .B(p_input[14978]), .Z(n11164) );
  AND U16746 ( .A(p_input[4978]), .B(p_input[34978]), .Z(n11163) );
  AND U16747 ( .A(n11165), .B(n11166), .Z(o[4977]) );
  AND U16748 ( .A(p_input[24977]), .B(p_input[14977]), .Z(n11166) );
  AND U16749 ( .A(p_input[4977]), .B(p_input[34977]), .Z(n11165) );
  AND U16750 ( .A(n11167), .B(n11168), .Z(o[4976]) );
  AND U16751 ( .A(p_input[24976]), .B(p_input[14976]), .Z(n11168) );
  AND U16752 ( .A(p_input[4976]), .B(p_input[34976]), .Z(n11167) );
  AND U16753 ( .A(n11169), .B(n11170), .Z(o[4975]) );
  AND U16754 ( .A(p_input[24975]), .B(p_input[14975]), .Z(n11170) );
  AND U16755 ( .A(p_input[4975]), .B(p_input[34975]), .Z(n11169) );
  AND U16756 ( .A(n11171), .B(n11172), .Z(o[4974]) );
  AND U16757 ( .A(p_input[24974]), .B(p_input[14974]), .Z(n11172) );
  AND U16758 ( .A(p_input[4974]), .B(p_input[34974]), .Z(n11171) );
  AND U16759 ( .A(n11173), .B(n11174), .Z(o[4973]) );
  AND U16760 ( .A(p_input[24973]), .B(p_input[14973]), .Z(n11174) );
  AND U16761 ( .A(p_input[4973]), .B(p_input[34973]), .Z(n11173) );
  AND U16762 ( .A(n11175), .B(n11176), .Z(o[4972]) );
  AND U16763 ( .A(p_input[24972]), .B(p_input[14972]), .Z(n11176) );
  AND U16764 ( .A(p_input[4972]), .B(p_input[34972]), .Z(n11175) );
  AND U16765 ( .A(n11177), .B(n11178), .Z(o[4971]) );
  AND U16766 ( .A(p_input[24971]), .B(p_input[14971]), .Z(n11178) );
  AND U16767 ( .A(p_input[4971]), .B(p_input[34971]), .Z(n11177) );
  AND U16768 ( .A(n11179), .B(n11180), .Z(o[4970]) );
  AND U16769 ( .A(p_input[24970]), .B(p_input[14970]), .Z(n11180) );
  AND U16770 ( .A(p_input[4970]), .B(p_input[34970]), .Z(n11179) );
  AND U16771 ( .A(n11181), .B(n11182), .Z(o[496]) );
  AND U16772 ( .A(p_input[20496]), .B(p_input[10496]), .Z(n11182) );
  AND U16773 ( .A(p_input[496]), .B(p_input[30496]), .Z(n11181) );
  AND U16774 ( .A(n11183), .B(n11184), .Z(o[4969]) );
  AND U16775 ( .A(p_input[24969]), .B(p_input[14969]), .Z(n11184) );
  AND U16776 ( .A(p_input[4969]), .B(p_input[34969]), .Z(n11183) );
  AND U16777 ( .A(n11185), .B(n11186), .Z(o[4968]) );
  AND U16778 ( .A(p_input[24968]), .B(p_input[14968]), .Z(n11186) );
  AND U16779 ( .A(p_input[4968]), .B(p_input[34968]), .Z(n11185) );
  AND U16780 ( .A(n11187), .B(n11188), .Z(o[4967]) );
  AND U16781 ( .A(p_input[24967]), .B(p_input[14967]), .Z(n11188) );
  AND U16782 ( .A(p_input[4967]), .B(p_input[34967]), .Z(n11187) );
  AND U16783 ( .A(n11189), .B(n11190), .Z(o[4966]) );
  AND U16784 ( .A(p_input[24966]), .B(p_input[14966]), .Z(n11190) );
  AND U16785 ( .A(p_input[4966]), .B(p_input[34966]), .Z(n11189) );
  AND U16786 ( .A(n11191), .B(n11192), .Z(o[4965]) );
  AND U16787 ( .A(p_input[24965]), .B(p_input[14965]), .Z(n11192) );
  AND U16788 ( .A(p_input[4965]), .B(p_input[34965]), .Z(n11191) );
  AND U16789 ( .A(n11193), .B(n11194), .Z(o[4964]) );
  AND U16790 ( .A(p_input[24964]), .B(p_input[14964]), .Z(n11194) );
  AND U16791 ( .A(p_input[4964]), .B(p_input[34964]), .Z(n11193) );
  AND U16792 ( .A(n11195), .B(n11196), .Z(o[4963]) );
  AND U16793 ( .A(p_input[24963]), .B(p_input[14963]), .Z(n11196) );
  AND U16794 ( .A(p_input[4963]), .B(p_input[34963]), .Z(n11195) );
  AND U16795 ( .A(n11197), .B(n11198), .Z(o[4962]) );
  AND U16796 ( .A(p_input[24962]), .B(p_input[14962]), .Z(n11198) );
  AND U16797 ( .A(p_input[4962]), .B(p_input[34962]), .Z(n11197) );
  AND U16798 ( .A(n11199), .B(n11200), .Z(o[4961]) );
  AND U16799 ( .A(p_input[24961]), .B(p_input[14961]), .Z(n11200) );
  AND U16800 ( .A(p_input[4961]), .B(p_input[34961]), .Z(n11199) );
  AND U16801 ( .A(n11201), .B(n11202), .Z(o[4960]) );
  AND U16802 ( .A(p_input[24960]), .B(p_input[14960]), .Z(n11202) );
  AND U16803 ( .A(p_input[4960]), .B(p_input[34960]), .Z(n11201) );
  AND U16804 ( .A(n11203), .B(n11204), .Z(o[495]) );
  AND U16805 ( .A(p_input[20495]), .B(p_input[10495]), .Z(n11204) );
  AND U16806 ( .A(p_input[495]), .B(p_input[30495]), .Z(n11203) );
  AND U16807 ( .A(n11205), .B(n11206), .Z(o[4959]) );
  AND U16808 ( .A(p_input[24959]), .B(p_input[14959]), .Z(n11206) );
  AND U16809 ( .A(p_input[4959]), .B(p_input[34959]), .Z(n11205) );
  AND U16810 ( .A(n11207), .B(n11208), .Z(o[4958]) );
  AND U16811 ( .A(p_input[24958]), .B(p_input[14958]), .Z(n11208) );
  AND U16812 ( .A(p_input[4958]), .B(p_input[34958]), .Z(n11207) );
  AND U16813 ( .A(n11209), .B(n11210), .Z(o[4957]) );
  AND U16814 ( .A(p_input[24957]), .B(p_input[14957]), .Z(n11210) );
  AND U16815 ( .A(p_input[4957]), .B(p_input[34957]), .Z(n11209) );
  AND U16816 ( .A(n11211), .B(n11212), .Z(o[4956]) );
  AND U16817 ( .A(p_input[24956]), .B(p_input[14956]), .Z(n11212) );
  AND U16818 ( .A(p_input[4956]), .B(p_input[34956]), .Z(n11211) );
  AND U16819 ( .A(n11213), .B(n11214), .Z(o[4955]) );
  AND U16820 ( .A(p_input[24955]), .B(p_input[14955]), .Z(n11214) );
  AND U16821 ( .A(p_input[4955]), .B(p_input[34955]), .Z(n11213) );
  AND U16822 ( .A(n11215), .B(n11216), .Z(o[4954]) );
  AND U16823 ( .A(p_input[24954]), .B(p_input[14954]), .Z(n11216) );
  AND U16824 ( .A(p_input[4954]), .B(p_input[34954]), .Z(n11215) );
  AND U16825 ( .A(n11217), .B(n11218), .Z(o[4953]) );
  AND U16826 ( .A(p_input[24953]), .B(p_input[14953]), .Z(n11218) );
  AND U16827 ( .A(p_input[4953]), .B(p_input[34953]), .Z(n11217) );
  AND U16828 ( .A(n11219), .B(n11220), .Z(o[4952]) );
  AND U16829 ( .A(p_input[24952]), .B(p_input[14952]), .Z(n11220) );
  AND U16830 ( .A(p_input[4952]), .B(p_input[34952]), .Z(n11219) );
  AND U16831 ( .A(n11221), .B(n11222), .Z(o[4951]) );
  AND U16832 ( .A(p_input[24951]), .B(p_input[14951]), .Z(n11222) );
  AND U16833 ( .A(p_input[4951]), .B(p_input[34951]), .Z(n11221) );
  AND U16834 ( .A(n11223), .B(n11224), .Z(o[4950]) );
  AND U16835 ( .A(p_input[24950]), .B(p_input[14950]), .Z(n11224) );
  AND U16836 ( .A(p_input[4950]), .B(p_input[34950]), .Z(n11223) );
  AND U16837 ( .A(n11225), .B(n11226), .Z(o[494]) );
  AND U16838 ( .A(p_input[20494]), .B(p_input[10494]), .Z(n11226) );
  AND U16839 ( .A(p_input[494]), .B(p_input[30494]), .Z(n11225) );
  AND U16840 ( .A(n11227), .B(n11228), .Z(o[4949]) );
  AND U16841 ( .A(p_input[24949]), .B(p_input[14949]), .Z(n11228) );
  AND U16842 ( .A(p_input[4949]), .B(p_input[34949]), .Z(n11227) );
  AND U16843 ( .A(n11229), .B(n11230), .Z(o[4948]) );
  AND U16844 ( .A(p_input[24948]), .B(p_input[14948]), .Z(n11230) );
  AND U16845 ( .A(p_input[4948]), .B(p_input[34948]), .Z(n11229) );
  AND U16846 ( .A(n11231), .B(n11232), .Z(o[4947]) );
  AND U16847 ( .A(p_input[24947]), .B(p_input[14947]), .Z(n11232) );
  AND U16848 ( .A(p_input[4947]), .B(p_input[34947]), .Z(n11231) );
  AND U16849 ( .A(n11233), .B(n11234), .Z(o[4946]) );
  AND U16850 ( .A(p_input[24946]), .B(p_input[14946]), .Z(n11234) );
  AND U16851 ( .A(p_input[4946]), .B(p_input[34946]), .Z(n11233) );
  AND U16852 ( .A(n11235), .B(n11236), .Z(o[4945]) );
  AND U16853 ( .A(p_input[24945]), .B(p_input[14945]), .Z(n11236) );
  AND U16854 ( .A(p_input[4945]), .B(p_input[34945]), .Z(n11235) );
  AND U16855 ( .A(n11237), .B(n11238), .Z(o[4944]) );
  AND U16856 ( .A(p_input[24944]), .B(p_input[14944]), .Z(n11238) );
  AND U16857 ( .A(p_input[4944]), .B(p_input[34944]), .Z(n11237) );
  AND U16858 ( .A(n11239), .B(n11240), .Z(o[4943]) );
  AND U16859 ( .A(p_input[24943]), .B(p_input[14943]), .Z(n11240) );
  AND U16860 ( .A(p_input[4943]), .B(p_input[34943]), .Z(n11239) );
  AND U16861 ( .A(n11241), .B(n11242), .Z(o[4942]) );
  AND U16862 ( .A(p_input[24942]), .B(p_input[14942]), .Z(n11242) );
  AND U16863 ( .A(p_input[4942]), .B(p_input[34942]), .Z(n11241) );
  AND U16864 ( .A(n11243), .B(n11244), .Z(o[4941]) );
  AND U16865 ( .A(p_input[24941]), .B(p_input[14941]), .Z(n11244) );
  AND U16866 ( .A(p_input[4941]), .B(p_input[34941]), .Z(n11243) );
  AND U16867 ( .A(n11245), .B(n11246), .Z(o[4940]) );
  AND U16868 ( .A(p_input[24940]), .B(p_input[14940]), .Z(n11246) );
  AND U16869 ( .A(p_input[4940]), .B(p_input[34940]), .Z(n11245) );
  AND U16870 ( .A(n11247), .B(n11248), .Z(o[493]) );
  AND U16871 ( .A(p_input[20493]), .B(p_input[10493]), .Z(n11248) );
  AND U16872 ( .A(p_input[493]), .B(p_input[30493]), .Z(n11247) );
  AND U16873 ( .A(n11249), .B(n11250), .Z(o[4939]) );
  AND U16874 ( .A(p_input[24939]), .B(p_input[14939]), .Z(n11250) );
  AND U16875 ( .A(p_input[4939]), .B(p_input[34939]), .Z(n11249) );
  AND U16876 ( .A(n11251), .B(n11252), .Z(o[4938]) );
  AND U16877 ( .A(p_input[24938]), .B(p_input[14938]), .Z(n11252) );
  AND U16878 ( .A(p_input[4938]), .B(p_input[34938]), .Z(n11251) );
  AND U16879 ( .A(n11253), .B(n11254), .Z(o[4937]) );
  AND U16880 ( .A(p_input[24937]), .B(p_input[14937]), .Z(n11254) );
  AND U16881 ( .A(p_input[4937]), .B(p_input[34937]), .Z(n11253) );
  AND U16882 ( .A(n11255), .B(n11256), .Z(o[4936]) );
  AND U16883 ( .A(p_input[24936]), .B(p_input[14936]), .Z(n11256) );
  AND U16884 ( .A(p_input[4936]), .B(p_input[34936]), .Z(n11255) );
  AND U16885 ( .A(n11257), .B(n11258), .Z(o[4935]) );
  AND U16886 ( .A(p_input[24935]), .B(p_input[14935]), .Z(n11258) );
  AND U16887 ( .A(p_input[4935]), .B(p_input[34935]), .Z(n11257) );
  AND U16888 ( .A(n11259), .B(n11260), .Z(o[4934]) );
  AND U16889 ( .A(p_input[24934]), .B(p_input[14934]), .Z(n11260) );
  AND U16890 ( .A(p_input[4934]), .B(p_input[34934]), .Z(n11259) );
  AND U16891 ( .A(n11261), .B(n11262), .Z(o[4933]) );
  AND U16892 ( .A(p_input[24933]), .B(p_input[14933]), .Z(n11262) );
  AND U16893 ( .A(p_input[4933]), .B(p_input[34933]), .Z(n11261) );
  AND U16894 ( .A(n11263), .B(n11264), .Z(o[4932]) );
  AND U16895 ( .A(p_input[24932]), .B(p_input[14932]), .Z(n11264) );
  AND U16896 ( .A(p_input[4932]), .B(p_input[34932]), .Z(n11263) );
  AND U16897 ( .A(n11265), .B(n11266), .Z(o[4931]) );
  AND U16898 ( .A(p_input[24931]), .B(p_input[14931]), .Z(n11266) );
  AND U16899 ( .A(p_input[4931]), .B(p_input[34931]), .Z(n11265) );
  AND U16900 ( .A(n11267), .B(n11268), .Z(o[4930]) );
  AND U16901 ( .A(p_input[24930]), .B(p_input[14930]), .Z(n11268) );
  AND U16902 ( .A(p_input[4930]), .B(p_input[34930]), .Z(n11267) );
  AND U16903 ( .A(n11269), .B(n11270), .Z(o[492]) );
  AND U16904 ( .A(p_input[20492]), .B(p_input[10492]), .Z(n11270) );
  AND U16905 ( .A(p_input[492]), .B(p_input[30492]), .Z(n11269) );
  AND U16906 ( .A(n11271), .B(n11272), .Z(o[4929]) );
  AND U16907 ( .A(p_input[24929]), .B(p_input[14929]), .Z(n11272) );
  AND U16908 ( .A(p_input[4929]), .B(p_input[34929]), .Z(n11271) );
  AND U16909 ( .A(n11273), .B(n11274), .Z(o[4928]) );
  AND U16910 ( .A(p_input[24928]), .B(p_input[14928]), .Z(n11274) );
  AND U16911 ( .A(p_input[4928]), .B(p_input[34928]), .Z(n11273) );
  AND U16912 ( .A(n11275), .B(n11276), .Z(o[4927]) );
  AND U16913 ( .A(p_input[24927]), .B(p_input[14927]), .Z(n11276) );
  AND U16914 ( .A(p_input[4927]), .B(p_input[34927]), .Z(n11275) );
  AND U16915 ( .A(n11277), .B(n11278), .Z(o[4926]) );
  AND U16916 ( .A(p_input[24926]), .B(p_input[14926]), .Z(n11278) );
  AND U16917 ( .A(p_input[4926]), .B(p_input[34926]), .Z(n11277) );
  AND U16918 ( .A(n11279), .B(n11280), .Z(o[4925]) );
  AND U16919 ( .A(p_input[24925]), .B(p_input[14925]), .Z(n11280) );
  AND U16920 ( .A(p_input[4925]), .B(p_input[34925]), .Z(n11279) );
  AND U16921 ( .A(n11281), .B(n11282), .Z(o[4924]) );
  AND U16922 ( .A(p_input[24924]), .B(p_input[14924]), .Z(n11282) );
  AND U16923 ( .A(p_input[4924]), .B(p_input[34924]), .Z(n11281) );
  AND U16924 ( .A(n11283), .B(n11284), .Z(o[4923]) );
  AND U16925 ( .A(p_input[24923]), .B(p_input[14923]), .Z(n11284) );
  AND U16926 ( .A(p_input[4923]), .B(p_input[34923]), .Z(n11283) );
  AND U16927 ( .A(n11285), .B(n11286), .Z(o[4922]) );
  AND U16928 ( .A(p_input[24922]), .B(p_input[14922]), .Z(n11286) );
  AND U16929 ( .A(p_input[4922]), .B(p_input[34922]), .Z(n11285) );
  AND U16930 ( .A(n11287), .B(n11288), .Z(o[4921]) );
  AND U16931 ( .A(p_input[24921]), .B(p_input[14921]), .Z(n11288) );
  AND U16932 ( .A(p_input[4921]), .B(p_input[34921]), .Z(n11287) );
  AND U16933 ( .A(n11289), .B(n11290), .Z(o[4920]) );
  AND U16934 ( .A(p_input[24920]), .B(p_input[14920]), .Z(n11290) );
  AND U16935 ( .A(p_input[4920]), .B(p_input[34920]), .Z(n11289) );
  AND U16936 ( .A(n11291), .B(n11292), .Z(o[491]) );
  AND U16937 ( .A(p_input[20491]), .B(p_input[10491]), .Z(n11292) );
  AND U16938 ( .A(p_input[491]), .B(p_input[30491]), .Z(n11291) );
  AND U16939 ( .A(n11293), .B(n11294), .Z(o[4919]) );
  AND U16940 ( .A(p_input[24919]), .B(p_input[14919]), .Z(n11294) );
  AND U16941 ( .A(p_input[4919]), .B(p_input[34919]), .Z(n11293) );
  AND U16942 ( .A(n11295), .B(n11296), .Z(o[4918]) );
  AND U16943 ( .A(p_input[24918]), .B(p_input[14918]), .Z(n11296) );
  AND U16944 ( .A(p_input[4918]), .B(p_input[34918]), .Z(n11295) );
  AND U16945 ( .A(n11297), .B(n11298), .Z(o[4917]) );
  AND U16946 ( .A(p_input[24917]), .B(p_input[14917]), .Z(n11298) );
  AND U16947 ( .A(p_input[4917]), .B(p_input[34917]), .Z(n11297) );
  AND U16948 ( .A(n11299), .B(n11300), .Z(o[4916]) );
  AND U16949 ( .A(p_input[24916]), .B(p_input[14916]), .Z(n11300) );
  AND U16950 ( .A(p_input[4916]), .B(p_input[34916]), .Z(n11299) );
  AND U16951 ( .A(n11301), .B(n11302), .Z(o[4915]) );
  AND U16952 ( .A(p_input[24915]), .B(p_input[14915]), .Z(n11302) );
  AND U16953 ( .A(p_input[4915]), .B(p_input[34915]), .Z(n11301) );
  AND U16954 ( .A(n11303), .B(n11304), .Z(o[4914]) );
  AND U16955 ( .A(p_input[24914]), .B(p_input[14914]), .Z(n11304) );
  AND U16956 ( .A(p_input[4914]), .B(p_input[34914]), .Z(n11303) );
  AND U16957 ( .A(n11305), .B(n11306), .Z(o[4913]) );
  AND U16958 ( .A(p_input[24913]), .B(p_input[14913]), .Z(n11306) );
  AND U16959 ( .A(p_input[4913]), .B(p_input[34913]), .Z(n11305) );
  AND U16960 ( .A(n11307), .B(n11308), .Z(o[4912]) );
  AND U16961 ( .A(p_input[24912]), .B(p_input[14912]), .Z(n11308) );
  AND U16962 ( .A(p_input[4912]), .B(p_input[34912]), .Z(n11307) );
  AND U16963 ( .A(n11309), .B(n11310), .Z(o[4911]) );
  AND U16964 ( .A(p_input[24911]), .B(p_input[14911]), .Z(n11310) );
  AND U16965 ( .A(p_input[4911]), .B(p_input[34911]), .Z(n11309) );
  AND U16966 ( .A(n11311), .B(n11312), .Z(o[4910]) );
  AND U16967 ( .A(p_input[24910]), .B(p_input[14910]), .Z(n11312) );
  AND U16968 ( .A(p_input[4910]), .B(p_input[34910]), .Z(n11311) );
  AND U16969 ( .A(n11313), .B(n11314), .Z(o[490]) );
  AND U16970 ( .A(p_input[20490]), .B(p_input[10490]), .Z(n11314) );
  AND U16971 ( .A(p_input[490]), .B(p_input[30490]), .Z(n11313) );
  AND U16972 ( .A(n11315), .B(n11316), .Z(o[4909]) );
  AND U16973 ( .A(p_input[24909]), .B(p_input[14909]), .Z(n11316) );
  AND U16974 ( .A(p_input[4909]), .B(p_input[34909]), .Z(n11315) );
  AND U16975 ( .A(n11317), .B(n11318), .Z(o[4908]) );
  AND U16976 ( .A(p_input[24908]), .B(p_input[14908]), .Z(n11318) );
  AND U16977 ( .A(p_input[4908]), .B(p_input[34908]), .Z(n11317) );
  AND U16978 ( .A(n11319), .B(n11320), .Z(o[4907]) );
  AND U16979 ( .A(p_input[24907]), .B(p_input[14907]), .Z(n11320) );
  AND U16980 ( .A(p_input[4907]), .B(p_input[34907]), .Z(n11319) );
  AND U16981 ( .A(n11321), .B(n11322), .Z(o[4906]) );
  AND U16982 ( .A(p_input[24906]), .B(p_input[14906]), .Z(n11322) );
  AND U16983 ( .A(p_input[4906]), .B(p_input[34906]), .Z(n11321) );
  AND U16984 ( .A(n11323), .B(n11324), .Z(o[4905]) );
  AND U16985 ( .A(p_input[24905]), .B(p_input[14905]), .Z(n11324) );
  AND U16986 ( .A(p_input[4905]), .B(p_input[34905]), .Z(n11323) );
  AND U16987 ( .A(n11325), .B(n11326), .Z(o[4904]) );
  AND U16988 ( .A(p_input[24904]), .B(p_input[14904]), .Z(n11326) );
  AND U16989 ( .A(p_input[4904]), .B(p_input[34904]), .Z(n11325) );
  AND U16990 ( .A(n11327), .B(n11328), .Z(o[4903]) );
  AND U16991 ( .A(p_input[24903]), .B(p_input[14903]), .Z(n11328) );
  AND U16992 ( .A(p_input[4903]), .B(p_input[34903]), .Z(n11327) );
  AND U16993 ( .A(n11329), .B(n11330), .Z(o[4902]) );
  AND U16994 ( .A(p_input[24902]), .B(p_input[14902]), .Z(n11330) );
  AND U16995 ( .A(p_input[4902]), .B(p_input[34902]), .Z(n11329) );
  AND U16996 ( .A(n11331), .B(n11332), .Z(o[4901]) );
  AND U16997 ( .A(p_input[24901]), .B(p_input[14901]), .Z(n11332) );
  AND U16998 ( .A(p_input[4901]), .B(p_input[34901]), .Z(n11331) );
  AND U16999 ( .A(n11333), .B(n11334), .Z(o[4900]) );
  AND U17000 ( .A(p_input[24900]), .B(p_input[14900]), .Z(n11334) );
  AND U17001 ( .A(p_input[4900]), .B(p_input[34900]), .Z(n11333) );
  AND U17002 ( .A(n11335), .B(n11336), .Z(o[48]) );
  AND U17003 ( .A(p_input[20048]), .B(p_input[10048]), .Z(n11336) );
  AND U17004 ( .A(p_input[48]), .B(p_input[30048]), .Z(n11335) );
  AND U17005 ( .A(n11337), .B(n11338), .Z(o[489]) );
  AND U17006 ( .A(p_input[20489]), .B(p_input[10489]), .Z(n11338) );
  AND U17007 ( .A(p_input[489]), .B(p_input[30489]), .Z(n11337) );
  AND U17008 ( .A(n11339), .B(n11340), .Z(o[4899]) );
  AND U17009 ( .A(p_input[24899]), .B(p_input[14899]), .Z(n11340) );
  AND U17010 ( .A(p_input[4899]), .B(p_input[34899]), .Z(n11339) );
  AND U17011 ( .A(n11341), .B(n11342), .Z(o[4898]) );
  AND U17012 ( .A(p_input[24898]), .B(p_input[14898]), .Z(n11342) );
  AND U17013 ( .A(p_input[4898]), .B(p_input[34898]), .Z(n11341) );
  AND U17014 ( .A(n11343), .B(n11344), .Z(o[4897]) );
  AND U17015 ( .A(p_input[24897]), .B(p_input[14897]), .Z(n11344) );
  AND U17016 ( .A(p_input[4897]), .B(p_input[34897]), .Z(n11343) );
  AND U17017 ( .A(n11345), .B(n11346), .Z(o[4896]) );
  AND U17018 ( .A(p_input[24896]), .B(p_input[14896]), .Z(n11346) );
  AND U17019 ( .A(p_input[4896]), .B(p_input[34896]), .Z(n11345) );
  AND U17020 ( .A(n11347), .B(n11348), .Z(o[4895]) );
  AND U17021 ( .A(p_input[24895]), .B(p_input[14895]), .Z(n11348) );
  AND U17022 ( .A(p_input[4895]), .B(p_input[34895]), .Z(n11347) );
  AND U17023 ( .A(n11349), .B(n11350), .Z(o[4894]) );
  AND U17024 ( .A(p_input[24894]), .B(p_input[14894]), .Z(n11350) );
  AND U17025 ( .A(p_input[4894]), .B(p_input[34894]), .Z(n11349) );
  AND U17026 ( .A(n11351), .B(n11352), .Z(o[4893]) );
  AND U17027 ( .A(p_input[24893]), .B(p_input[14893]), .Z(n11352) );
  AND U17028 ( .A(p_input[4893]), .B(p_input[34893]), .Z(n11351) );
  AND U17029 ( .A(n11353), .B(n11354), .Z(o[4892]) );
  AND U17030 ( .A(p_input[24892]), .B(p_input[14892]), .Z(n11354) );
  AND U17031 ( .A(p_input[4892]), .B(p_input[34892]), .Z(n11353) );
  AND U17032 ( .A(n11355), .B(n11356), .Z(o[4891]) );
  AND U17033 ( .A(p_input[24891]), .B(p_input[14891]), .Z(n11356) );
  AND U17034 ( .A(p_input[4891]), .B(p_input[34891]), .Z(n11355) );
  AND U17035 ( .A(n11357), .B(n11358), .Z(o[4890]) );
  AND U17036 ( .A(p_input[24890]), .B(p_input[14890]), .Z(n11358) );
  AND U17037 ( .A(p_input[4890]), .B(p_input[34890]), .Z(n11357) );
  AND U17038 ( .A(n11359), .B(n11360), .Z(o[488]) );
  AND U17039 ( .A(p_input[20488]), .B(p_input[10488]), .Z(n11360) );
  AND U17040 ( .A(p_input[488]), .B(p_input[30488]), .Z(n11359) );
  AND U17041 ( .A(n11361), .B(n11362), .Z(o[4889]) );
  AND U17042 ( .A(p_input[24889]), .B(p_input[14889]), .Z(n11362) );
  AND U17043 ( .A(p_input[4889]), .B(p_input[34889]), .Z(n11361) );
  AND U17044 ( .A(n11363), .B(n11364), .Z(o[4888]) );
  AND U17045 ( .A(p_input[24888]), .B(p_input[14888]), .Z(n11364) );
  AND U17046 ( .A(p_input[4888]), .B(p_input[34888]), .Z(n11363) );
  AND U17047 ( .A(n11365), .B(n11366), .Z(o[4887]) );
  AND U17048 ( .A(p_input[24887]), .B(p_input[14887]), .Z(n11366) );
  AND U17049 ( .A(p_input[4887]), .B(p_input[34887]), .Z(n11365) );
  AND U17050 ( .A(n11367), .B(n11368), .Z(o[4886]) );
  AND U17051 ( .A(p_input[24886]), .B(p_input[14886]), .Z(n11368) );
  AND U17052 ( .A(p_input[4886]), .B(p_input[34886]), .Z(n11367) );
  AND U17053 ( .A(n11369), .B(n11370), .Z(o[4885]) );
  AND U17054 ( .A(p_input[24885]), .B(p_input[14885]), .Z(n11370) );
  AND U17055 ( .A(p_input[4885]), .B(p_input[34885]), .Z(n11369) );
  AND U17056 ( .A(n11371), .B(n11372), .Z(o[4884]) );
  AND U17057 ( .A(p_input[24884]), .B(p_input[14884]), .Z(n11372) );
  AND U17058 ( .A(p_input[4884]), .B(p_input[34884]), .Z(n11371) );
  AND U17059 ( .A(n11373), .B(n11374), .Z(o[4883]) );
  AND U17060 ( .A(p_input[24883]), .B(p_input[14883]), .Z(n11374) );
  AND U17061 ( .A(p_input[4883]), .B(p_input[34883]), .Z(n11373) );
  AND U17062 ( .A(n11375), .B(n11376), .Z(o[4882]) );
  AND U17063 ( .A(p_input[24882]), .B(p_input[14882]), .Z(n11376) );
  AND U17064 ( .A(p_input[4882]), .B(p_input[34882]), .Z(n11375) );
  AND U17065 ( .A(n11377), .B(n11378), .Z(o[4881]) );
  AND U17066 ( .A(p_input[24881]), .B(p_input[14881]), .Z(n11378) );
  AND U17067 ( .A(p_input[4881]), .B(p_input[34881]), .Z(n11377) );
  AND U17068 ( .A(n11379), .B(n11380), .Z(o[4880]) );
  AND U17069 ( .A(p_input[24880]), .B(p_input[14880]), .Z(n11380) );
  AND U17070 ( .A(p_input[4880]), .B(p_input[34880]), .Z(n11379) );
  AND U17071 ( .A(n11381), .B(n11382), .Z(o[487]) );
  AND U17072 ( .A(p_input[20487]), .B(p_input[10487]), .Z(n11382) );
  AND U17073 ( .A(p_input[487]), .B(p_input[30487]), .Z(n11381) );
  AND U17074 ( .A(n11383), .B(n11384), .Z(o[4879]) );
  AND U17075 ( .A(p_input[24879]), .B(p_input[14879]), .Z(n11384) );
  AND U17076 ( .A(p_input[4879]), .B(p_input[34879]), .Z(n11383) );
  AND U17077 ( .A(n11385), .B(n11386), .Z(o[4878]) );
  AND U17078 ( .A(p_input[24878]), .B(p_input[14878]), .Z(n11386) );
  AND U17079 ( .A(p_input[4878]), .B(p_input[34878]), .Z(n11385) );
  AND U17080 ( .A(n11387), .B(n11388), .Z(o[4877]) );
  AND U17081 ( .A(p_input[24877]), .B(p_input[14877]), .Z(n11388) );
  AND U17082 ( .A(p_input[4877]), .B(p_input[34877]), .Z(n11387) );
  AND U17083 ( .A(n11389), .B(n11390), .Z(o[4876]) );
  AND U17084 ( .A(p_input[24876]), .B(p_input[14876]), .Z(n11390) );
  AND U17085 ( .A(p_input[4876]), .B(p_input[34876]), .Z(n11389) );
  AND U17086 ( .A(n11391), .B(n11392), .Z(o[4875]) );
  AND U17087 ( .A(p_input[24875]), .B(p_input[14875]), .Z(n11392) );
  AND U17088 ( .A(p_input[4875]), .B(p_input[34875]), .Z(n11391) );
  AND U17089 ( .A(n11393), .B(n11394), .Z(o[4874]) );
  AND U17090 ( .A(p_input[24874]), .B(p_input[14874]), .Z(n11394) );
  AND U17091 ( .A(p_input[4874]), .B(p_input[34874]), .Z(n11393) );
  AND U17092 ( .A(n11395), .B(n11396), .Z(o[4873]) );
  AND U17093 ( .A(p_input[24873]), .B(p_input[14873]), .Z(n11396) );
  AND U17094 ( .A(p_input[4873]), .B(p_input[34873]), .Z(n11395) );
  AND U17095 ( .A(n11397), .B(n11398), .Z(o[4872]) );
  AND U17096 ( .A(p_input[24872]), .B(p_input[14872]), .Z(n11398) );
  AND U17097 ( .A(p_input[4872]), .B(p_input[34872]), .Z(n11397) );
  AND U17098 ( .A(n11399), .B(n11400), .Z(o[4871]) );
  AND U17099 ( .A(p_input[24871]), .B(p_input[14871]), .Z(n11400) );
  AND U17100 ( .A(p_input[4871]), .B(p_input[34871]), .Z(n11399) );
  AND U17101 ( .A(n11401), .B(n11402), .Z(o[4870]) );
  AND U17102 ( .A(p_input[24870]), .B(p_input[14870]), .Z(n11402) );
  AND U17103 ( .A(p_input[4870]), .B(p_input[34870]), .Z(n11401) );
  AND U17104 ( .A(n11403), .B(n11404), .Z(o[486]) );
  AND U17105 ( .A(p_input[20486]), .B(p_input[10486]), .Z(n11404) );
  AND U17106 ( .A(p_input[486]), .B(p_input[30486]), .Z(n11403) );
  AND U17107 ( .A(n11405), .B(n11406), .Z(o[4869]) );
  AND U17108 ( .A(p_input[24869]), .B(p_input[14869]), .Z(n11406) );
  AND U17109 ( .A(p_input[4869]), .B(p_input[34869]), .Z(n11405) );
  AND U17110 ( .A(n11407), .B(n11408), .Z(o[4868]) );
  AND U17111 ( .A(p_input[24868]), .B(p_input[14868]), .Z(n11408) );
  AND U17112 ( .A(p_input[4868]), .B(p_input[34868]), .Z(n11407) );
  AND U17113 ( .A(n11409), .B(n11410), .Z(o[4867]) );
  AND U17114 ( .A(p_input[24867]), .B(p_input[14867]), .Z(n11410) );
  AND U17115 ( .A(p_input[4867]), .B(p_input[34867]), .Z(n11409) );
  AND U17116 ( .A(n11411), .B(n11412), .Z(o[4866]) );
  AND U17117 ( .A(p_input[24866]), .B(p_input[14866]), .Z(n11412) );
  AND U17118 ( .A(p_input[4866]), .B(p_input[34866]), .Z(n11411) );
  AND U17119 ( .A(n11413), .B(n11414), .Z(o[4865]) );
  AND U17120 ( .A(p_input[24865]), .B(p_input[14865]), .Z(n11414) );
  AND U17121 ( .A(p_input[4865]), .B(p_input[34865]), .Z(n11413) );
  AND U17122 ( .A(n11415), .B(n11416), .Z(o[4864]) );
  AND U17123 ( .A(p_input[24864]), .B(p_input[14864]), .Z(n11416) );
  AND U17124 ( .A(p_input[4864]), .B(p_input[34864]), .Z(n11415) );
  AND U17125 ( .A(n11417), .B(n11418), .Z(o[4863]) );
  AND U17126 ( .A(p_input[24863]), .B(p_input[14863]), .Z(n11418) );
  AND U17127 ( .A(p_input[4863]), .B(p_input[34863]), .Z(n11417) );
  AND U17128 ( .A(n11419), .B(n11420), .Z(o[4862]) );
  AND U17129 ( .A(p_input[24862]), .B(p_input[14862]), .Z(n11420) );
  AND U17130 ( .A(p_input[4862]), .B(p_input[34862]), .Z(n11419) );
  AND U17131 ( .A(n11421), .B(n11422), .Z(o[4861]) );
  AND U17132 ( .A(p_input[24861]), .B(p_input[14861]), .Z(n11422) );
  AND U17133 ( .A(p_input[4861]), .B(p_input[34861]), .Z(n11421) );
  AND U17134 ( .A(n11423), .B(n11424), .Z(o[4860]) );
  AND U17135 ( .A(p_input[24860]), .B(p_input[14860]), .Z(n11424) );
  AND U17136 ( .A(p_input[4860]), .B(p_input[34860]), .Z(n11423) );
  AND U17137 ( .A(n11425), .B(n11426), .Z(o[485]) );
  AND U17138 ( .A(p_input[20485]), .B(p_input[10485]), .Z(n11426) );
  AND U17139 ( .A(p_input[485]), .B(p_input[30485]), .Z(n11425) );
  AND U17140 ( .A(n11427), .B(n11428), .Z(o[4859]) );
  AND U17141 ( .A(p_input[24859]), .B(p_input[14859]), .Z(n11428) );
  AND U17142 ( .A(p_input[4859]), .B(p_input[34859]), .Z(n11427) );
  AND U17143 ( .A(n11429), .B(n11430), .Z(o[4858]) );
  AND U17144 ( .A(p_input[24858]), .B(p_input[14858]), .Z(n11430) );
  AND U17145 ( .A(p_input[4858]), .B(p_input[34858]), .Z(n11429) );
  AND U17146 ( .A(n11431), .B(n11432), .Z(o[4857]) );
  AND U17147 ( .A(p_input[24857]), .B(p_input[14857]), .Z(n11432) );
  AND U17148 ( .A(p_input[4857]), .B(p_input[34857]), .Z(n11431) );
  AND U17149 ( .A(n11433), .B(n11434), .Z(o[4856]) );
  AND U17150 ( .A(p_input[24856]), .B(p_input[14856]), .Z(n11434) );
  AND U17151 ( .A(p_input[4856]), .B(p_input[34856]), .Z(n11433) );
  AND U17152 ( .A(n11435), .B(n11436), .Z(o[4855]) );
  AND U17153 ( .A(p_input[24855]), .B(p_input[14855]), .Z(n11436) );
  AND U17154 ( .A(p_input[4855]), .B(p_input[34855]), .Z(n11435) );
  AND U17155 ( .A(n11437), .B(n11438), .Z(o[4854]) );
  AND U17156 ( .A(p_input[24854]), .B(p_input[14854]), .Z(n11438) );
  AND U17157 ( .A(p_input[4854]), .B(p_input[34854]), .Z(n11437) );
  AND U17158 ( .A(n11439), .B(n11440), .Z(o[4853]) );
  AND U17159 ( .A(p_input[24853]), .B(p_input[14853]), .Z(n11440) );
  AND U17160 ( .A(p_input[4853]), .B(p_input[34853]), .Z(n11439) );
  AND U17161 ( .A(n11441), .B(n11442), .Z(o[4852]) );
  AND U17162 ( .A(p_input[24852]), .B(p_input[14852]), .Z(n11442) );
  AND U17163 ( .A(p_input[4852]), .B(p_input[34852]), .Z(n11441) );
  AND U17164 ( .A(n11443), .B(n11444), .Z(o[4851]) );
  AND U17165 ( .A(p_input[24851]), .B(p_input[14851]), .Z(n11444) );
  AND U17166 ( .A(p_input[4851]), .B(p_input[34851]), .Z(n11443) );
  AND U17167 ( .A(n11445), .B(n11446), .Z(o[4850]) );
  AND U17168 ( .A(p_input[24850]), .B(p_input[14850]), .Z(n11446) );
  AND U17169 ( .A(p_input[4850]), .B(p_input[34850]), .Z(n11445) );
  AND U17170 ( .A(n11447), .B(n11448), .Z(o[484]) );
  AND U17171 ( .A(p_input[20484]), .B(p_input[10484]), .Z(n11448) );
  AND U17172 ( .A(p_input[484]), .B(p_input[30484]), .Z(n11447) );
  AND U17173 ( .A(n11449), .B(n11450), .Z(o[4849]) );
  AND U17174 ( .A(p_input[24849]), .B(p_input[14849]), .Z(n11450) );
  AND U17175 ( .A(p_input[4849]), .B(p_input[34849]), .Z(n11449) );
  AND U17176 ( .A(n11451), .B(n11452), .Z(o[4848]) );
  AND U17177 ( .A(p_input[24848]), .B(p_input[14848]), .Z(n11452) );
  AND U17178 ( .A(p_input[4848]), .B(p_input[34848]), .Z(n11451) );
  AND U17179 ( .A(n11453), .B(n11454), .Z(o[4847]) );
  AND U17180 ( .A(p_input[24847]), .B(p_input[14847]), .Z(n11454) );
  AND U17181 ( .A(p_input[4847]), .B(p_input[34847]), .Z(n11453) );
  AND U17182 ( .A(n11455), .B(n11456), .Z(o[4846]) );
  AND U17183 ( .A(p_input[24846]), .B(p_input[14846]), .Z(n11456) );
  AND U17184 ( .A(p_input[4846]), .B(p_input[34846]), .Z(n11455) );
  AND U17185 ( .A(n11457), .B(n11458), .Z(o[4845]) );
  AND U17186 ( .A(p_input[24845]), .B(p_input[14845]), .Z(n11458) );
  AND U17187 ( .A(p_input[4845]), .B(p_input[34845]), .Z(n11457) );
  AND U17188 ( .A(n11459), .B(n11460), .Z(o[4844]) );
  AND U17189 ( .A(p_input[24844]), .B(p_input[14844]), .Z(n11460) );
  AND U17190 ( .A(p_input[4844]), .B(p_input[34844]), .Z(n11459) );
  AND U17191 ( .A(n11461), .B(n11462), .Z(o[4843]) );
  AND U17192 ( .A(p_input[24843]), .B(p_input[14843]), .Z(n11462) );
  AND U17193 ( .A(p_input[4843]), .B(p_input[34843]), .Z(n11461) );
  AND U17194 ( .A(n11463), .B(n11464), .Z(o[4842]) );
  AND U17195 ( .A(p_input[24842]), .B(p_input[14842]), .Z(n11464) );
  AND U17196 ( .A(p_input[4842]), .B(p_input[34842]), .Z(n11463) );
  AND U17197 ( .A(n11465), .B(n11466), .Z(o[4841]) );
  AND U17198 ( .A(p_input[24841]), .B(p_input[14841]), .Z(n11466) );
  AND U17199 ( .A(p_input[4841]), .B(p_input[34841]), .Z(n11465) );
  AND U17200 ( .A(n11467), .B(n11468), .Z(o[4840]) );
  AND U17201 ( .A(p_input[24840]), .B(p_input[14840]), .Z(n11468) );
  AND U17202 ( .A(p_input[4840]), .B(p_input[34840]), .Z(n11467) );
  AND U17203 ( .A(n11469), .B(n11470), .Z(o[483]) );
  AND U17204 ( .A(p_input[20483]), .B(p_input[10483]), .Z(n11470) );
  AND U17205 ( .A(p_input[483]), .B(p_input[30483]), .Z(n11469) );
  AND U17206 ( .A(n11471), .B(n11472), .Z(o[4839]) );
  AND U17207 ( .A(p_input[24839]), .B(p_input[14839]), .Z(n11472) );
  AND U17208 ( .A(p_input[4839]), .B(p_input[34839]), .Z(n11471) );
  AND U17209 ( .A(n11473), .B(n11474), .Z(o[4838]) );
  AND U17210 ( .A(p_input[24838]), .B(p_input[14838]), .Z(n11474) );
  AND U17211 ( .A(p_input[4838]), .B(p_input[34838]), .Z(n11473) );
  AND U17212 ( .A(n11475), .B(n11476), .Z(o[4837]) );
  AND U17213 ( .A(p_input[24837]), .B(p_input[14837]), .Z(n11476) );
  AND U17214 ( .A(p_input[4837]), .B(p_input[34837]), .Z(n11475) );
  AND U17215 ( .A(n11477), .B(n11478), .Z(o[4836]) );
  AND U17216 ( .A(p_input[24836]), .B(p_input[14836]), .Z(n11478) );
  AND U17217 ( .A(p_input[4836]), .B(p_input[34836]), .Z(n11477) );
  AND U17218 ( .A(n11479), .B(n11480), .Z(o[4835]) );
  AND U17219 ( .A(p_input[24835]), .B(p_input[14835]), .Z(n11480) );
  AND U17220 ( .A(p_input[4835]), .B(p_input[34835]), .Z(n11479) );
  AND U17221 ( .A(n11481), .B(n11482), .Z(o[4834]) );
  AND U17222 ( .A(p_input[24834]), .B(p_input[14834]), .Z(n11482) );
  AND U17223 ( .A(p_input[4834]), .B(p_input[34834]), .Z(n11481) );
  AND U17224 ( .A(n11483), .B(n11484), .Z(o[4833]) );
  AND U17225 ( .A(p_input[24833]), .B(p_input[14833]), .Z(n11484) );
  AND U17226 ( .A(p_input[4833]), .B(p_input[34833]), .Z(n11483) );
  AND U17227 ( .A(n11485), .B(n11486), .Z(o[4832]) );
  AND U17228 ( .A(p_input[24832]), .B(p_input[14832]), .Z(n11486) );
  AND U17229 ( .A(p_input[4832]), .B(p_input[34832]), .Z(n11485) );
  AND U17230 ( .A(n11487), .B(n11488), .Z(o[4831]) );
  AND U17231 ( .A(p_input[24831]), .B(p_input[14831]), .Z(n11488) );
  AND U17232 ( .A(p_input[4831]), .B(p_input[34831]), .Z(n11487) );
  AND U17233 ( .A(n11489), .B(n11490), .Z(o[4830]) );
  AND U17234 ( .A(p_input[24830]), .B(p_input[14830]), .Z(n11490) );
  AND U17235 ( .A(p_input[4830]), .B(p_input[34830]), .Z(n11489) );
  AND U17236 ( .A(n11491), .B(n11492), .Z(o[482]) );
  AND U17237 ( .A(p_input[20482]), .B(p_input[10482]), .Z(n11492) );
  AND U17238 ( .A(p_input[482]), .B(p_input[30482]), .Z(n11491) );
  AND U17239 ( .A(n11493), .B(n11494), .Z(o[4829]) );
  AND U17240 ( .A(p_input[24829]), .B(p_input[14829]), .Z(n11494) );
  AND U17241 ( .A(p_input[4829]), .B(p_input[34829]), .Z(n11493) );
  AND U17242 ( .A(n11495), .B(n11496), .Z(o[4828]) );
  AND U17243 ( .A(p_input[24828]), .B(p_input[14828]), .Z(n11496) );
  AND U17244 ( .A(p_input[4828]), .B(p_input[34828]), .Z(n11495) );
  AND U17245 ( .A(n11497), .B(n11498), .Z(o[4827]) );
  AND U17246 ( .A(p_input[24827]), .B(p_input[14827]), .Z(n11498) );
  AND U17247 ( .A(p_input[4827]), .B(p_input[34827]), .Z(n11497) );
  AND U17248 ( .A(n11499), .B(n11500), .Z(o[4826]) );
  AND U17249 ( .A(p_input[24826]), .B(p_input[14826]), .Z(n11500) );
  AND U17250 ( .A(p_input[4826]), .B(p_input[34826]), .Z(n11499) );
  AND U17251 ( .A(n11501), .B(n11502), .Z(o[4825]) );
  AND U17252 ( .A(p_input[24825]), .B(p_input[14825]), .Z(n11502) );
  AND U17253 ( .A(p_input[4825]), .B(p_input[34825]), .Z(n11501) );
  AND U17254 ( .A(n11503), .B(n11504), .Z(o[4824]) );
  AND U17255 ( .A(p_input[24824]), .B(p_input[14824]), .Z(n11504) );
  AND U17256 ( .A(p_input[4824]), .B(p_input[34824]), .Z(n11503) );
  AND U17257 ( .A(n11505), .B(n11506), .Z(o[4823]) );
  AND U17258 ( .A(p_input[24823]), .B(p_input[14823]), .Z(n11506) );
  AND U17259 ( .A(p_input[4823]), .B(p_input[34823]), .Z(n11505) );
  AND U17260 ( .A(n11507), .B(n11508), .Z(o[4822]) );
  AND U17261 ( .A(p_input[24822]), .B(p_input[14822]), .Z(n11508) );
  AND U17262 ( .A(p_input[4822]), .B(p_input[34822]), .Z(n11507) );
  AND U17263 ( .A(n11509), .B(n11510), .Z(o[4821]) );
  AND U17264 ( .A(p_input[24821]), .B(p_input[14821]), .Z(n11510) );
  AND U17265 ( .A(p_input[4821]), .B(p_input[34821]), .Z(n11509) );
  AND U17266 ( .A(n11511), .B(n11512), .Z(o[4820]) );
  AND U17267 ( .A(p_input[24820]), .B(p_input[14820]), .Z(n11512) );
  AND U17268 ( .A(p_input[4820]), .B(p_input[34820]), .Z(n11511) );
  AND U17269 ( .A(n11513), .B(n11514), .Z(o[481]) );
  AND U17270 ( .A(p_input[20481]), .B(p_input[10481]), .Z(n11514) );
  AND U17271 ( .A(p_input[481]), .B(p_input[30481]), .Z(n11513) );
  AND U17272 ( .A(n11515), .B(n11516), .Z(o[4819]) );
  AND U17273 ( .A(p_input[24819]), .B(p_input[14819]), .Z(n11516) );
  AND U17274 ( .A(p_input[4819]), .B(p_input[34819]), .Z(n11515) );
  AND U17275 ( .A(n11517), .B(n11518), .Z(o[4818]) );
  AND U17276 ( .A(p_input[24818]), .B(p_input[14818]), .Z(n11518) );
  AND U17277 ( .A(p_input[4818]), .B(p_input[34818]), .Z(n11517) );
  AND U17278 ( .A(n11519), .B(n11520), .Z(o[4817]) );
  AND U17279 ( .A(p_input[24817]), .B(p_input[14817]), .Z(n11520) );
  AND U17280 ( .A(p_input[4817]), .B(p_input[34817]), .Z(n11519) );
  AND U17281 ( .A(n11521), .B(n11522), .Z(o[4816]) );
  AND U17282 ( .A(p_input[24816]), .B(p_input[14816]), .Z(n11522) );
  AND U17283 ( .A(p_input[4816]), .B(p_input[34816]), .Z(n11521) );
  AND U17284 ( .A(n11523), .B(n11524), .Z(o[4815]) );
  AND U17285 ( .A(p_input[24815]), .B(p_input[14815]), .Z(n11524) );
  AND U17286 ( .A(p_input[4815]), .B(p_input[34815]), .Z(n11523) );
  AND U17287 ( .A(n11525), .B(n11526), .Z(o[4814]) );
  AND U17288 ( .A(p_input[24814]), .B(p_input[14814]), .Z(n11526) );
  AND U17289 ( .A(p_input[4814]), .B(p_input[34814]), .Z(n11525) );
  AND U17290 ( .A(n11527), .B(n11528), .Z(o[4813]) );
  AND U17291 ( .A(p_input[24813]), .B(p_input[14813]), .Z(n11528) );
  AND U17292 ( .A(p_input[4813]), .B(p_input[34813]), .Z(n11527) );
  AND U17293 ( .A(n11529), .B(n11530), .Z(o[4812]) );
  AND U17294 ( .A(p_input[24812]), .B(p_input[14812]), .Z(n11530) );
  AND U17295 ( .A(p_input[4812]), .B(p_input[34812]), .Z(n11529) );
  AND U17296 ( .A(n11531), .B(n11532), .Z(o[4811]) );
  AND U17297 ( .A(p_input[24811]), .B(p_input[14811]), .Z(n11532) );
  AND U17298 ( .A(p_input[4811]), .B(p_input[34811]), .Z(n11531) );
  AND U17299 ( .A(n11533), .B(n11534), .Z(o[4810]) );
  AND U17300 ( .A(p_input[24810]), .B(p_input[14810]), .Z(n11534) );
  AND U17301 ( .A(p_input[4810]), .B(p_input[34810]), .Z(n11533) );
  AND U17302 ( .A(n11535), .B(n11536), .Z(o[480]) );
  AND U17303 ( .A(p_input[20480]), .B(p_input[10480]), .Z(n11536) );
  AND U17304 ( .A(p_input[480]), .B(p_input[30480]), .Z(n11535) );
  AND U17305 ( .A(n11537), .B(n11538), .Z(o[4809]) );
  AND U17306 ( .A(p_input[24809]), .B(p_input[14809]), .Z(n11538) );
  AND U17307 ( .A(p_input[4809]), .B(p_input[34809]), .Z(n11537) );
  AND U17308 ( .A(n11539), .B(n11540), .Z(o[4808]) );
  AND U17309 ( .A(p_input[24808]), .B(p_input[14808]), .Z(n11540) );
  AND U17310 ( .A(p_input[4808]), .B(p_input[34808]), .Z(n11539) );
  AND U17311 ( .A(n11541), .B(n11542), .Z(o[4807]) );
  AND U17312 ( .A(p_input[24807]), .B(p_input[14807]), .Z(n11542) );
  AND U17313 ( .A(p_input[4807]), .B(p_input[34807]), .Z(n11541) );
  AND U17314 ( .A(n11543), .B(n11544), .Z(o[4806]) );
  AND U17315 ( .A(p_input[24806]), .B(p_input[14806]), .Z(n11544) );
  AND U17316 ( .A(p_input[4806]), .B(p_input[34806]), .Z(n11543) );
  AND U17317 ( .A(n11545), .B(n11546), .Z(o[4805]) );
  AND U17318 ( .A(p_input[24805]), .B(p_input[14805]), .Z(n11546) );
  AND U17319 ( .A(p_input[4805]), .B(p_input[34805]), .Z(n11545) );
  AND U17320 ( .A(n11547), .B(n11548), .Z(o[4804]) );
  AND U17321 ( .A(p_input[24804]), .B(p_input[14804]), .Z(n11548) );
  AND U17322 ( .A(p_input[4804]), .B(p_input[34804]), .Z(n11547) );
  AND U17323 ( .A(n11549), .B(n11550), .Z(o[4803]) );
  AND U17324 ( .A(p_input[24803]), .B(p_input[14803]), .Z(n11550) );
  AND U17325 ( .A(p_input[4803]), .B(p_input[34803]), .Z(n11549) );
  AND U17326 ( .A(n11551), .B(n11552), .Z(o[4802]) );
  AND U17327 ( .A(p_input[24802]), .B(p_input[14802]), .Z(n11552) );
  AND U17328 ( .A(p_input[4802]), .B(p_input[34802]), .Z(n11551) );
  AND U17329 ( .A(n11553), .B(n11554), .Z(o[4801]) );
  AND U17330 ( .A(p_input[24801]), .B(p_input[14801]), .Z(n11554) );
  AND U17331 ( .A(p_input[4801]), .B(p_input[34801]), .Z(n11553) );
  AND U17332 ( .A(n11555), .B(n11556), .Z(o[4800]) );
  AND U17333 ( .A(p_input[24800]), .B(p_input[14800]), .Z(n11556) );
  AND U17334 ( .A(p_input[4800]), .B(p_input[34800]), .Z(n11555) );
  AND U17335 ( .A(n11557), .B(n11558), .Z(o[47]) );
  AND U17336 ( .A(p_input[20047]), .B(p_input[10047]), .Z(n11558) );
  AND U17337 ( .A(p_input[47]), .B(p_input[30047]), .Z(n11557) );
  AND U17338 ( .A(n11559), .B(n11560), .Z(o[479]) );
  AND U17339 ( .A(p_input[20479]), .B(p_input[10479]), .Z(n11560) );
  AND U17340 ( .A(p_input[479]), .B(p_input[30479]), .Z(n11559) );
  AND U17341 ( .A(n11561), .B(n11562), .Z(o[4799]) );
  AND U17342 ( .A(p_input[24799]), .B(p_input[14799]), .Z(n11562) );
  AND U17343 ( .A(p_input[4799]), .B(p_input[34799]), .Z(n11561) );
  AND U17344 ( .A(n11563), .B(n11564), .Z(o[4798]) );
  AND U17345 ( .A(p_input[24798]), .B(p_input[14798]), .Z(n11564) );
  AND U17346 ( .A(p_input[4798]), .B(p_input[34798]), .Z(n11563) );
  AND U17347 ( .A(n11565), .B(n11566), .Z(o[4797]) );
  AND U17348 ( .A(p_input[24797]), .B(p_input[14797]), .Z(n11566) );
  AND U17349 ( .A(p_input[4797]), .B(p_input[34797]), .Z(n11565) );
  AND U17350 ( .A(n11567), .B(n11568), .Z(o[4796]) );
  AND U17351 ( .A(p_input[24796]), .B(p_input[14796]), .Z(n11568) );
  AND U17352 ( .A(p_input[4796]), .B(p_input[34796]), .Z(n11567) );
  AND U17353 ( .A(n11569), .B(n11570), .Z(o[4795]) );
  AND U17354 ( .A(p_input[24795]), .B(p_input[14795]), .Z(n11570) );
  AND U17355 ( .A(p_input[4795]), .B(p_input[34795]), .Z(n11569) );
  AND U17356 ( .A(n11571), .B(n11572), .Z(o[4794]) );
  AND U17357 ( .A(p_input[24794]), .B(p_input[14794]), .Z(n11572) );
  AND U17358 ( .A(p_input[4794]), .B(p_input[34794]), .Z(n11571) );
  AND U17359 ( .A(n11573), .B(n11574), .Z(o[4793]) );
  AND U17360 ( .A(p_input[24793]), .B(p_input[14793]), .Z(n11574) );
  AND U17361 ( .A(p_input[4793]), .B(p_input[34793]), .Z(n11573) );
  AND U17362 ( .A(n11575), .B(n11576), .Z(o[4792]) );
  AND U17363 ( .A(p_input[24792]), .B(p_input[14792]), .Z(n11576) );
  AND U17364 ( .A(p_input[4792]), .B(p_input[34792]), .Z(n11575) );
  AND U17365 ( .A(n11577), .B(n11578), .Z(o[4791]) );
  AND U17366 ( .A(p_input[24791]), .B(p_input[14791]), .Z(n11578) );
  AND U17367 ( .A(p_input[4791]), .B(p_input[34791]), .Z(n11577) );
  AND U17368 ( .A(n11579), .B(n11580), .Z(o[4790]) );
  AND U17369 ( .A(p_input[24790]), .B(p_input[14790]), .Z(n11580) );
  AND U17370 ( .A(p_input[4790]), .B(p_input[34790]), .Z(n11579) );
  AND U17371 ( .A(n11581), .B(n11582), .Z(o[478]) );
  AND U17372 ( .A(p_input[20478]), .B(p_input[10478]), .Z(n11582) );
  AND U17373 ( .A(p_input[478]), .B(p_input[30478]), .Z(n11581) );
  AND U17374 ( .A(n11583), .B(n11584), .Z(o[4789]) );
  AND U17375 ( .A(p_input[24789]), .B(p_input[14789]), .Z(n11584) );
  AND U17376 ( .A(p_input[4789]), .B(p_input[34789]), .Z(n11583) );
  AND U17377 ( .A(n11585), .B(n11586), .Z(o[4788]) );
  AND U17378 ( .A(p_input[24788]), .B(p_input[14788]), .Z(n11586) );
  AND U17379 ( .A(p_input[4788]), .B(p_input[34788]), .Z(n11585) );
  AND U17380 ( .A(n11587), .B(n11588), .Z(o[4787]) );
  AND U17381 ( .A(p_input[24787]), .B(p_input[14787]), .Z(n11588) );
  AND U17382 ( .A(p_input[4787]), .B(p_input[34787]), .Z(n11587) );
  AND U17383 ( .A(n11589), .B(n11590), .Z(o[4786]) );
  AND U17384 ( .A(p_input[24786]), .B(p_input[14786]), .Z(n11590) );
  AND U17385 ( .A(p_input[4786]), .B(p_input[34786]), .Z(n11589) );
  AND U17386 ( .A(n11591), .B(n11592), .Z(o[4785]) );
  AND U17387 ( .A(p_input[24785]), .B(p_input[14785]), .Z(n11592) );
  AND U17388 ( .A(p_input[4785]), .B(p_input[34785]), .Z(n11591) );
  AND U17389 ( .A(n11593), .B(n11594), .Z(o[4784]) );
  AND U17390 ( .A(p_input[24784]), .B(p_input[14784]), .Z(n11594) );
  AND U17391 ( .A(p_input[4784]), .B(p_input[34784]), .Z(n11593) );
  AND U17392 ( .A(n11595), .B(n11596), .Z(o[4783]) );
  AND U17393 ( .A(p_input[24783]), .B(p_input[14783]), .Z(n11596) );
  AND U17394 ( .A(p_input[4783]), .B(p_input[34783]), .Z(n11595) );
  AND U17395 ( .A(n11597), .B(n11598), .Z(o[4782]) );
  AND U17396 ( .A(p_input[24782]), .B(p_input[14782]), .Z(n11598) );
  AND U17397 ( .A(p_input[4782]), .B(p_input[34782]), .Z(n11597) );
  AND U17398 ( .A(n11599), .B(n11600), .Z(o[4781]) );
  AND U17399 ( .A(p_input[24781]), .B(p_input[14781]), .Z(n11600) );
  AND U17400 ( .A(p_input[4781]), .B(p_input[34781]), .Z(n11599) );
  AND U17401 ( .A(n11601), .B(n11602), .Z(o[4780]) );
  AND U17402 ( .A(p_input[24780]), .B(p_input[14780]), .Z(n11602) );
  AND U17403 ( .A(p_input[4780]), .B(p_input[34780]), .Z(n11601) );
  AND U17404 ( .A(n11603), .B(n11604), .Z(o[477]) );
  AND U17405 ( .A(p_input[20477]), .B(p_input[10477]), .Z(n11604) );
  AND U17406 ( .A(p_input[477]), .B(p_input[30477]), .Z(n11603) );
  AND U17407 ( .A(n11605), .B(n11606), .Z(o[4779]) );
  AND U17408 ( .A(p_input[24779]), .B(p_input[14779]), .Z(n11606) );
  AND U17409 ( .A(p_input[4779]), .B(p_input[34779]), .Z(n11605) );
  AND U17410 ( .A(n11607), .B(n11608), .Z(o[4778]) );
  AND U17411 ( .A(p_input[24778]), .B(p_input[14778]), .Z(n11608) );
  AND U17412 ( .A(p_input[4778]), .B(p_input[34778]), .Z(n11607) );
  AND U17413 ( .A(n11609), .B(n11610), .Z(o[4777]) );
  AND U17414 ( .A(p_input[24777]), .B(p_input[14777]), .Z(n11610) );
  AND U17415 ( .A(p_input[4777]), .B(p_input[34777]), .Z(n11609) );
  AND U17416 ( .A(n11611), .B(n11612), .Z(o[4776]) );
  AND U17417 ( .A(p_input[24776]), .B(p_input[14776]), .Z(n11612) );
  AND U17418 ( .A(p_input[4776]), .B(p_input[34776]), .Z(n11611) );
  AND U17419 ( .A(n11613), .B(n11614), .Z(o[4775]) );
  AND U17420 ( .A(p_input[24775]), .B(p_input[14775]), .Z(n11614) );
  AND U17421 ( .A(p_input[4775]), .B(p_input[34775]), .Z(n11613) );
  AND U17422 ( .A(n11615), .B(n11616), .Z(o[4774]) );
  AND U17423 ( .A(p_input[24774]), .B(p_input[14774]), .Z(n11616) );
  AND U17424 ( .A(p_input[4774]), .B(p_input[34774]), .Z(n11615) );
  AND U17425 ( .A(n11617), .B(n11618), .Z(o[4773]) );
  AND U17426 ( .A(p_input[24773]), .B(p_input[14773]), .Z(n11618) );
  AND U17427 ( .A(p_input[4773]), .B(p_input[34773]), .Z(n11617) );
  AND U17428 ( .A(n11619), .B(n11620), .Z(o[4772]) );
  AND U17429 ( .A(p_input[24772]), .B(p_input[14772]), .Z(n11620) );
  AND U17430 ( .A(p_input[4772]), .B(p_input[34772]), .Z(n11619) );
  AND U17431 ( .A(n11621), .B(n11622), .Z(o[4771]) );
  AND U17432 ( .A(p_input[24771]), .B(p_input[14771]), .Z(n11622) );
  AND U17433 ( .A(p_input[4771]), .B(p_input[34771]), .Z(n11621) );
  AND U17434 ( .A(n11623), .B(n11624), .Z(o[4770]) );
  AND U17435 ( .A(p_input[24770]), .B(p_input[14770]), .Z(n11624) );
  AND U17436 ( .A(p_input[4770]), .B(p_input[34770]), .Z(n11623) );
  AND U17437 ( .A(n11625), .B(n11626), .Z(o[476]) );
  AND U17438 ( .A(p_input[20476]), .B(p_input[10476]), .Z(n11626) );
  AND U17439 ( .A(p_input[476]), .B(p_input[30476]), .Z(n11625) );
  AND U17440 ( .A(n11627), .B(n11628), .Z(o[4769]) );
  AND U17441 ( .A(p_input[24769]), .B(p_input[14769]), .Z(n11628) );
  AND U17442 ( .A(p_input[4769]), .B(p_input[34769]), .Z(n11627) );
  AND U17443 ( .A(n11629), .B(n11630), .Z(o[4768]) );
  AND U17444 ( .A(p_input[24768]), .B(p_input[14768]), .Z(n11630) );
  AND U17445 ( .A(p_input[4768]), .B(p_input[34768]), .Z(n11629) );
  AND U17446 ( .A(n11631), .B(n11632), .Z(o[4767]) );
  AND U17447 ( .A(p_input[24767]), .B(p_input[14767]), .Z(n11632) );
  AND U17448 ( .A(p_input[4767]), .B(p_input[34767]), .Z(n11631) );
  AND U17449 ( .A(n11633), .B(n11634), .Z(o[4766]) );
  AND U17450 ( .A(p_input[24766]), .B(p_input[14766]), .Z(n11634) );
  AND U17451 ( .A(p_input[4766]), .B(p_input[34766]), .Z(n11633) );
  AND U17452 ( .A(n11635), .B(n11636), .Z(o[4765]) );
  AND U17453 ( .A(p_input[24765]), .B(p_input[14765]), .Z(n11636) );
  AND U17454 ( .A(p_input[4765]), .B(p_input[34765]), .Z(n11635) );
  AND U17455 ( .A(n11637), .B(n11638), .Z(o[4764]) );
  AND U17456 ( .A(p_input[24764]), .B(p_input[14764]), .Z(n11638) );
  AND U17457 ( .A(p_input[4764]), .B(p_input[34764]), .Z(n11637) );
  AND U17458 ( .A(n11639), .B(n11640), .Z(o[4763]) );
  AND U17459 ( .A(p_input[24763]), .B(p_input[14763]), .Z(n11640) );
  AND U17460 ( .A(p_input[4763]), .B(p_input[34763]), .Z(n11639) );
  AND U17461 ( .A(n11641), .B(n11642), .Z(o[4762]) );
  AND U17462 ( .A(p_input[24762]), .B(p_input[14762]), .Z(n11642) );
  AND U17463 ( .A(p_input[4762]), .B(p_input[34762]), .Z(n11641) );
  AND U17464 ( .A(n11643), .B(n11644), .Z(o[4761]) );
  AND U17465 ( .A(p_input[24761]), .B(p_input[14761]), .Z(n11644) );
  AND U17466 ( .A(p_input[4761]), .B(p_input[34761]), .Z(n11643) );
  AND U17467 ( .A(n11645), .B(n11646), .Z(o[4760]) );
  AND U17468 ( .A(p_input[24760]), .B(p_input[14760]), .Z(n11646) );
  AND U17469 ( .A(p_input[4760]), .B(p_input[34760]), .Z(n11645) );
  AND U17470 ( .A(n11647), .B(n11648), .Z(o[475]) );
  AND U17471 ( .A(p_input[20475]), .B(p_input[10475]), .Z(n11648) );
  AND U17472 ( .A(p_input[475]), .B(p_input[30475]), .Z(n11647) );
  AND U17473 ( .A(n11649), .B(n11650), .Z(o[4759]) );
  AND U17474 ( .A(p_input[24759]), .B(p_input[14759]), .Z(n11650) );
  AND U17475 ( .A(p_input[4759]), .B(p_input[34759]), .Z(n11649) );
  AND U17476 ( .A(n11651), .B(n11652), .Z(o[4758]) );
  AND U17477 ( .A(p_input[24758]), .B(p_input[14758]), .Z(n11652) );
  AND U17478 ( .A(p_input[4758]), .B(p_input[34758]), .Z(n11651) );
  AND U17479 ( .A(n11653), .B(n11654), .Z(o[4757]) );
  AND U17480 ( .A(p_input[24757]), .B(p_input[14757]), .Z(n11654) );
  AND U17481 ( .A(p_input[4757]), .B(p_input[34757]), .Z(n11653) );
  AND U17482 ( .A(n11655), .B(n11656), .Z(o[4756]) );
  AND U17483 ( .A(p_input[24756]), .B(p_input[14756]), .Z(n11656) );
  AND U17484 ( .A(p_input[4756]), .B(p_input[34756]), .Z(n11655) );
  AND U17485 ( .A(n11657), .B(n11658), .Z(o[4755]) );
  AND U17486 ( .A(p_input[24755]), .B(p_input[14755]), .Z(n11658) );
  AND U17487 ( .A(p_input[4755]), .B(p_input[34755]), .Z(n11657) );
  AND U17488 ( .A(n11659), .B(n11660), .Z(o[4754]) );
  AND U17489 ( .A(p_input[24754]), .B(p_input[14754]), .Z(n11660) );
  AND U17490 ( .A(p_input[4754]), .B(p_input[34754]), .Z(n11659) );
  AND U17491 ( .A(n11661), .B(n11662), .Z(o[4753]) );
  AND U17492 ( .A(p_input[24753]), .B(p_input[14753]), .Z(n11662) );
  AND U17493 ( .A(p_input[4753]), .B(p_input[34753]), .Z(n11661) );
  AND U17494 ( .A(n11663), .B(n11664), .Z(o[4752]) );
  AND U17495 ( .A(p_input[24752]), .B(p_input[14752]), .Z(n11664) );
  AND U17496 ( .A(p_input[4752]), .B(p_input[34752]), .Z(n11663) );
  AND U17497 ( .A(n11665), .B(n11666), .Z(o[4751]) );
  AND U17498 ( .A(p_input[24751]), .B(p_input[14751]), .Z(n11666) );
  AND U17499 ( .A(p_input[4751]), .B(p_input[34751]), .Z(n11665) );
  AND U17500 ( .A(n11667), .B(n11668), .Z(o[4750]) );
  AND U17501 ( .A(p_input[24750]), .B(p_input[14750]), .Z(n11668) );
  AND U17502 ( .A(p_input[4750]), .B(p_input[34750]), .Z(n11667) );
  AND U17503 ( .A(n11669), .B(n11670), .Z(o[474]) );
  AND U17504 ( .A(p_input[20474]), .B(p_input[10474]), .Z(n11670) );
  AND U17505 ( .A(p_input[474]), .B(p_input[30474]), .Z(n11669) );
  AND U17506 ( .A(n11671), .B(n11672), .Z(o[4749]) );
  AND U17507 ( .A(p_input[24749]), .B(p_input[14749]), .Z(n11672) );
  AND U17508 ( .A(p_input[4749]), .B(p_input[34749]), .Z(n11671) );
  AND U17509 ( .A(n11673), .B(n11674), .Z(o[4748]) );
  AND U17510 ( .A(p_input[24748]), .B(p_input[14748]), .Z(n11674) );
  AND U17511 ( .A(p_input[4748]), .B(p_input[34748]), .Z(n11673) );
  AND U17512 ( .A(n11675), .B(n11676), .Z(o[4747]) );
  AND U17513 ( .A(p_input[24747]), .B(p_input[14747]), .Z(n11676) );
  AND U17514 ( .A(p_input[4747]), .B(p_input[34747]), .Z(n11675) );
  AND U17515 ( .A(n11677), .B(n11678), .Z(o[4746]) );
  AND U17516 ( .A(p_input[24746]), .B(p_input[14746]), .Z(n11678) );
  AND U17517 ( .A(p_input[4746]), .B(p_input[34746]), .Z(n11677) );
  AND U17518 ( .A(n11679), .B(n11680), .Z(o[4745]) );
  AND U17519 ( .A(p_input[24745]), .B(p_input[14745]), .Z(n11680) );
  AND U17520 ( .A(p_input[4745]), .B(p_input[34745]), .Z(n11679) );
  AND U17521 ( .A(n11681), .B(n11682), .Z(o[4744]) );
  AND U17522 ( .A(p_input[24744]), .B(p_input[14744]), .Z(n11682) );
  AND U17523 ( .A(p_input[4744]), .B(p_input[34744]), .Z(n11681) );
  AND U17524 ( .A(n11683), .B(n11684), .Z(o[4743]) );
  AND U17525 ( .A(p_input[24743]), .B(p_input[14743]), .Z(n11684) );
  AND U17526 ( .A(p_input[4743]), .B(p_input[34743]), .Z(n11683) );
  AND U17527 ( .A(n11685), .B(n11686), .Z(o[4742]) );
  AND U17528 ( .A(p_input[24742]), .B(p_input[14742]), .Z(n11686) );
  AND U17529 ( .A(p_input[4742]), .B(p_input[34742]), .Z(n11685) );
  AND U17530 ( .A(n11687), .B(n11688), .Z(o[4741]) );
  AND U17531 ( .A(p_input[24741]), .B(p_input[14741]), .Z(n11688) );
  AND U17532 ( .A(p_input[4741]), .B(p_input[34741]), .Z(n11687) );
  AND U17533 ( .A(n11689), .B(n11690), .Z(o[4740]) );
  AND U17534 ( .A(p_input[24740]), .B(p_input[14740]), .Z(n11690) );
  AND U17535 ( .A(p_input[4740]), .B(p_input[34740]), .Z(n11689) );
  AND U17536 ( .A(n11691), .B(n11692), .Z(o[473]) );
  AND U17537 ( .A(p_input[20473]), .B(p_input[10473]), .Z(n11692) );
  AND U17538 ( .A(p_input[473]), .B(p_input[30473]), .Z(n11691) );
  AND U17539 ( .A(n11693), .B(n11694), .Z(o[4739]) );
  AND U17540 ( .A(p_input[24739]), .B(p_input[14739]), .Z(n11694) );
  AND U17541 ( .A(p_input[4739]), .B(p_input[34739]), .Z(n11693) );
  AND U17542 ( .A(n11695), .B(n11696), .Z(o[4738]) );
  AND U17543 ( .A(p_input[24738]), .B(p_input[14738]), .Z(n11696) );
  AND U17544 ( .A(p_input[4738]), .B(p_input[34738]), .Z(n11695) );
  AND U17545 ( .A(n11697), .B(n11698), .Z(o[4737]) );
  AND U17546 ( .A(p_input[24737]), .B(p_input[14737]), .Z(n11698) );
  AND U17547 ( .A(p_input[4737]), .B(p_input[34737]), .Z(n11697) );
  AND U17548 ( .A(n11699), .B(n11700), .Z(o[4736]) );
  AND U17549 ( .A(p_input[24736]), .B(p_input[14736]), .Z(n11700) );
  AND U17550 ( .A(p_input[4736]), .B(p_input[34736]), .Z(n11699) );
  AND U17551 ( .A(n11701), .B(n11702), .Z(o[4735]) );
  AND U17552 ( .A(p_input[24735]), .B(p_input[14735]), .Z(n11702) );
  AND U17553 ( .A(p_input[4735]), .B(p_input[34735]), .Z(n11701) );
  AND U17554 ( .A(n11703), .B(n11704), .Z(o[4734]) );
  AND U17555 ( .A(p_input[24734]), .B(p_input[14734]), .Z(n11704) );
  AND U17556 ( .A(p_input[4734]), .B(p_input[34734]), .Z(n11703) );
  AND U17557 ( .A(n11705), .B(n11706), .Z(o[4733]) );
  AND U17558 ( .A(p_input[24733]), .B(p_input[14733]), .Z(n11706) );
  AND U17559 ( .A(p_input[4733]), .B(p_input[34733]), .Z(n11705) );
  AND U17560 ( .A(n11707), .B(n11708), .Z(o[4732]) );
  AND U17561 ( .A(p_input[24732]), .B(p_input[14732]), .Z(n11708) );
  AND U17562 ( .A(p_input[4732]), .B(p_input[34732]), .Z(n11707) );
  AND U17563 ( .A(n11709), .B(n11710), .Z(o[4731]) );
  AND U17564 ( .A(p_input[24731]), .B(p_input[14731]), .Z(n11710) );
  AND U17565 ( .A(p_input[4731]), .B(p_input[34731]), .Z(n11709) );
  AND U17566 ( .A(n11711), .B(n11712), .Z(o[4730]) );
  AND U17567 ( .A(p_input[24730]), .B(p_input[14730]), .Z(n11712) );
  AND U17568 ( .A(p_input[4730]), .B(p_input[34730]), .Z(n11711) );
  AND U17569 ( .A(n11713), .B(n11714), .Z(o[472]) );
  AND U17570 ( .A(p_input[20472]), .B(p_input[10472]), .Z(n11714) );
  AND U17571 ( .A(p_input[472]), .B(p_input[30472]), .Z(n11713) );
  AND U17572 ( .A(n11715), .B(n11716), .Z(o[4729]) );
  AND U17573 ( .A(p_input[24729]), .B(p_input[14729]), .Z(n11716) );
  AND U17574 ( .A(p_input[4729]), .B(p_input[34729]), .Z(n11715) );
  AND U17575 ( .A(n11717), .B(n11718), .Z(o[4728]) );
  AND U17576 ( .A(p_input[24728]), .B(p_input[14728]), .Z(n11718) );
  AND U17577 ( .A(p_input[4728]), .B(p_input[34728]), .Z(n11717) );
  AND U17578 ( .A(n11719), .B(n11720), .Z(o[4727]) );
  AND U17579 ( .A(p_input[24727]), .B(p_input[14727]), .Z(n11720) );
  AND U17580 ( .A(p_input[4727]), .B(p_input[34727]), .Z(n11719) );
  AND U17581 ( .A(n11721), .B(n11722), .Z(o[4726]) );
  AND U17582 ( .A(p_input[24726]), .B(p_input[14726]), .Z(n11722) );
  AND U17583 ( .A(p_input[4726]), .B(p_input[34726]), .Z(n11721) );
  AND U17584 ( .A(n11723), .B(n11724), .Z(o[4725]) );
  AND U17585 ( .A(p_input[24725]), .B(p_input[14725]), .Z(n11724) );
  AND U17586 ( .A(p_input[4725]), .B(p_input[34725]), .Z(n11723) );
  AND U17587 ( .A(n11725), .B(n11726), .Z(o[4724]) );
  AND U17588 ( .A(p_input[24724]), .B(p_input[14724]), .Z(n11726) );
  AND U17589 ( .A(p_input[4724]), .B(p_input[34724]), .Z(n11725) );
  AND U17590 ( .A(n11727), .B(n11728), .Z(o[4723]) );
  AND U17591 ( .A(p_input[24723]), .B(p_input[14723]), .Z(n11728) );
  AND U17592 ( .A(p_input[4723]), .B(p_input[34723]), .Z(n11727) );
  AND U17593 ( .A(n11729), .B(n11730), .Z(o[4722]) );
  AND U17594 ( .A(p_input[24722]), .B(p_input[14722]), .Z(n11730) );
  AND U17595 ( .A(p_input[4722]), .B(p_input[34722]), .Z(n11729) );
  AND U17596 ( .A(n11731), .B(n11732), .Z(o[4721]) );
  AND U17597 ( .A(p_input[24721]), .B(p_input[14721]), .Z(n11732) );
  AND U17598 ( .A(p_input[4721]), .B(p_input[34721]), .Z(n11731) );
  AND U17599 ( .A(n11733), .B(n11734), .Z(o[4720]) );
  AND U17600 ( .A(p_input[24720]), .B(p_input[14720]), .Z(n11734) );
  AND U17601 ( .A(p_input[4720]), .B(p_input[34720]), .Z(n11733) );
  AND U17602 ( .A(n11735), .B(n11736), .Z(o[471]) );
  AND U17603 ( .A(p_input[20471]), .B(p_input[10471]), .Z(n11736) );
  AND U17604 ( .A(p_input[471]), .B(p_input[30471]), .Z(n11735) );
  AND U17605 ( .A(n11737), .B(n11738), .Z(o[4719]) );
  AND U17606 ( .A(p_input[24719]), .B(p_input[14719]), .Z(n11738) );
  AND U17607 ( .A(p_input[4719]), .B(p_input[34719]), .Z(n11737) );
  AND U17608 ( .A(n11739), .B(n11740), .Z(o[4718]) );
  AND U17609 ( .A(p_input[24718]), .B(p_input[14718]), .Z(n11740) );
  AND U17610 ( .A(p_input[4718]), .B(p_input[34718]), .Z(n11739) );
  AND U17611 ( .A(n11741), .B(n11742), .Z(o[4717]) );
  AND U17612 ( .A(p_input[24717]), .B(p_input[14717]), .Z(n11742) );
  AND U17613 ( .A(p_input[4717]), .B(p_input[34717]), .Z(n11741) );
  AND U17614 ( .A(n11743), .B(n11744), .Z(o[4716]) );
  AND U17615 ( .A(p_input[24716]), .B(p_input[14716]), .Z(n11744) );
  AND U17616 ( .A(p_input[4716]), .B(p_input[34716]), .Z(n11743) );
  AND U17617 ( .A(n11745), .B(n11746), .Z(o[4715]) );
  AND U17618 ( .A(p_input[24715]), .B(p_input[14715]), .Z(n11746) );
  AND U17619 ( .A(p_input[4715]), .B(p_input[34715]), .Z(n11745) );
  AND U17620 ( .A(n11747), .B(n11748), .Z(o[4714]) );
  AND U17621 ( .A(p_input[24714]), .B(p_input[14714]), .Z(n11748) );
  AND U17622 ( .A(p_input[4714]), .B(p_input[34714]), .Z(n11747) );
  AND U17623 ( .A(n11749), .B(n11750), .Z(o[4713]) );
  AND U17624 ( .A(p_input[24713]), .B(p_input[14713]), .Z(n11750) );
  AND U17625 ( .A(p_input[4713]), .B(p_input[34713]), .Z(n11749) );
  AND U17626 ( .A(n11751), .B(n11752), .Z(o[4712]) );
  AND U17627 ( .A(p_input[24712]), .B(p_input[14712]), .Z(n11752) );
  AND U17628 ( .A(p_input[4712]), .B(p_input[34712]), .Z(n11751) );
  AND U17629 ( .A(n11753), .B(n11754), .Z(o[4711]) );
  AND U17630 ( .A(p_input[24711]), .B(p_input[14711]), .Z(n11754) );
  AND U17631 ( .A(p_input[4711]), .B(p_input[34711]), .Z(n11753) );
  AND U17632 ( .A(n11755), .B(n11756), .Z(o[4710]) );
  AND U17633 ( .A(p_input[24710]), .B(p_input[14710]), .Z(n11756) );
  AND U17634 ( .A(p_input[4710]), .B(p_input[34710]), .Z(n11755) );
  AND U17635 ( .A(n11757), .B(n11758), .Z(o[470]) );
  AND U17636 ( .A(p_input[20470]), .B(p_input[10470]), .Z(n11758) );
  AND U17637 ( .A(p_input[470]), .B(p_input[30470]), .Z(n11757) );
  AND U17638 ( .A(n11759), .B(n11760), .Z(o[4709]) );
  AND U17639 ( .A(p_input[24709]), .B(p_input[14709]), .Z(n11760) );
  AND U17640 ( .A(p_input[4709]), .B(p_input[34709]), .Z(n11759) );
  AND U17641 ( .A(n11761), .B(n11762), .Z(o[4708]) );
  AND U17642 ( .A(p_input[24708]), .B(p_input[14708]), .Z(n11762) );
  AND U17643 ( .A(p_input[4708]), .B(p_input[34708]), .Z(n11761) );
  AND U17644 ( .A(n11763), .B(n11764), .Z(o[4707]) );
  AND U17645 ( .A(p_input[24707]), .B(p_input[14707]), .Z(n11764) );
  AND U17646 ( .A(p_input[4707]), .B(p_input[34707]), .Z(n11763) );
  AND U17647 ( .A(n11765), .B(n11766), .Z(o[4706]) );
  AND U17648 ( .A(p_input[24706]), .B(p_input[14706]), .Z(n11766) );
  AND U17649 ( .A(p_input[4706]), .B(p_input[34706]), .Z(n11765) );
  AND U17650 ( .A(n11767), .B(n11768), .Z(o[4705]) );
  AND U17651 ( .A(p_input[24705]), .B(p_input[14705]), .Z(n11768) );
  AND U17652 ( .A(p_input[4705]), .B(p_input[34705]), .Z(n11767) );
  AND U17653 ( .A(n11769), .B(n11770), .Z(o[4704]) );
  AND U17654 ( .A(p_input[24704]), .B(p_input[14704]), .Z(n11770) );
  AND U17655 ( .A(p_input[4704]), .B(p_input[34704]), .Z(n11769) );
  AND U17656 ( .A(n11771), .B(n11772), .Z(o[4703]) );
  AND U17657 ( .A(p_input[24703]), .B(p_input[14703]), .Z(n11772) );
  AND U17658 ( .A(p_input[4703]), .B(p_input[34703]), .Z(n11771) );
  AND U17659 ( .A(n11773), .B(n11774), .Z(o[4702]) );
  AND U17660 ( .A(p_input[24702]), .B(p_input[14702]), .Z(n11774) );
  AND U17661 ( .A(p_input[4702]), .B(p_input[34702]), .Z(n11773) );
  AND U17662 ( .A(n11775), .B(n11776), .Z(o[4701]) );
  AND U17663 ( .A(p_input[24701]), .B(p_input[14701]), .Z(n11776) );
  AND U17664 ( .A(p_input[4701]), .B(p_input[34701]), .Z(n11775) );
  AND U17665 ( .A(n11777), .B(n11778), .Z(o[4700]) );
  AND U17666 ( .A(p_input[24700]), .B(p_input[14700]), .Z(n11778) );
  AND U17667 ( .A(p_input[4700]), .B(p_input[34700]), .Z(n11777) );
  AND U17668 ( .A(n11779), .B(n11780), .Z(o[46]) );
  AND U17669 ( .A(p_input[20046]), .B(p_input[10046]), .Z(n11780) );
  AND U17670 ( .A(p_input[46]), .B(p_input[30046]), .Z(n11779) );
  AND U17671 ( .A(n11781), .B(n11782), .Z(o[469]) );
  AND U17672 ( .A(p_input[20469]), .B(p_input[10469]), .Z(n11782) );
  AND U17673 ( .A(p_input[469]), .B(p_input[30469]), .Z(n11781) );
  AND U17674 ( .A(n11783), .B(n11784), .Z(o[4699]) );
  AND U17675 ( .A(p_input[24699]), .B(p_input[14699]), .Z(n11784) );
  AND U17676 ( .A(p_input[4699]), .B(p_input[34699]), .Z(n11783) );
  AND U17677 ( .A(n11785), .B(n11786), .Z(o[4698]) );
  AND U17678 ( .A(p_input[24698]), .B(p_input[14698]), .Z(n11786) );
  AND U17679 ( .A(p_input[4698]), .B(p_input[34698]), .Z(n11785) );
  AND U17680 ( .A(n11787), .B(n11788), .Z(o[4697]) );
  AND U17681 ( .A(p_input[24697]), .B(p_input[14697]), .Z(n11788) );
  AND U17682 ( .A(p_input[4697]), .B(p_input[34697]), .Z(n11787) );
  AND U17683 ( .A(n11789), .B(n11790), .Z(o[4696]) );
  AND U17684 ( .A(p_input[24696]), .B(p_input[14696]), .Z(n11790) );
  AND U17685 ( .A(p_input[4696]), .B(p_input[34696]), .Z(n11789) );
  AND U17686 ( .A(n11791), .B(n11792), .Z(o[4695]) );
  AND U17687 ( .A(p_input[24695]), .B(p_input[14695]), .Z(n11792) );
  AND U17688 ( .A(p_input[4695]), .B(p_input[34695]), .Z(n11791) );
  AND U17689 ( .A(n11793), .B(n11794), .Z(o[4694]) );
  AND U17690 ( .A(p_input[24694]), .B(p_input[14694]), .Z(n11794) );
  AND U17691 ( .A(p_input[4694]), .B(p_input[34694]), .Z(n11793) );
  AND U17692 ( .A(n11795), .B(n11796), .Z(o[4693]) );
  AND U17693 ( .A(p_input[24693]), .B(p_input[14693]), .Z(n11796) );
  AND U17694 ( .A(p_input[4693]), .B(p_input[34693]), .Z(n11795) );
  AND U17695 ( .A(n11797), .B(n11798), .Z(o[4692]) );
  AND U17696 ( .A(p_input[24692]), .B(p_input[14692]), .Z(n11798) );
  AND U17697 ( .A(p_input[4692]), .B(p_input[34692]), .Z(n11797) );
  AND U17698 ( .A(n11799), .B(n11800), .Z(o[4691]) );
  AND U17699 ( .A(p_input[24691]), .B(p_input[14691]), .Z(n11800) );
  AND U17700 ( .A(p_input[4691]), .B(p_input[34691]), .Z(n11799) );
  AND U17701 ( .A(n11801), .B(n11802), .Z(o[4690]) );
  AND U17702 ( .A(p_input[24690]), .B(p_input[14690]), .Z(n11802) );
  AND U17703 ( .A(p_input[4690]), .B(p_input[34690]), .Z(n11801) );
  AND U17704 ( .A(n11803), .B(n11804), .Z(o[468]) );
  AND U17705 ( .A(p_input[20468]), .B(p_input[10468]), .Z(n11804) );
  AND U17706 ( .A(p_input[468]), .B(p_input[30468]), .Z(n11803) );
  AND U17707 ( .A(n11805), .B(n11806), .Z(o[4689]) );
  AND U17708 ( .A(p_input[24689]), .B(p_input[14689]), .Z(n11806) );
  AND U17709 ( .A(p_input[4689]), .B(p_input[34689]), .Z(n11805) );
  AND U17710 ( .A(n11807), .B(n11808), .Z(o[4688]) );
  AND U17711 ( .A(p_input[24688]), .B(p_input[14688]), .Z(n11808) );
  AND U17712 ( .A(p_input[4688]), .B(p_input[34688]), .Z(n11807) );
  AND U17713 ( .A(n11809), .B(n11810), .Z(o[4687]) );
  AND U17714 ( .A(p_input[24687]), .B(p_input[14687]), .Z(n11810) );
  AND U17715 ( .A(p_input[4687]), .B(p_input[34687]), .Z(n11809) );
  AND U17716 ( .A(n11811), .B(n11812), .Z(o[4686]) );
  AND U17717 ( .A(p_input[24686]), .B(p_input[14686]), .Z(n11812) );
  AND U17718 ( .A(p_input[4686]), .B(p_input[34686]), .Z(n11811) );
  AND U17719 ( .A(n11813), .B(n11814), .Z(o[4685]) );
  AND U17720 ( .A(p_input[24685]), .B(p_input[14685]), .Z(n11814) );
  AND U17721 ( .A(p_input[4685]), .B(p_input[34685]), .Z(n11813) );
  AND U17722 ( .A(n11815), .B(n11816), .Z(o[4684]) );
  AND U17723 ( .A(p_input[24684]), .B(p_input[14684]), .Z(n11816) );
  AND U17724 ( .A(p_input[4684]), .B(p_input[34684]), .Z(n11815) );
  AND U17725 ( .A(n11817), .B(n11818), .Z(o[4683]) );
  AND U17726 ( .A(p_input[24683]), .B(p_input[14683]), .Z(n11818) );
  AND U17727 ( .A(p_input[4683]), .B(p_input[34683]), .Z(n11817) );
  AND U17728 ( .A(n11819), .B(n11820), .Z(o[4682]) );
  AND U17729 ( .A(p_input[24682]), .B(p_input[14682]), .Z(n11820) );
  AND U17730 ( .A(p_input[4682]), .B(p_input[34682]), .Z(n11819) );
  AND U17731 ( .A(n11821), .B(n11822), .Z(o[4681]) );
  AND U17732 ( .A(p_input[24681]), .B(p_input[14681]), .Z(n11822) );
  AND U17733 ( .A(p_input[4681]), .B(p_input[34681]), .Z(n11821) );
  AND U17734 ( .A(n11823), .B(n11824), .Z(o[4680]) );
  AND U17735 ( .A(p_input[24680]), .B(p_input[14680]), .Z(n11824) );
  AND U17736 ( .A(p_input[4680]), .B(p_input[34680]), .Z(n11823) );
  AND U17737 ( .A(n11825), .B(n11826), .Z(o[467]) );
  AND U17738 ( .A(p_input[20467]), .B(p_input[10467]), .Z(n11826) );
  AND U17739 ( .A(p_input[467]), .B(p_input[30467]), .Z(n11825) );
  AND U17740 ( .A(n11827), .B(n11828), .Z(o[4679]) );
  AND U17741 ( .A(p_input[24679]), .B(p_input[14679]), .Z(n11828) );
  AND U17742 ( .A(p_input[4679]), .B(p_input[34679]), .Z(n11827) );
  AND U17743 ( .A(n11829), .B(n11830), .Z(o[4678]) );
  AND U17744 ( .A(p_input[24678]), .B(p_input[14678]), .Z(n11830) );
  AND U17745 ( .A(p_input[4678]), .B(p_input[34678]), .Z(n11829) );
  AND U17746 ( .A(n11831), .B(n11832), .Z(o[4677]) );
  AND U17747 ( .A(p_input[24677]), .B(p_input[14677]), .Z(n11832) );
  AND U17748 ( .A(p_input[4677]), .B(p_input[34677]), .Z(n11831) );
  AND U17749 ( .A(n11833), .B(n11834), .Z(o[4676]) );
  AND U17750 ( .A(p_input[24676]), .B(p_input[14676]), .Z(n11834) );
  AND U17751 ( .A(p_input[4676]), .B(p_input[34676]), .Z(n11833) );
  AND U17752 ( .A(n11835), .B(n11836), .Z(o[4675]) );
  AND U17753 ( .A(p_input[24675]), .B(p_input[14675]), .Z(n11836) );
  AND U17754 ( .A(p_input[4675]), .B(p_input[34675]), .Z(n11835) );
  AND U17755 ( .A(n11837), .B(n11838), .Z(o[4674]) );
  AND U17756 ( .A(p_input[24674]), .B(p_input[14674]), .Z(n11838) );
  AND U17757 ( .A(p_input[4674]), .B(p_input[34674]), .Z(n11837) );
  AND U17758 ( .A(n11839), .B(n11840), .Z(o[4673]) );
  AND U17759 ( .A(p_input[24673]), .B(p_input[14673]), .Z(n11840) );
  AND U17760 ( .A(p_input[4673]), .B(p_input[34673]), .Z(n11839) );
  AND U17761 ( .A(n11841), .B(n11842), .Z(o[4672]) );
  AND U17762 ( .A(p_input[24672]), .B(p_input[14672]), .Z(n11842) );
  AND U17763 ( .A(p_input[4672]), .B(p_input[34672]), .Z(n11841) );
  AND U17764 ( .A(n11843), .B(n11844), .Z(o[4671]) );
  AND U17765 ( .A(p_input[24671]), .B(p_input[14671]), .Z(n11844) );
  AND U17766 ( .A(p_input[4671]), .B(p_input[34671]), .Z(n11843) );
  AND U17767 ( .A(n11845), .B(n11846), .Z(o[4670]) );
  AND U17768 ( .A(p_input[24670]), .B(p_input[14670]), .Z(n11846) );
  AND U17769 ( .A(p_input[4670]), .B(p_input[34670]), .Z(n11845) );
  AND U17770 ( .A(n11847), .B(n11848), .Z(o[466]) );
  AND U17771 ( .A(p_input[20466]), .B(p_input[10466]), .Z(n11848) );
  AND U17772 ( .A(p_input[466]), .B(p_input[30466]), .Z(n11847) );
  AND U17773 ( .A(n11849), .B(n11850), .Z(o[4669]) );
  AND U17774 ( .A(p_input[24669]), .B(p_input[14669]), .Z(n11850) );
  AND U17775 ( .A(p_input[4669]), .B(p_input[34669]), .Z(n11849) );
  AND U17776 ( .A(n11851), .B(n11852), .Z(o[4668]) );
  AND U17777 ( .A(p_input[24668]), .B(p_input[14668]), .Z(n11852) );
  AND U17778 ( .A(p_input[4668]), .B(p_input[34668]), .Z(n11851) );
  AND U17779 ( .A(n11853), .B(n11854), .Z(o[4667]) );
  AND U17780 ( .A(p_input[24667]), .B(p_input[14667]), .Z(n11854) );
  AND U17781 ( .A(p_input[4667]), .B(p_input[34667]), .Z(n11853) );
  AND U17782 ( .A(n11855), .B(n11856), .Z(o[4666]) );
  AND U17783 ( .A(p_input[24666]), .B(p_input[14666]), .Z(n11856) );
  AND U17784 ( .A(p_input[4666]), .B(p_input[34666]), .Z(n11855) );
  AND U17785 ( .A(n11857), .B(n11858), .Z(o[4665]) );
  AND U17786 ( .A(p_input[24665]), .B(p_input[14665]), .Z(n11858) );
  AND U17787 ( .A(p_input[4665]), .B(p_input[34665]), .Z(n11857) );
  AND U17788 ( .A(n11859), .B(n11860), .Z(o[4664]) );
  AND U17789 ( .A(p_input[24664]), .B(p_input[14664]), .Z(n11860) );
  AND U17790 ( .A(p_input[4664]), .B(p_input[34664]), .Z(n11859) );
  AND U17791 ( .A(n11861), .B(n11862), .Z(o[4663]) );
  AND U17792 ( .A(p_input[24663]), .B(p_input[14663]), .Z(n11862) );
  AND U17793 ( .A(p_input[4663]), .B(p_input[34663]), .Z(n11861) );
  AND U17794 ( .A(n11863), .B(n11864), .Z(o[4662]) );
  AND U17795 ( .A(p_input[24662]), .B(p_input[14662]), .Z(n11864) );
  AND U17796 ( .A(p_input[4662]), .B(p_input[34662]), .Z(n11863) );
  AND U17797 ( .A(n11865), .B(n11866), .Z(o[4661]) );
  AND U17798 ( .A(p_input[24661]), .B(p_input[14661]), .Z(n11866) );
  AND U17799 ( .A(p_input[4661]), .B(p_input[34661]), .Z(n11865) );
  AND U17800 ( .A(n11867), .B(n11868), .Z(o[4660]) );
  AND U17801 ( .A(p_input[24660]), .B(p_input[14660]), .Z(n11868) );
  AND U17802 ( .A(p_input[4660]), .B(p_input[34660]), .Z(n11867) );
  AND U17803 ( .A(n11869), .B(n11870), .Z(o[465]) );
  AND U17804 ( .A(p_input[20465]), .B(p_input[10465]), .Z(n11870) );
  AND U17805 ( .A(p_input[465]), .B(p_input[30465]), .Z(n11869) );
  AND U17806 ( .A(n11871), .B(n11872), .Z(o[4659]) );
  AND U17807 ( .A(p_input[24659]), .B(p_input[14659]), .Z(n11872) );
  AND U17808 ( .A(p_input[4659]), .B(p_input[34659]), .Z(n11871) );
  AND U17809 ( .A(n11873), .B(n11874), .Z(o[4658]) );
  AND U17810 ( .A(p_input[24658]), .B(p_input[14658]), .Z(n11874) );
  AND U17811 ( .A(p_input[4658]), .B(p_input[34658]), .Z(n11873) );
  AND U17812 ( .A(n11875), .B(n11876), .Z(o[4657]) );
  AND U17813 ( .A(p_input[24657]), .B(p_input[14657]), .Z(n11876) );
  AND U17814 ( .A(p_input[4657]), .B(p_input[34657]), .Z(n11875) );
  AND U17815 ( .A(n11877), .B(n11878), .Z(o[4656]) );
  AND U17816 ( .A(p_input[24656]), .B(p_input[14656]), .Z(n11878) );
  AND U17817 ( .A(p_input[4656]), .B(p_input[34656]), .Z(n11877) );
  AND U17818 ( .A(n11879), .B(n11880), .Z(o[4655]) );
  AND U17819 ( .A(p_input[24655]), .B(p_input[14655]), .Z(n11880) );
  AND U17820 ( .A(p_input[4655]), .B(p_input[34655]), .Z(n11879) );
  AND U17821 ( .A(n11881), .B(n11882), .Z(o[4654]) );
  AND U17822 ( .A(p_input[24654]), .B(p_input[14654]), .Z(n11882) );
  AND U17823 ( .A(p_input[4654]), .B(p_input[34654]), .Z(n11881) );
  AND U17824 ( .A(n11883), .B(n11884), .Z(o[4653]) );
  AND U17825 ( .A(p_input[24653]), .B(p_input[14653]), .Z(n11884) );
  AND U17826 ( .A(p_input[4653]), .B(p_input[34653]), .Z(n11883) );
  AND U17827 ( .A(n11885), .B(n11886), .Z(o[4652]) );
  AND U17828 ( .A(p_input[24652]), .B(p_input[14652]), .Z(n11886) );
  AND U17829 ( .A(p_input[4652]), .B(p_input[34652]), .Z(n11885) );
  AND U17830 ( .A(n11887), .B(n11888), .Z(o[4651]) );
  AND U17831 ( .A(p_input[24651]), .B(p_input[14651]), .Z(n11888) );
  AND U17832 ( .A(p_input[4651]), .B(p_input[34651]), .Z(n11887) );
  AND U17833 ( .A(n11889), .B(n11890), .Z(o[4650]) );
  AND U17834 ( .A(p_input[24650]), .B(p_input[14650]), .Z(n11890) );
  AND U17835 ( .A(p_input[4650]), .B(p_input[34650]), .Z(n11889) );
  AND U17836 ( .A(n11891), .B(n11892), .Z(o[464]) );
  AND U17837 ( .A(p_input[20464]), .B(p_input[10464]), .Z(n11892) );
  AND U17838 ( .A(p_input[464]), .B(p_input[30464]), .Z(n11891) );
  AND U17839 ( .A(n11893), .B(n11894), .Z(o[4649]) );
  AND U17840 ( .A(p_input[24649]), .B(p_input[14649]), .Z(n11894) );
  AND U17841 ( .A(p_input[4649]), .B(p_input[34649]), .Z(n11893) );
  AND U17842 ( .A(n11895), .B(n11896), .Z(o[4648]) );
  AND U17843 ( .A(p_input[24648]), .B(p_input[14648]), .Z(n11896) );
  AND U17844 ( .A(p_input[4648]), .B(p_input[34648]), .Z(n11895) );
  AND U17845 ( .A(n11897), .B(n11898), .Z(o[4647]) );
  AND U17846 ( .A(p_input[24647]), .B(p_input[14647]), .Z(n11898) );
  AND U17847 ( .A(p_input[4647]), .B(p_input[34647]), .Z(n11897) );
  AND U17848 ( .A(n11899), .B(n11900), .Z(o[4646]) );
  AND U17849 ( .A(p_input[24646]), .B(p_input[14646]), .Z(n11900) );
  AND U17850 ( .A(p_input[4646]), .B(p_input[34646]), .Z(n11899) );
  AND U17851 ( .A(n11901), .B(n11902), .Z(o[4645]) );
  AND U17852 ( .A(p_input[24645]), .B(p_input[14645]), .Z(n11902) );
  AND U17853 ( .A(p_input[4645]), .B(p_input[34645]), .Z(n11901) );
  AND U17854 ( .A(n11903), .B(n11904), .Z(o[4644]) );
  AND U17855 ( .A(p_input[24644]), .B(p_input[14644]), .Z(n11904) );
  AND U17856 ( .A(p_input[4644]), .B(p_input[34644]), .Z(n11903) );
  AND U17857 ( .A(n11905), .B(n11906), .Z(o[4643]) );
  AND U17858 ( .A(p_input[24643]), .B(p_input[14643]), .Z(n11906) );
  AND U17859 ( .A(p_input[4643]), .B(p_input[34643]), .Z(n11905) );
  AND U17860 ( .A(n11907), .B(n11908), .Z(o[4642]) );
  AND U17861 ( .A(p_input[24642]), .B(p_input[14642]), .Z(n11908) );
  AND U17862 ( .A(p_input[4642]), .B(p_input[34642]), .Z(n11907) );
  AND U17863 ( .A(n11909), .B(n11910), .Z(o[4641]) );
  AND U17864 ( .A(p_input[24641]), .B(p_input[14641]), .Z(n11910) );
  AND U17865 ( .A(p_input[4641]), .B(p_input[34641]), .Z(n11909) );
  AND U17866 ( .A(n11911), .B(n11912), .Z(o[4640]) );
  AND U17867 ( .A(p_input[24640]), .B(p_input[14640]), .Z(n11912) );
  AND U17868 ( .A(p_input[4640]), .B(p_input[34640]), .Z(n11911) );
  AND U17869 ( .A(n11913), .B(n11914), .Z(o[463]) );
  AND U17870 ( .A(p_input[20463]), .B(p_input[10463]), .Z(n11914) );
  AND U17871 ( .A(p_input[463]), .B(p_input[30463]), .Z(n11913) );
  AND U17872 ( .A(n11915), .B(n11916), .Z(o[4639]) );
  AND U17873 ( .A(p_input[24639]), .B(p_input[14639]), .Z(n11916) );
  AND U17874 ( .A(p_input[4639]), .B(p_input[34639]), .Z(n11915) );
  AND U17875 ( .A(n11917), .B(n11918), .Z(o[4638]) );
  AND U17876 ( .A(p_input[24638]), .B(p_input[14638]), .Z(n11918) );
  AND U17877 ( .A(p_input[4638]), .B(p_input[34638]), .Z(n11917) );
  AND U17878 ( .A(n11919), .B(n11920), .Z(o[4637]) );
  AND U17879 ( .A(p_input[24637]), .B(p_input[14637]), .Z(n11920) );
  AND U17880 ( .A(p_input[4637]), .B(p_input[34637]), .Z(n11919) );
  AND U17881 ( .A(n11921), .B(n11922), .Z(o[4636]) );
  AND U17882 ( .A(p_input[24636]), .B(p_input[14636]), .Z(n11922) );
  AND U17883 ( .A(p_input[4636]), .B(p_input[34636]), .Z(n11921) );
  AND U17884 ( .A(n11923), .B(n11924), .Z(o[4635]) );
  AND U17885 ( .A(p_input[24635]), .B(p_input[14635]), .Z(n11924) );
  AND U17886 ( .A(p_input[4635]), .B(p_input[34635]), .Z(n11923) );
  AND U17887 ( .A(n11925), .B(n11926), .Z(o[4634]) );
  AND U17888 ( .A(p_input[24634]), .B(p_input[14634]), .Z(n11926) );
  AND U17889 ( .A(p_input[4634]), .B(p_input[34634]), .Z(n11925) );
  AND U17890 ( .A(n11927), .B(n11928), .Z(o[4633]) );
  AND U17891 ( .A(p_input[24633]), .B(p_input[14633]), .Z(n11928) );
  AND U17892 ( .A(p_input[4633]), .B(p_input[34633]), .Z(n11927) );
  AND U17893 ( .A(n11929), .B(n11930), .Z(o[4632]) );
  AND U17894 ( .A(p_input[24632]), .B(p_input[14632]), .Z(n11930) );
  AND U17895 ( .A(p_input[4632]), .B(p_input[34632]), .Z(n11929) );
  AND U17896 ( .A(n11931), .B(n11932), .Z(o[4631]) );
  AND U17897 ( .A(p_input[24631]), .B(p_input[14631]), .Z(n11932) );
  AND U17898 ( .A(p_input[4631]), .B(p_input[34631]), .Z(n11931) );
  AND U17899 ( .A(n11933), .B(n11934), .Z(o[4630]) );
  AND U17900 ( .A(p_input[24630]), .B(p_input[14630]), .Z(n11934) );
  AND U17901 ( .A(p_input[4630]), .B(p_input[34630]), .Z(n11933) );
  AND U17902 ( .A(n11935), .B(n11936), .Z(o[462]) );
  AND U17903 ( .A(p_input[20462]), .B(p_input[10462]), .Z(n11936) );
  AND U17904 ( .A(p_input[462]), .B(p_input[30462]), .Z(n11935) );
  AND U17905 ( .A(n11937), .B(n11938), .Z(o[4629]) );
  AND U17906 ( .A(p_input[24629]), .B(p_input[14629]), .Z(n11938) );
  AND U17907 ( .A(p_input[4629]), .B(p_input[34629]), .Z(n11937) );
  AND U17908 ( .A(n11939), .B(n11940), .Z(o[4628]) );
  AND U17909 ( .A(p_input[24628]), .B(p_input[14628]), .Z(n11940) );
  AND U17910 ( .A(p_input[4628]), .B(p_input[34628]), .Z(n11939) );
  AND U17911 ( .A(n11941), .B(n11942), .Z(o[4627]) );
  AND U17912 ( .A(p_input[24627]), .B(p_input[14627]), .Z(n11942) );
  AND U17913 ( .A(p_input[4627]), .B(p_input[34627]), .Z(n11941) );
  AND U17914 ( .A(n11943), .B(n11944), .Z(o[4626]) );
  AND U17915 ( .A(p_input[24626]), .B(p_input[14626]), .Z(n11944) );
  AND U17916 ( .A(p_input[4626]), .B(p_input[34626]), .Z(n11943) );
  AND U17917 ( .A(n11945), .B(n11946), .Z(o[4625]) );
  AND U17918 ( .A(p_input[24625]), .B(p_input[14625]), .Z(n11946) );
  AND U17919 ( .A(p_input[4625]), .B(p_input[34625]), .Z(n11945) );
  AND U17920 ( .A(n11947), .B(n11948), .Z(o[4624]) );
  AND U17921 ( .A(p_input[24624]), .B(p_input[14624]), .Z(n11948) );
  AND U17922 ( .A(p_input[4624]), .B(p_input[34624]), .Z(n11947) );
  AND U17923 ( .A(n11949), .B(n11950), .Z(o[4623]) );
  AND U17924 ( .A(p_input[24623]), .B(p_input[14623]), .Z(n11950) );
  AND U17925 ( .A(p_input[4623]), .B(p_input[34623]), .Z(n11949) );
  AND U17926 ( .A(n11951), .B(n11952), .Z(o[4622]) );
  AND U17927 ( .A(p_input[24622]), .B(p_input[14622]), .Z(n11952) );
  AND U17928 ( .A(p_input[4622]), .B(p_input[34622]), .Z(n11951) );
  AND U17929 ( .A(n11953), .B(n11954), .Z(o[4621]) );
  AND U17930 ( .A(p_input[24621]), .B(p_input[14621]), .Z(n11954) );
  AND U17931 ( .A(p_input[4621]), .B(p_input[34621]), .Z(n11953) );
  AND U17932 ( .A(n11955), .B(n11956), .Z(o[4620]) );
  AND U17933 ( .A(p_input[24620]), .B(p_input[14620]), .Z(n11956) );
  AND U17934 ( .A(p_input[4620]), .B(p_input[34620]), .Z(n11955) );
  AND U17935 ( .A(n11957), .B(n11958), .Z(o[461]) );
  AND U17936 ( .A(p_input[20461]), .B(p_input[10461]), .Z(n11958) );
  AND U17937 ( .A(p_input[461]), .B(p_input[30461]), .Z(n11957) );
  AND U17938 ( .A(n11959), .B(n11960), .Z(o[4619]) );
  AND U17939 ( .A(p_input[24619]), .B(p_input[14619]), .Z(n11960) );
  AND U17940 ( .A(p_input[4619]), .B(p_input[34619]), .Z(n11959) );
  AND U17941 ( .A(n11961), .B(n11962), .Z(o[4618]) );
  AND U17942 ( .A(p_input[24618]), .B(p_input[14618]), .Z(n11962) );
  AND U17943 ( .A(p_input[4618]), .B(p_input[34618]), .Z(n11961) );
  AND U17944 ( .A(n11963), .B(n11964), .Z(o[4617]) );
  AND U17945 ( .A(p_input[24617]), .B(p_input[14617]), .Z(n11964) );
  AND U17946 ( .A(p_input[4617]), .B(p_input[34617]), .Z(n11963) );
  AND U17947 ( .A(n11965), .B(n11966), .Z(o[4616]) );
  AND U17948 ( .A(p_input[24616]), .B(p_input[14616]), .Z(n11966) );
  AND U17949 ( .A(p_input[4616]), .B(p_input[34616]), .Z(n11965) );
  AND U17950 ( .A(n11967), .B(n11968), .Z(o[4615]) );
  AND U17951 ( .A(p_input[24615]), .B(p_input[14615]), .Z(n11968) );
  AND U17952 ( .A(p_input[4615]), .B(p_input[34615]), .Z(n11967) );
  AND U17953 ( .A(n11969), .B(n11970), .Z(o[4614]) );
  AND U17954 ( .A(p_input[24614]), .B(p_input[14614]), .Z(n11970) );
  AND U17955 ( .A(p_input[4614]), .B(p_input[34614]), .Z(n11969) );
  AND U17956 ( .A(n11971), .B(n11972), .Z(o[4613]) );
  AND U17957 ( .A(p_input[24613]), .B(p_input[14613]), .Z(n11972) );
  AND U17958 ( .A(p_input[4613]), .B(p_input[34613]), .Z(n11971) );
  AND U17959 ( .A(n11973), .B(n11974), .Z(o[4612]) );
  AND U17960 ( .A(p_input[24612]), .B(p_input[14612]), .Z(n11974) );
  AND U17961 ( .A(p_input[4612]), .B(p_input[34612]), .Z(n11973) );
  AND U17962 ( .A(n11975), .B(n11976), .Z(o[4611]) );
  AND U17963 ( .A(p_input[24611]), .B(p_input[14611]), .Z(n11976) );
  AND U17964 ( .A(p_input[4611]), .B(p_input[34611]), .Z(n11975) );
  AND U17965 ( .A(n11977), .B(n11978), .Z(o[4610]) );
  AND U17966 ( .A(p_input[24610]), .B(p_input[14610]), .Z(n11978) );
  AND U17967 ( .A(p_input[4610]), .B(p_input[34610]), .Z(n11977) );
  AND U17968 ( .A(n11979), .B(n11980), .Z(o[460]) );
  AND U17969 ( .A(p_input[20460]), .B(p_input[10460]), .Z(n11980) );
  AND U17970 ( .A(p_input[460]), .B(p_input[30460]), .Z(n11979) );
  AND U17971 ( .A(n11981), .B(n11982), .Z(o[4609]) );
  AND U17972 ( .A(p_input[24609]), .B(p_input[14609]), .Z(n11982) );
  AND U17973 ( .A(p_input[4609]), .B(p_input[34609]), .Z(n11981) );
  AND U17974 ( .A(n11983), .B(n11984), .Z(o[4608]) );
  AND U17975 ( .A(p_input[24608]), .B(p_input[14608]), .Z(n11984) );
  AND U17976 ( .A(p_input[4608]), .B(p_input[34608]), .Z(n11983) );
  AND U17977 ( .A(n11985), .B(n11986), .Z(o[4607]) );
  AND U17978 ( .A(p_input[24607]), .B(p_input[14607]), .Z(n11986) );
  AND U17979 ( .A(p_input[4607]), .B(p_input[34607]), .Z(n11985) );
  AND U17980 ( .A(n11987), .B(n11988), .Z(o[4606]) );
  AND U17981 ( .A(p_input[24606]), .B(p_input[14606]), .Z(n11988) );
  AND U17982 ( .A(p_input[4606]), .B(p_input[34606]), .Z(n11987) );
  AND U17983 ( .A(n11989), .B(n11990), .Z(o[4605]) );
  AND U17984 ( .A(p_input[24605]), .B(p_input[14605]), .Z(n11990) );
  AND U17985 ( .A(p_input[4605]), .B(p_input[34605]), .Z(n11989) );
  AND U17986 ( .A(n11991), .B(n11992), .Z(o[4604]) );
  AND U17987 ( .A(p_input[24604]), .B(p_input[14604]), .Z(n11992) );
  AND U17988 ( .A(p_input[4604]), .B(p_input[34604]), .Z(n11991) );
  AND U17989 ( .A(n11993), .B(n11994), .Z(o[4603]) );
  AND U17990 ( .A(p_input[24603]), .B(p_input[14603]), .Z(n11994) );
  AND U17991 ( .A(p_input[4603]), .B(p_input[34603]), .Z(n11993) );
  AND U17992 ( .A(n11995), .B(n11996), .Z(o[4602]) );
  AND U17993 ( .A(p_input[24602]), .B(p_input[14602]), .Z(n11996) );
  AND U17994 ( .A(p_input[4602]), .B(p_input[34602]), .Z(n11995) );
  AND U17995 ( .A(n11997), .B(n11998), .Z(o[4601]) );
  AND U17996 ( .A(p_input[24601]), .B(p_input[14601]), .Z(n11998) );
  AND U17997 ( .A(p_input[4601]), .B(p_input[34601]), .Z(n11997) );
  AND U17998 ( .A(n11999), .B(n12000), .Z(o[4600]) );
  AND U17999 ( .A(p_input[24600]), .B(p_input[14600]), .Z(n12000) );
  AND U18000 ( .A(p_input[4600]), .B(p_input[34600]), .Z(n11999) );
  AND U18001 ( .A(n12001), .B(n12002), .Z(o[45]) );
  AND U18002 ( .A(p_input[20045]), .B(p_input[10045]), .Z(n12002) );
  AND U18003 ( .A(p_input[45]), .B(p_input[30045]), .Z(n12001) );
  AND U18004 ( .A(n12003), .B(n12004), .Z(o[459]) );
  AND U18005 ( .A(p_input[20459]), .B(p_input[10459]), .Z(n12004) );
  AND U18006 ( .A(p_input[459]), .B(p_input[30459]), .Z(n12003) );
  AND U18007 ( .A(n12005), .B(n12006), .Z(o[4599]) );
  AND U18008 ( .A(p_input[24599]), .B(p_input[14599]), .Z(n12006) );
  AND U18009 ( .A(p_input[4599]), .B(p_input[34599]), .Z(n12005) );
  AND U18010 ( .A(n12007), .B(n12008), .Z(o[4598]) );
  AND U18011 ( .A(p_input[24598]), .B(p_input[14598]), .Z(n12008) );
  AND U18012 ( .A(p_input[4598]), .B(p_input[34598]), .Z(n12007) );
  AND U18013 ( .A(n12009), .B(n12010), .Z(o[4597]) );
  AND U18014 ( .A(p_input[24597]), .B(p_input[14597]), .Z(n12010) );
  AND U18015 ( .A(p_input[4597]), .B(p_input[34597]), .Z(n12009) );
  AND U18016 ( .A(n12011), .B(n12012), .Z(o[4596]) );
  AND U18017 ( .A(p_input[24596]), .B(p_input[14596]), .Z(n12012) );
  AND U18018 ( .A(p_input[4596]), .B(p_input[34596]), .Z(n12011) );
  AND U18019 ( .A(n12013), .B(n12014), .Z(o[4595]) );
  AND U18020 ( .A(p_input[24595]), .B(p_input[14595]), .Z(n12014) );
  AND U18021 ( .A(p_input[4595]), .B(p_input[34595]), .Z(n12013) );
  AND U18022 ( .A(n12015), .B(n12016), .Z(o[4594]) );
  AND U18023 ( .A(p_input[24594]), .B(p_input[14594]), .Z(n12016) );
  AND U18024 ( .A(p_input[4594]), .B(p_input[34594]), .Z(n12015) );
  AND U18025 ( .A(n12017), .B(n12018), .Z(o[4593]) );
  AND U18026 ( .A(p_input[24593]), .B(p_input[14593]), .Z(n12018) );
  AND U18027 ( .A(p_input[4593]), .B(p_input[34593]), .Z(n12017) );
  AND U18028 ( .A(n12019), .B(n12020), .Z(o[4592]) );
  AND U18029 ( .A(p_input[24592]), .B(p_input[14592]), .Z(n12020) );
  AND U18030 ( .A(p_input[4592]), .B(p_input[34592]), .Z(n12019) );
  AND U18031 ( .A(n12021), .B(n12022), .Z(o[4591]) );
  AND U18032 ( .A(p_input[24591]), .B(p_input[14591]), .Z(n12022) );
  AND U18033 ( .A(p_input[4591]), .B(p_input[34591]), .Z(n12021) );
  AND U18034 ( .A(n12023), .B(n12024), .Z(o[4590]) );
  AND U18035 ( .A(p_input[24590]), .B(p_input[14590]), .Z(n12024) );
  AND U18036 ( .A(p_input[4590]), .B(p_input[34590]), .Z(n12023) );
  AND U18037 ( .A(n12025), .B(n12026), .Z(o[458]) );
  AND U18038 ( .A(p_input[20458]), .B(p_input[10458]), .Z(n12026) );
  AND U18039 ( .A(p_input[458]), .B(p_input[30458]), .Z(n12025) );
  AND U18040 ( .A(n12027), .B(n12028), .Z(o[4589]) );
  AND U18041 ( .A(p_input[24589]), .B(p_input[14589]), .Z(n12028) );
  AND U18042 ( .A(p_input[4589]), .B(p_input[34589]), .Z(n12027) );
  AND U18043 ( .A(n12029), .B(n12030), .Z(o[4588]) );
  AND U18044 ( .A(p_input[24588]), .B(p_input[14588]), .Z(n12030) );
  AND U18045 ( .A(p_input[4588]), .B(p_input[34588]), .Z(n12029) );
  AND U18046 ( .A(n12031), .B(n12032), .Z(o[4587]) );
  AND U18047 ( .A(p_input[24587]), .B(p_input[14587]), .Z(n12032) );
  AND U18048 ( .A(p_input[4587]), .B(p_input[34587]), .Z(n12031) );
  AND U18049 ( .A(n12033), .B(n12034), .Z(o[4586]) );
  AND U18050 ( .A(p_input[24586]), .B(p_input[14586]), .Z(n12034) );
  AND U18051 ( .A(p_input[4586]), .B(p_input[34586]), .Z(n12033) );
  AND U18052 ( .A(n12035), .B(n12036), .Z(o[4585]) );
  AND U18053 ( .A(p_input[24585]), .B(p_input[14585]), .Z(n12036) );
  AND U18054 ( .A(p_input[4585]), .B(p_input[34585]), .Z(n12035) );
  AND U18055 ( .A(n12037), .B(n12038), .Z(o[4584]) );
  AND U18056 ( .A(p_input[24584]), .B(p_input[14584]), .Z(n12038) );
  AND U18057 ( .A(p_input[4584]), .B(p_input[34584]), .Z(n12037) );
  AND U18058 ( .A(n12039), .B(n12040), .Z(o[4583]) );
  AND U18059 ( .A(p_input[24583]), .B(p_input[14583]), .Z(n12040) );
  AND U18060 ( .A(p_input[4583]), .B(p_input[34583]), .Z(n12039) );
  AND U18061 ( .A(n12041), .B(n12042), .Z(o[4582]) );
  AND U18062 ( .A(p_input[24582]), .B(p_input[14582]), .Z(n12042) );
  AND U18063 ( .A(p_input[4582]), .B(p_input[34582]), .Z(n12041) );
  AND U18064 ( .A(n12043), .B(n12044), .Z(o[4581]) );
  AND U18065 ( .A(p_input[24581]), .B(p_input[14581]), .Z(n12044) );
  AND U18066 ( .A(p_input[4581]), .B(p_input[34581]), .Z(n12043) );
  AND U18067 ( .A(n12045), .B(n12046), .Z(o[4580]) );
  AND U18068 ( .A(p_input[24580]), .B(p_input[14580]), .Z(n12046) );
  AND U18069 ( .A(p_input[4580]), .B(p_input[34580]), .Z(n12045) );
  AND U18070 ( .A(n12047), .B(n12048), .Z(o[457]) );
  AND U18071 ( .A(p_input[20457]), .B(p_input[10457]), .Z(n12048) );
  AND U18072 ( .A(p_input[457]), .B(p_input[30457]), .Z(n12047) );
  AND U18073 ( .A(n12049), .B(n12050), .Z(o[4579]) );
  AND U18074 ( .A(p_input[24579]), .B(p_input[14579]), .Z(n12050) );
  AND U18075 ( .A(p_input[4579]), .B(p_input[34579]), .Z(n12049) );
  AND U18076 ( .A(n12051), .B(n12052), .Z(o[4578]) );
  AND U18077 ( .A(p_input[24578]), .B(p_input[14578]), .Z(n12052) );
  AND U18078 ( .A(p_input[4578]), .B(p_input[34578]), .Z(n12051) );
  AND U18079 ( .A(n12053), .B(n12054), .Z(o[4577]) );
  AND U18080 ( .A(p_input[24577]), .B(p_input[14577]), .Z(n12054) );
  AND U18081 ( .A(p_input[4577]), .B(p_input[34577]), .Z(n12053) );
  AND U18082 ( .A(n12055), .B(n12056), .Z(o[4576]) );
  AND U18083 ( .A(p_input[24576]), .B(p_input[14576]), .Z(n12056) );
  AND U18084 ( .A(p_input[4576]), .B(p_input[34576]), .Z(n12055) );
  AND U18085 ( .A(n12057), .B(n12058), .Z(o[4575]) );
  AND U18086 ( .A(p_input[24575]), .B(p_input[14575]), .Z(n12058) );
  AND U18087 ( .A(p_input[4575]), .B(p_input[34575]), .Z(n12057) );
  AND U18088 ( .A(n12059), .B(n12060), .Z(o[4574]) );
  AND U18089 ( .A(p_input[24574]), .B(p_input[14574]), .Z(n12060) );
  AND U18090 ( .A(p_input[4574]), .B(p_input[34574]), .Z(n12059) );
  AND U18091 ( .A(n12061), .B(n12062), .Z(o[4573]) );
  AND U18092 ( .A(p_input[24573]), .B(p_input[14573]), .Z(n12062) );
  AND U18093 ( .A(p_input[4573]), .B(p_input[34573]), .Z(n12061) );
  AND U18094 ( .A(n12063), .B(n12064), .Z(o[4572]) );
  AND U18095 ( .A(p_input[24572]), .B(p_input[14572]), .Z(n12064) );
  AND U18096 ( .A(p_input[4572]), .B(p_input[34572]), .Z(n12063) );
  AND U18097 ( .A(n12065), .B(n12066), .Z(o[4571]) );
  AND U18098 ( .A(p_input[24571]), .B(p_input[14571]), .Z(n12066) );
  AND U18099 ( .A(p_input[4571]), .B(p_input[34571]), .Z(n12065) );
  AND U18100 ( .A(n12067), .B(n12068), .Z(o[4570]) );
  AND U18101 ( .A(p_input[24570]), .B(p_input[14570]), .Z(n12068) );
  AND U18102 ( .A(p_input[4570]), .B(p_input[34570]), .Z(n12067) );
  AND U18103 ( .A(n12069), .B(n12070), .Z(o[456]) );
  AND U18104 ( .A(p_input[20456]), .B(p_input[10456]), .Z(n12070) );
  AND U18105 ( .A(p_input[456]), .B(p_input[30456]), .Z(n12069) );
  AND U18106 ( .A(n12071), .B(n12072), .Z(o[4569]) );
  AND U18107 ( .A(p_input[24569]), .B(p_input[14569]), .Z(n12072) );
  AND U18108 ( .A(p_input[4569]), .B(p_input[34569]), .Z(n12071) );
  AND U18109 ( .A(n12073), .B(n12074), .Z(o[4568]) );
  AND U18110 ( .A(p_input[24568]), .B(p_input[14568]), .Z(n12074) );
  AND U18111 ( .A(p_input[4568]), .B(p_input[34568]), .Z(n12073) );
  AND U18112 ( .A(n12075), .B(n12076), .Z(o[4567]) );
  AND U18113 ( .A(p_input[24567]), .B(p_input[14567]), .Z(n12076) );
  AND U18114 ( .A(p_input[4567]), .B(p_input[34567]), .Z(n12075) );
  AND U18115 ( .A(n12077), .B(n12078), .Z(o[4566]) );
  AND U18116 ( .A(p_input[24566]), .B(p_input[14566]), .Z(n12078) );
  AND U18117 ( .A(p_input[4566]), .B(p_input[34566]), .Z(n12077) );
  AND U18118 ( .A(n12079), .B(n12080), .Z(o[4565]) );
  AND U18119 ( .A(p_input[24565]), .B(p_input[14565]), .Z(n12080) );
  AND U18120 ( .A(p_input[4565]), .B(p_input[34565]), .Z(n12079) );
  AND U18121 ( .A(n12081), .B(n12082), .Z(o[4564]) );
  AND U18122 ( .A(p_input[24564]), .B(p_input[14564]), .Z(n12082) );
  AND U18123 ( .A(p_input[4564]), .B(p_input[34564]), .Z(n12081) );
  AND U18124 ( .A(n12083), .B(n12084), .Z(o[4563]) );
  AND U18125 ( .A(p_input[24563]), .B(p_input[14563]), .Z(n12084) );
  AND U18126 ( .A(p_input[4563]), .B(p_input[34563]), .Z(n12083) );
  AND U18127 ( .A(n12085), .B(n12086), .Z(o[4562]) );
  AND U18128 ( .A(p_input[24562]), .B(p_input[14562]), .Z(n12086) );
  AND U18129 ( .A(p_input[4562]), .B(p_input[34562]), .Z(n12085) );
  AND U18130 ( .A(n12087), .B(n12088), .Z(o[4561]) );
  AND U18131 ( .A(p_input[24561]), .B(p_input[14561]), .Z(n12088) );
  AND U18132 ( .A(p_input[4561]), .B(p_input[34561]), .Z(n12087) );
  AND U18133 ( .A(n12089), .B(n12090), .Z(o[4560]) );
  AND U18134 ( .A(p_input[24560]), .B(p_input[14560]), .Z(n12090) );
  AND U18135 ( .A(p_input[4560]), .B(p_input[34560]), .Z(n12089) );
  AND U18136 ( .A(n12091), .B(n12092), .Z(o[455]) );
  AND U18137 ( .A(p_input[20455]), .B(p_input[10455]), .Z(n12092) );
  AND U18138 ( .A(p_input[455]), .B(p_input[30455]), .Z(n12091) );
  AND U18139 ( .A(n12093), .B(n12094), .Z(o[4559]) );
  AND U18140 ( .A(p_input[24559]), .B(p_input[14559]), .Z(n12094) );
  AND U18141 ( .A(p_input[4559]), .B(p_input[34559]), .Z(n12093) );
  AND U18142 ( .A(n12095), .B(n12096), .Z(o[4558]) );
  AND U18143 ( .A(p_input[24558]), .B(p_input[14558]), .Z(n12096) );
  AND U18144 ( .A(p_input[4558]), .B(p_input[34558]), .Z(n12095) );
  AND U18145 ( .A(n12097), .B(n12098), .Z(o[4557]) );
  AND U18146 ( .A(p_input[24557]), .B(p_input[14557]), .Z(n12098) );
  AND U18147 ( .A(p_input[4557]), .B(p_input[34557]), .Z(n12097) );
  AND U18148 ( .A(n12099), .B(n12100), .Z(o[4556]) );
  AND U18149 ( .A(p_input[24556]), .B(p_input[14556]), .Z(n12100) );
  AND U18150 ( .A(p_input[4556]), .B(p_input[34556]), .Z(n12099) );
  AND U18151 ( .A(n12101), .B(n12102), .Z(o[4555]) );
  AND U18152 ( .A(p_input[24555]), .B(p_input[14555]), .Z(n12102) );
  AND U18153 ( .A(p_input[4555]), .B(p_input[34555]), .Z(n12101) );
  AND U18154 ( .A(n12103), .B(n12104), .Z(o[4554]) );
  AND U18155 ( .A(p_input[24554]), .B(p_input[14554]), .Z(n12104) );
  AND U18156 ( .A(p_input[4554]), .B(p_input[34554]), .Z(n12103) );
  AND U18157 ( .A(n12105), .B(n12106), .Z(o[4553]) );
  AND U18158 ( .A(p_input[24553]), .B(p_input[14553]), .Z(n12106) );
  AND U18159 ( .A(p_input[4553]), .B(p_input[34553]), .Z(n12105) );
  AND U18160 ( .A(n12107), .B(n12108), .Z(o[4552]) );
  AND U18161 ( .A(p_input[24552]), .B(p_input[14552]), .Z(n12108) );
  AND U18162 ( .A(p_input[4552]), .B(p_input[34552]), .Z(n12107) );
  AND U18163 ( .A(n12109), .B(n12110), .Z(o[4551]) );
  AND U18164 ( .A(p_input[24551]), .B(p_input[14551]), .Z(n12110) );
  AND U18165 ( .A(p_input[4551]), .B(p_input[34551]), .Z(n12109) );
  AND U18166 ( .A(n12111), .B(n12112), .Z(o[4550]) );
  AND U18167 ( .A(p_input[24550]), .B(p_input[14550]), .Z(n12112) );
  AND U18168 ( .A(p_input[4550]), .B(p_input[34550]), .Z(n12111) );
  AND U18169 ( .A(n12113), .B(n12114), .Z(o[454]) );
  AND U18170 ( .A(p_input[20454]), .B(p_input[10454]), .Z(n12114) );
  AND U18171 ( .A(p_input[454]), .B(p_input[30454]), .Z(n12113) );
  AND U18172 ( .A(n12115), .B(n12116), .Z(o[4549]) );
  AND U18173 ( .A(p_input[24549]), .B(p_input[14549]), .Z(n12116) );
  AND U18174 ( .A(p_input[4549]), .B(p_input[34549]), .Z(n12115) );
  AND U18175 ( .A(n12117), .B(n12118), .Z(o[4548]) );
  AND U18176 ( .A(p_input[24548]), .B(p_input[14548]), .Z(n12118) );
  AND U18177 ( .A(p_input[4548]), .B(p_input[34548]), .Z(n12117) );
  AND U18178 ( .A(n12119), .B(n12120), .Z(o[4547]) );
  AND U18179 ( .A(p_input[24547]), .B(p_input[14547]), .Z(n12120) );
  AND U18180 ( .A(p_input[4547]), .B(p_input[34547]), .Z(n12119) );
  AND U18181 ( .A(n12121), .B(n12122), .Z(o[4546]) );
  AND U18182 ( .A(p_input[24546]), .B(p_input[14546]), .Z(n12122) );
  AND U18183 ( .A(p_input[4546]), .B(p_input[34546]), .Z(n12121) );
  AND U18184 ( .A(n12123), .B(n12124), .Z(o[4545]) );
  AND U18185 ( .A(p_input[24545]), .B(p_input[14545]), .Z(n12124) );
  AND U18186 ( .A(p_input[4545]), .B(p_input[34545]), .Z(n12123) );
  AND U18187 ( .A(n12125), .B(n12126), .Z(o[4544]) );
  AND U18188 ( .A(p_input[24544]), .B(p_input[14544]), .Z(n12126) );
  AND U18189 ( .A(p_input[4544]), .B(p_input[34544]), .Z(n12125) );
  AND U18190 ( .A(n12127), .B(n12128), .Z(o[4543]) );
  AND U18191 ( .A(p_input[24543]), .B(p_input[14543]), .Z(n12128) );
  AND U18192 ( .A(p_input[4543]), .B(p_input[34543]), .Z(n12127) );
  AND U18193 ( .A(n12129), .B(n12130), .Z(o[4542]) );
  AND U18194 ( .A(p_input[24542]), .B(p_input[14542]), .Z(n12130) );
  AND U18195 ( .A(p_input[4542]), .B(p_input[34542]), .Z(n12129) );
  AND U18196 ( .A(n12131), .B(n12132), .Z(o[4541]) );
  AND U18197 ( .A(p_input[24541]), .B(p_input[14541]), .Z(n12132) );
  AND U18198 ( .A(p_input[4541]), .B(p_input[34541]), .Z(n12131) );
  AND U18199 ( .A(n12133), .B(n12134), .Z(o[4540]) );
  AND U18200 ( .A(p_input[24540]), .B(p_input[14540]), .Z(n12134) );
  AND U18201 ( .A(p_input[4540]), .B(p_input[34540]), .Z(n12133) );
  AND U18202 ( .A(n12135), .B(n12136), .Z(o[453]) );
  AND U18203 ( .A(p_input[20453]), .B(p_input[10453]), .Z(n12136) );
  AND U18204 ( .A(p_input[453]), .B(p_input[30453]), .Z(n12135) );
  AND U18205 ( .A(n12137), .B(n12138), .Z(o[4539]) );
  AND U18206 ( .A(p_input[24539]), .B(p_input[14539]), .Z(n12138) );
  AND U18207 ( .A(p_input[4539]), .B(p_input[34539]), .Z(n12137) );
  AND U18208 ( .A(n12139), .B(n12140), .Z(o[4538]) );
  AND U18209 ( .A(p_input[24538]), .B(p_input[14538]), .Z(n12140) );
  AND U18210 ( .A(p_input[4538]), .B(p_input[34538]), .Z(n12139) );
  AND U18211 ( .A(n12141), .B(n12142), .Z(o[4537]) );
  AND U18212 ( .A(p_input[24537]), .B(p_input[14537]), .Z(n12142) );
  AND U18213 ( .A(p_input[4537]), .B(p_input[34537]), .Z(n12141) );
  AND U18214 ( .A(n12143), .B(n12144), .Z(o[4536]) );
  AND U18215 ( .A(p_input[24536]), .B(p_input[14536]), .Z(n12144) );
  AND U18216 ( .A(p_input[4536]), .B(p_input[34536]), .Z(n12143) );
  AND U18217 ( .A(n12145), .B(n12146), .Z(o[4535]) );
  AND U18218 ( .A(p_input[24535]), .B(p_input[14535]), .Z(n12146) );
  AND U18219 ( .A(p_input[4535]), .B(p_input[34535]), .Z(n12145) );
  AND U18220 ( .A(n12147), .B(n12148), .Z(o[4534]) );
  AND U18221 ( .A(p_input[24534]), .B(p_input[14534]), .Z(n12148) );
  AND U18222 ( .A(p_input[4534]), .B(p_input[34534]), .Z(n12147) );
  AND U18223 ( .A(n12149), .B(n12150), .Z(o[4533]) );
  AND U18224 ( .A(p_input[24533]), .B(p_input[14533]), .Z(n12150) );
  AND U18225 ( .A(p_input[4533]), .B(p_input[34533]), .Z(n12149) );
  AND U18226 ( .A(n12151), .B(n12152), .Z(o[4532]) );
  AND U18227 ( .A(p_input[24532]), .B(p_input[14532]), .Z(n12152) );
  AND U18228 ( .A(p_input[4532]), .B(p_input[34532]), .Z(n12151) );
  AND U18229 ( .A(n12153), .B(n12154), .Z(o[4531]) );
  AND U18230 ( .A(p_input[24531]), .B(p_input[14531]), .Z(n12154) );
  AND U18231 ( .A(p_input[4531]), .B(p_input[34531]), .Z(n12153) );
  AND U18232 ( .A(n12155), .B(n12156), .Z(o[4530]) );
  AND U18233 ( .A(p_input[24530]), .B(p_input[14530]), .Z(n12156) );
  AND U18234 ( .A(p_input[4530]), .B(p_input[34530]), .Z(n12155) );
  AND U18235 ( .A(n12157), .B(n12158), .Z(o[452]) );
  AND U18236 ( .A(p_input[20452]), .B(p_input[10452]), .Z(n12158) );
  AND U18237 ( .A(p_input[452]), .B(p_input[30452]), .Z(n12157) );
  AND U18238 ( .A(n12159), .B(n12160), .Z(o[4529]) );
  AND U18239 ( .A(p_input[24529]), .B(p_input[14529]), .Z(n12160) );
  AND U18240 ( .A(p_input[4529]), .B(p_input[34529]), .Z(n12159) );
  AND U18241 ( .A(n12161), .B(n12162), .Z(o[4528]) );
  AND U18242 ( .A(p_input[24528]), .B(p_input[14528]), .Z(n12162) );
  AND U18243 ( .A(p_input[4528]), .B(p_input[34528]), .Z(n12161) );
  AND U18244 ( .A(n12163), .B(n12164), .Z(o[4527]) );
  AND U18245 ( .A(p_input[24527]), .B(p_input[14527]), .Z(n12164) );
  AND U18246 ( .A(p_input[4527]), .B(p_input[34527]), .Z(n12163) );
  AND U18247 ( .A(n12165), .B(n12166), .Z(o[4526]) );
  AND U18248 ( .A(p_input[24526]), .B(p_input[14526]), .Z(n12166) );
  AND U18249 ( .A(p_input[4526]), .B(p_input[34526]), .Z(n12165) );
  AND U18250 ( .A(n12167), .B(n12168), .Z(o[4525]) );
  AND U18251 ( .A(p_input[24525]), .B(p_input[14525]), .Z(n12168) );
  AND U18252 ( .A(p_input[4525]), .B(p_input[34525]), .Z(n12167) );
  AND U18253 ( .A(n12169), .B(n12170), .Z(o[4524]) );
  AND U18254 ( .A(p_input[24524]), .B(p_input[14524]), .Z(n12170) );
  AND U18255 ( .A(p_input[4524]), .B(p_input[34524]), .Z(n12169) );
  AND U18256 ( .A(n12171), .B(n12172), .Z(o[4523]) );
  AND U18257 ( .A(p_input[24523]), .B(p_input[14523]), .Z(n12172) );
  AND U18258 ( .A(p_input[4523]), .B(p_input[34523]), .Z(n12171) );
  AND U18259 ( .A(n12173), .B(n12174), .Z(o[4522]) );
  AND U18260 ( .A(p_input[24522]), .B(p_input[14522]), .Z(n12174) );
  AND U18261 ( .A(p_input[4522]), .B(p_input[34522]), .Z(n12173) );
  AND U18262 ( .A(n12175), .B(n12176), .Z(o[4521]) );
  AND U18263 ( .A(p_input[24521]), .B(p_input[14521]), .Z(n12176) );
  AND U18264 ( .A(p_input[4521]), .B(p_input[34521]), .Z(n12175) );
  AND U18265 ( .A(n12177), .B(n12178), .Z(o[4520]) );
  AND U18266 ( .A(p_input[24520]), .B(p_input[14520]), .Z(n12178) );
  AND U18267 ( .A(p_input[4520]), .B(p_input[34520]), .Z(n12177) );
  AND U18268 ( .A(n12179), .B(n12180), .Z(o[451]) );
  AND U18269 ( .A(p_input[20451]), .B(p_input[10451]), .Z(n12180) );
  AND U18270 ( .A(p_input[451]), .B(p_input[30451]), .Z(n12179) );
  AND U18271 ( .A(n12181), .B(n12182), .Z(o[4519]) );
  AND U18272 ( .A(p_input[24519]), .B(p_input[14519]), .Z(n12182) );
  AND U18273 ( .A(p_input[4519]), .B(p_input[34519]), .Z(n12181) );
  AND U18274 ( .A(n12183), .B(n12184), .Z(o[4518]) );
  AND U18275 ( .A(p_input[24518]), .B(p_input[14518]), .Z(n12184) );
  AND U18276 ( .A(p_input[4518]), .B(p_input[34518]), .Z(n12183) );
  AND U18277 ( .A(n12185), .B(n12186), .Z(o[4517]) );
  AND U18278 ( .A(p_input[24517]), .B(p_input[14517]), .Z(n12186) );
  AND U18279 ( .A(p_input[4517]), .B(p_input[34517]), .Z(n12185) );
  AND U18280 ( .A(n12187), .B(n12188), .Z(o[4516]) );
  AND U18281 ( .A(p_input[24516]), .B(p_input[14516]), .Z(n12188) );
  AND U18282 ( .A(p_input[4516]), .B(p_input[34516]), .Z(n12187) );
  AND U18283 ( .A(n12189), .B(n12190), .Z(o[4515]) );
  AND U18284 ( .A(p_input[24515]), .B(p_input[14515]), .Z(n12190) );
  AND U18285 ( .A(p_input[4515]), .B(p_input[34515]), .Z(n12189) );
  AND U18286 ( .A(n12191), .B(n12192), .Z(o[4514]) );
  AND U18287 ( .A(p_input[24514]), .B(p_input[14514]), .Z(n12192) );
  AND U18288 ( .A(p_input[4514]), .B(p_input[34514]), .Z(n12191) );
  AND U18289 ( .A(n12193), .B(n12194), .Z(o[4513]) );
  AND U18290 ( .A(p_input[24513]), .B(p_input[14513]), .Z(n12194) );
  AND U18291 ( .A(p_input[4513]), .B(p_input[34513]), .Z(n12193) );
  AND U18292 ( .A(n12195), .B(n12196), .Z(o[4512]) );
  AND U18293 ( .A(p_input[24512]), .B(p_input[14512]), .Z(n12196) );
  AND U18294 ( .A(p_input[4512]), .B(p_input[34512]), .Z(n12195) );
  AND U18295 ( .A(n12197), .B(n12198), .Z(o[4511]) );
  AND U18296 ( .A(p_input[24511]), .B(p_input[14511]), .Z(n12198) );
  AND U18297 ( .A(p_input[4511]), .B(p_input[34511]), .Z(n12197) );
  AND U18298 ( .A(n12199), .B(n12200), .Z(o[4510]) );
  AND U18299 ( .A(p_input[24510]), .B(p_input[14510]), .Z(n12200) );
  AND U18300 ( .A(p_input[4510]), .B(p_input[34510]), .Z(n12199) );
  AND U18301 ( .A(n12201), .B(n12202), .Z(o[450]) );
  AND U18302 ( .A(p_input[20450]), .B(p_input[10450]), .Z(n12202) );
  AND U18303 ( .A(p_input[450]), .B(p_input[30450]), .Z(n12201) );
  AND U18304 ( .A(n12203), .B(n12204), .Z(o[4509]) );
  AND U18305 ( .A(p_input[24509]), .B(p_input[14509]), .Z(n12204) );
  AND U18306 ( .A(p_input[4509]), .B(p_input[34509]), .Z(n12203) );
  AND U18307 ( .A(n12205), .B(n12206), .Z(o[4508]) );
  AND U18308 ( .A(p_input[24508]), .B(p_input[14508]), .Z(n12206) );
  AND U18309 ( .A(p_input[4508]), .B(p_input[34508]), .Z(n12205) );
  AND U18310 ( .A(n12207), .B(n12208), .Z(o[4507]) );
  AND U18311 ( .A(p_input[24507]), .B(p_input[14507]), .Z(n12208) );
  AND U18312 ( .A(p_input[4507]), .B(p_input[34507]), .Z(n12207) );
  AND U18313 ( .A(n12209), .B(n12210), .Z(o[4506]) );
  AND U18314 ( .A(p_input[24506]), .B(p_input[14506]), .Z(n12210) );
  AND U18315 ( .A(p_input[4506]), .B(p_input[34506]), .Z(n12209) );
  AND U18316 ( .A(n12211), .B(n12212), .Z(o[4505]) );
  AND U18317 ( .A(p_input[24505]), .B(p_input[14505]), .Z(n12212) );
  AND U18318 ( .A(p_input[4505]), .B(p_input[34505]), .Z(n12211) );
  AND U18319 ( .A(n12213), .B(n12214), .Z(o[4504]) );
  AND U18320 ( .A(p_input[24504]), .B(p_input[14504]), .Z(n12214) );
  AND U18321 ( .A(p_input[4504]), .B(p_input[34504]), .Z(n12213) );
  AND U18322 ( .A(n12215), .B(n12216), .Z(o[4503]) );
  AND U18323 ( .A(p_input[24503]), .B(p_input[14503]), .Z(n12216) );
  AND U18324 ( .A(p_input[4503]), .B(p_input[34503]), .Z(n12215) );
  AND U18325 ( .A(n12217), .B(n12218), .Z(o[4502]) );
  AND U18326 ( .A(p_input[24502]), .B(p_input[14502]), .Z(n12218) );
  AND U18327 ( .A(p_input[4502]), .B(p_input[34502]), .Z(n12217) );
  AND U18328 ( .A(n12219), .B(n12220), .Z(o[4501]) );
  AND U18329 ( .A(p_input[24501]), .B(p_input[14501]), .Z(n12220) );
  AND U18330 ( .A(p_input[4501]), .B(p_input[34501]), .Z(n12219) );
  AND U18331 ( .A(n12221), .B(n12222), .Z(o[4500]) );
  AND U18332 ( .A(p_input[24500]), .B(p_input[14500]), .Z(n12222) );
  AND U18333 ( .A(p_input[4500]), .B(p_input[34500]), .Z(n12221) );
  AND U18334 ( .A(n12223), .B(n12224), .Z(o[44]) );
  AND U18335 ( .A(p_input[20044]), .B(p_input[10044]), .Z(n12224) );
  AND U18336 ( .A(p_input[44]), .B(p_input[30044]), .Z(n12223) );
  AND U18337 ( .A(n12225), .B(n12226), .Z(o[449]) );
  AND U18338 ( .A(p_input[20449]), .B(p_input[10449]), .Z(n12226) );
  AND U18339 ( .A(p_input[449]), .B(p_input[30449]), .Z(n12225) );
  AND U18340 ( .A(n12227), .B(n12228), .Z(o[4499]) );
  AND U18341 ( .A(p_input[24499]), .B(p_input[14499]), .Z(n12228) );
  AND U18342 ( .A(p_input[4499]), .B(p_input[34499]), .Z(n12227) );
  AND U18343 ( .A(n12229), .B(n12230), .Z(o[4498]) );
  AND U18344 ( .A(p_input[24498]), .B(p_input[14498]), .Z(n12230) );
  AND U18345 ( .A(p_input[4498]), .B(p_input[34498]), .Z(n12229) );
  AND U18346 ( .A(n12231), .B(n12232), .Z(o[4497]) );
  AND U18347 ( .A(p_input[24497]), .B(p_input[14497]), .Z(n12232) );
  AND U18348 ( .A(p_input[4497]), .B(p_input[34497]), .Z(n12231) );
  AND U18349 ( .A(n12233), .B(n12234), .Z(o[4496]) );
  AND U18350 ( .A(p_input[24496]), .B(p_input[14496]), .Z(n12234) );
  AND U18351 ( .A(p_input[4496]), .B(p_input[34496]), .Z(n12233) );
  AND U18352 ( .A(n12235), .B(n12236), .Z(o[4495]) );
  AND U18353 ( .A(p_input[24495]), .B(p_input[14495]), .Z(n12236) );
  AND U18354 ( .A(p_input[4495]), .B(p_input[34495]), .Z(n12235) );
  AND U18355 ( .A(n12237), .B(n12238), .Z(o[4494]) );
  AND U18356 ( .A(p_input[24494]), .B(p_input[14494]), .Z(n12238) );
  AND U18357 ( .A(p_input[4494]), .B(p_input[34494]), .Z(n12237) );
  AND U18358 ( .A(n12239), .B(n12240), .Z(o[4493]) );
  AND U18359 ( .A(p_input[24493]), .B(p_input[14493]), .Z(n12240) );
  AND U18360 ( .A(p_input[4493]), .B(p_input[34493]), .Z(n12239) );
  AND U18361 ( .A(n12241), .B(n12242), .Z(o[4492]) );
  AND U18362 ( .A(p_input[24492]), .B(p_input[14492]), .Z(n12242) );
  AND U18363 ( .A(p_input[4492]), .B(p_input[34492]), .Z(n12241) );
  AND U18364 ( .A(n12243), .B(n12244), .Z(o[4491]) );
  AND U18365 ( .A(p_input[24491]), .B(p_input[14491]), .Z(n12244) );
  AND U18366 ( .A(p_input[4491]), .B(p_input[34491]), .Z(n12243) );
  AND U18367 ( .A(n12245), .B(n12246), .Z(o[4490]) );
  AND U18368 ( .A(p_input[24490]), .B(p_input[14490]), .Z(n12246) );
  AND U18369 ( .A(p_input[4490]), .B(p_input[34490]), .Z(n12245) );
  AND U18370 ( .A(n12247), .B(n12248), .Z(o[448]) );
  AND U18371 ( .A(p_input[20448]), .B(p_input[10448]), .Z(n12248) );
  AND U18372 ( .A(p_input[448]), .B(p_input[30448]), .Z(n12247) );
  AND U18373 ( .A(n12249), .B(n12250), .Z(o[4489]) );
  AND U18374 ( .A(p_input[24489]), .B(p_input[14489]), .Z(n12250) );
  AND U18375 ( .A(p_input[4489]), .B(p_input[34489]), .Z(n12249) );
  AND U18376 ( .A(n12251), .B(n12252), .Z(o[4488]) );
  AND U18377 ( .A(p_input[24488]), .B(p_input[14488]), .Z(n12252) );
  AND U18378 ( .A(p_input[4488]), .B(p_input[34488]), .Z(n12251) );
  AND U18379 ( .A(n12253), .B(n12254), .Z(o[4487]) );
  AND U18380 ( .A(p_input[24487]), .B(p_input[14487]), .Z(n12254) );
  AND U18381 ( .A(p_input[4487]), .B(p_input[34487]), .Z(n12253) );
  AND U18382 ( .A(n12255), .B(n12256), .Z(o[4486]) );
  AND U18383 ( .A(p_input[24486]), .B(p_input[14486]), .Z(n12256) );
  AND U18384 ( .A(p_input[4486]), .B(p_input[34486]), .Z(n12255) );
  AND U18385 ( .A(n12257), .B(n12258), .Z(o[4485]) );
  AND U18386 ( .A(p_input[24485]), .B(p_input[14485]), .Z(n12258) );
  AND U18387 ( .A(p_input[4485]), .B(p_input[34485]), .Z(n12257) );
  AND U18388 ( .A(n12259), .B(n12260), .Z(o[4484]) );
  AND U18389 ( .A(p_input[24484]), .B(p_input[14484]), .Z(n12260) );
  AND U18390 ( .A(p_input[4484]), .B(p_input[34484]), .Z(n12259) );
  AND U18391 ( .A(n12261), .B(n12262), .Z(o[4483]) );
  AND U18392 ( .A(p_input[24483]), .B(p_input[14483]), .Z(n12262) );
  AND U18393 ( .A(p_input[4483]), .B(p_input[34483]), .Z(n12261) );
  AND U18394 ( .A(n12263), .B(n12264), .Z(o[4482]) );
  AND U18395 ( .A(p_input[24482]), .B(p_input[14482]), .Z(n12264) );
  AND U18396 ( .A(p_input[4482]), .B(p_input[34482]), .Z(n12263) );
  AND U18397 ( .A(n12265), .B(n12266), .Z(o[4481]) );
  AND U18398 ( .A(p_input[24481]), .B(p_input[14481]), .Z(n12266) );
  AND U18399 ( .A(p_input[4481]), .B(p_input[34481]), .Z(n12265) );
  AND U18400 ( .A(n12267), .B(n12268), .Z(o[4480]) );
  AND U18401 ( .A(p_input[24480]), .B(p_input[14480]), .Z(n12268) );
  AND U18402 ( .A(p_input[4480]), .B(p_input[34480]), .Z(n12267) );
  AND U18403 ( .A(n12269), .B(n12270), .Z(o[447]) );
  AND U18404 ( .A(p_input[20447]), .B(p_input[10447]), .Z(n12270) );
  AND U18405 ( .A(p_input[447]), .B(p_input[30447]), .Z(n12269) );
  AND U18406 ( .A(n12271), .B(n12272), .Z(o[4479]) );
  AND U18407 ( .A(p_input[24479]), .B(p_input[14479]), .Z(n12272) );
  AND U18408 ( .A(p_input[4479]), .B(p_input[34479]), .Z(n12271) );
  AND U18409 ( .A(n12273), .B(n12274), .Z(o[4478]) );
  AND U18410 ( .A(p_input[24478]), .B(p_input[14478]), .Z(n12274) );
  AND U18411 ( .A(p_input[4478]), .B(p_input[34478]), .Z(n12273) );
  AND U18412 ( .A(n12275), .B(n12276), .Z(o[4477]) );
  AND U18413 ( .A(p_input[24477]), .B(p_input[14477]), .Z(n12276) );
  AND U18414 ( .A(p_input[4477]), .B(p_input[34477]), .Z(n12275) );
  AND U18415 ( .A(n12277), .B(n12278), .Z(o[4476]) );
  AND U18416 ( .A(p_input[24476]), .B(p_input[14476]), .Z(n12278) );
  AND U18417 ( .A(p_input[4476]), .B(p_input[34476]), .Z(n12277) );
  AND U18418 ( .A(n12279), .B(n12280), .Z(o[4475]) );
  AND U18419 ( .A(p_input[24475]), .B(p_input[14475]), .Z(n12280) );
  AND U18420 ( .A(p_input[4475]), .B(p_input[34475]), .Z(n12279) );
  AND U18421 ( .A(n12281), .B(n12282), .Z(o[4474]) );
  AND U18422 ( .A(p_input[24474]), .B(p_input[14474]), .Z(n12282) );
  AND U18423 ( .A(p_input[4474]), .B(p_input[34474]), .Z(n12281) );
  AND U18424 ( .A(n12283), .B(n12284), .Z(o[4473]) );
  AND U18425 ( .A(p_input[24473]), .B(p_input[14473]), .Z(n12284) );
  AND U18426 ( .A(p_input[4473]), .B(p_input[34473]), .Z(n12283) );
  AND U18427 ( .A(n12285), .B(n12286), .Z(o[4472]) );
  AND U18428 ( .A(p_input[24472]), .B(p_input[14472]), .Z(n12286) );
  AND U18429 ( .A(p_input[4472]), .B(p_input[34472]), .Z(n12285) );
  AND U18430 ( .A(n12287), .B(n12288), .Z(o[4471]) );
  AND U18431 ( .A(p_input[24471]), .B(p_input[14471]), .Z(n12288) );
  AND U18432 ( .A(p_input[4471]), .B(p_input[34471]), .Z(n12287) );
  AND U18433 ( .A(n12289), .B(n12290), .Z(o[4470]) );
  AND U18434 ( .A(p_input[24470]), .B(p_input[14470]), .Z(n12290) );
  AND U18435 ( .A(p_input[4470]), .B(p_input[34470]), .Z(n12289) );
  AND U18436 ( .A(n12291), .B(n12292), .Z(o[446]) );
  AND U18437 ( .A(p_input[20446]), .B(p_input[10446]), .Z(n12292) );
  AND U18438 ( .A(p_input[446]), .B(p_input[30446]), .Z(n12291) );
  AND U18439 ( .A(n12293), .B(n12294), .Z(o[4469]) );
  AND U18440 ( .A(p_input[24469]), .B(p_input[14469]), .Z(n12294) );
  AND U18441 ( .A(p_input[4469]), .B(p_input[34469]), .Z(n12293) );
  AND U18442 ( .A(n12295), .B(n12296), .Z(o[4468]) );
  AND U18443 ( .A(p_input[24468]), .B(p_input[14468]), .Z(n12296) );
  AND U18444 ( .A(p_input[4468]), .B(p_input[34468]), .Z(n12295) );
  AND U18445 ( .A(n12297), .B(n12298), .Z(o[4467]) );
  AND U18446 ( .A(p_input[24467]), .B(p_input[14467]), .Z(n12298) );
  AND U18447 ( .A(p_input[4467]), .B(p_input[34467]), .Z(n12297) );
  AND U18448 ( .A(n12299), .B(n12300), .Z(o[4466]) );
  AND U18449 ( .A(p_input[24466]), .B(p_input[14466]), .Z(n12300) );
  AND U18450 ( .A(p_input[4466]), .B(p_input[34466]), .Z(n12299) );
  AND U18451 ( .A(n12301), .B(n12302), .Z(o[4465]) );
  AND U18452 ( .A(p_input[24465]), .B(p_input[14465]), .Z(n12302) );
  AND U18453 ( .A(p_input[4465]), .B(p_input[34465]), .Z(n12301) );
  AND U18454 ( .A(n12303), .B(n12304), .Z(o[4464]) );
  AND U18455 ( .A(p_input[24464]), .B(p_input[14464]), .Z(n12304) );
  AND U18456 ( .A(p_input[4464]), .B(p_input[34464]), .Z(n12303) );
  AND U18457 ( .A(n12305), .B(n12306), .Z(o[4463]) );
  AND U18458 ( .A(p_input[24463]), .B(p_input[14463]), .Z(n12306) );
  AND U18459 ( .A(p_input[4463]), .B(p_input[34463]), .Z(n12305) );
  AND U18460 ( .A(n12307), .B(n12308), .Z(o[4462]) );
  AND U18461 ( .A(p_input[24462]), .B(p_input[14462]), .Z(n12308) );
  AND U18462 ( .A(p_input[4462]), .B(p_input[34462]), .Z(n12307) );
  AND U18463 ( .A(n12309), .B(n12310), .Z(o[4461]) );
  AND U18464 ( .A(p_input[24461]), .B(p_input[14461]), .Z(n12310) );
  AND U18465 ( .A(p_input[4461]), .B(p_input[34461]), .Z(n12309) );
  AND U18466 ( .A(n12311), .B(n12312), .Z(o[4460]) );
  AND U18467 ( .A(p_input[24460]), .B(p_input[14460]), .Z(n12312) );
  AND U18468 ( .A(p_input[4460]), .B(p_input[34460]), .Z(n12311) );
  AND U18469 ( .A(n12313), .B(n12314), .Z(o[445]) );
  AND U18470 ( .A(p_input[20445]), .B(p_input[10445]), .Z(n12314) );
  AND U18471 ( .A(p_input[445]), .B(p_input[30445]), .Z(n12313) );
  AND U18472 ( .A(n12315), .B(n12316), .Z(o[4459]) );
  AND U18473 ( .A(p_input[24459]), .B(p_input[14459]), .Z(n12316) );
  AND U18474 ( .A(p_input[4459]), .B(p_input[34459]), .Z(n12315) );
  AND U18475 ( .A(n12317), .B(n12318), .Z(o[4458]) );
  AND U18476 ( .A(p_input[24458]), .B(p_input[14458]), .Z(n12318) );
  AND U18477 ( .A(p_input[4458]), .B(p_input[34458]), .Z(n12317) );
  AND U18478 ( .A(n12319), .B(n12320), .Z(o[4457]) );
  AND U18479 ( .A(p_input[24457]), .B(p_input[14457]), .Z(n12320) );
  AND U18480 ( .A(p_input[4457]), .B(p_input[34457]), .Z(n12319) );
  AND U18481 ( .A(n12321), .B(n12322), .Z(o[4456]) );
  AND U18482 ( .A(p_input[24456]), .B(p_input[14456]), .Z(n12322) );
  AND U18483 ( .A(p_input[4456]), .B(p_input[34456]), .Z(n12321) );
  AND U18484 ( .A(n12323), .B(n12324), .Z(o[4455]) );
  AND U18485 ( .A(p_input[24455]), .B(p_input[14455]), .Z(n12324) );
  AND U18486 ( .A(p_input[4455]), .B(p_input[34455]), .Z(n12323) );
  AND U18487 ( .A(n12325), .B(n12326), .Z(o[4454]) );
  AND U18488 ( .A(p_input[24454]), .B(p_input[14454]), .Z(n12326) );
  AND U18489 ( .A(p_input[4454]), .B(p_input[34454]), .Z(n12325) );
  AND U18490 ( .A(n12327), .B(n12328), .Z(o[4453]) );
  AND U18491 ( .A(p_input[24453]), .B(p_input[14453]), .Z(n12328) );
  AND U18492 ( .A(p_input[4453]), .B(p_input[34453]), .Z(n12327) );
  AND U18493 ( .A(n12329), .B(n12330), .Z(o[4452]) );
  AND U18494 ( .A(p_input[24452]), .B(p_input[14452]), .Z(n12330) );
  AND U18495 ( .A(p_input[4452]), .B(p_input[34452]), .Z(n12329) );
  AND U18496 ( .A(n12331), .B(n12332), .Z(o[4451]) );
  AND U18497 ( .A(p_input[24451]), .B(p_input[14451]), .Z(n12332) );
  AND U18498 ( .A(p_input[4451]), .B(p_input[34451]), .Z(n12331) );
  AND U18499 ( .A(n12333), .B(n12334), .Z(o[4450]) );
  AND U18500 ( .A(p_input[24450]), .B(p_input[14450]), .Z(n12334) );
  AND U18501 ( .A(p_input[4450]), .B(p_input[34450]), .Z(n12333) );
  AND U18502 ( .A(n12335), .B(n12336), .Z(o[444]) );
  AND U18503 ( .A(p_input[20444]), .B(p_input[10444]), .Z(n12336) );
  AND U18504 ( .A(p_input[444]), .B(p_input[30444]), .Z(n12335) );
  AND U18505 ( .A(n12337), .B(n12338), .Z(o[4449]) );
  AND U18506 ( .A(p_input[24449]), .B(p_input[14449]), .Z(n12338) );
  AND U18507 ( .A(p_input[4449]), .B(p_input[34449]), .Z(n12337) );
  AND U18508 ( .A(n12339), .B(n12340), .Z(o[4448]) );
  AND U18509 ( .A(p_input[24448]), .B(p_input[14448]), .Z(n12340) );
  AND U18510 ( .A(p_input[4448]), .B(p_input[34448]), .Z(n12339) );
  AND U18511 ( .A(n12341), .B(n12342), .Z(o[4447]) );
  AND U18512 ( .A(p_input[24447]), .B(p_input[14447]), .Z(n12342) );
  AND U18513 ( .A(p_input[4447]), .B(p_input[34447]), .Z(n12341) );
  AND U18514 ( .A(n12343), .B(n12344), .Z(o[4446]) );
  AND U18515 ( .A(p_input[24446]), .B(p_input[14446]), .Z(n12344) );
  AND U18516 ( .A(p_input[4446]), .B(p_input[34446]), .Z(n12343) );
  AND U18517 ( .A(n12345), .B(n12346), .Z(o[4445]) );
  AND U18518 ( .A(p_input[24445]), .B(p_input[14445]), .Z(n12346) );
  AND U18519 ( .A(p_input[4445]), .B(p_input[34445]), .Z(n12345) );
  AND U18520 ( .A(n12347), .B(n12348), .Z(o[4444]) );
  AND U18521 ( .A(p_input[24444]), .B(p_input[14444]), .Z(n12348) );
  AND U18522 ( .A(p_input[4444]), .B(p_input[34444]), .Z(n12347) );
  AND U18523 ( .A(n12349), .B(n12350), .Z(o[4443]) );
  AND U18524 ( .A(p_input[24443]), .B(p_input[14443]), .Z(n12350) );
  AND U18525 ( .A(p_input[4443]), .B(p_input[34443]), .Z(n12349) );
  AND U18526 ( .A(n12351), .B(n12352), .Z(o[4442]) );
  AND U18527 ( .A(p_input[24442]), .B(p_input[14442]), .Z(n12352) );
  AND U18528 ( .A(p_input[4442]), .B(p_input[34442]), .Z(n12351) );
  AND U18529 ( .A(n12353), .B(n12354), .Z(o[4441]) );
  AND U18530 ( .A(p_input[24441]), .B(p_input[14441]), .Z(n12354) );
  AND U18531 ( .A(p_input[4441]), .B(p_input[34441]), .Z(n12353) );
  AND U18532 ( .A(n12355), .B(n12356), .Z(o[4440]) );
  AND U18533 ( .A(p_input[24440]), .B(p_input[14440]), .Z(n12356) );
  AND U18534 ( .A(p_input[4440]), .B(p_input[34440]), .Z(n12355) );
  AND U18535 ( .A(n12357), .B(n12358), .Z(o[443]) );
  AND U18536 ( .A(p_input[20443]), .B(p_input[10443]), .Z(n12358) );
  AND U18537 ( .A(p_input[443]), .B(p_input[30443]), .Z(n12357) );
  AND U18538 ( .A(n12359), .B(n12360), .Z(o[4439]) );
  AND U18539 ( .A(p_input[24439]), .B(p_input[14439]), .Z(n12360) );
  AND U18540 ( .A(p_input[4439]), .B(p_input[34439]), .Z(n12359) );
  AND U18541 ( .A(n12361), .B(n12362), .Z(o[4438]) );
  AND U18542 ( .A(p_input[24438]), .B(p_input[14438]), .Z(n12362) );
  AND U18543 ( .A(p_input[4438]), .B(p_input[34438]), .Z(n12361) );
  AND U18544 ( .A(n12363), .B(n12364), .Z(o[4437]) );
  AND U18545 ( .A(p_input[24437]), .B(p_input[14437]), .Z(n12364) );
  AND U18546 ( .A(p_input[4437]), .B(p_input[34437]), .Z(n12363) );
  AND U18547 ( .A(n12365), .B(n12366), .Z(o[4436]) );
  AND U18548 ( .A(p_input[24436]), .B(p_input[14436]), .Z(n12366) );
  AND U18549 ( .A(p_input[4436]), .B(p_input[34436]), .Z(n12365) );
  AND U18550 ( .A(n12367), .B(n12368), .Z(o[4435]) );
  AND U18551 ( .A(p_input[24435]), .B(p_input[14435]), .Z(n12368) );
  AND U18552 ( .A(p_input[4435]), .B(p_input[34435]), .Z(n12367) );
  AND U18553 ( .A(n12369), .B(n12370), .Z(o[4434]) );
  AND U18554 ( .A(p_input[24434]), .B(p_input[14434]), .Z(n12370) );
  AND U18555 ( .A(p_input[4434]), .B(p_input[34434]), .Z(n12369) );
  AND U18556 ( .A(n12371), .B(n12372), .Z(o[4433]) );
  AND U18557 ( .A(p_input[24433]), .B(p_input[14433]), .Z(n12372) );
  AND U18558 ( .A(p_input[4433]), .B(p_input[34433]), .Z(n12371) );
  AND U18559 ( .A(n12373), .B(n12374), .Z(o[4432]) );
  AND U18560 ( .A(p_input[24432]), .B(p_input[14432]), .Z(n12374) );
  AND U18561 ( .A(p_input[4432]), .B(p_input[34432]), .Z(n12373) );
  AND U18562 ( .A(n12375), .B(n12376), .Z(o[4431]) );
  AND U18563 ( .A(p_input[24431]), .B(p_input[14431]), .Z(n12376) );
  AND U18564 ( .A(p_input[4431]), .B(p_input[34431]), .Z(n12375) );
  AND U18565 ( .A(n12377), .B(n12378), .Z(o[4430]) );
  AND U18566 ( .A(p_input[24430]), .B(p_input[14430]), .Z(n12378) );
  AND U18567 ( .A(p_input[4430]), .B(p_input[34430]), .Z(n12377) );
  AND U18568 ( .A(n12379), .B(n12380), .Z(o[442]) );
  AND U18569 ( .A(p_input[20442]), .B(p_input[10442]), .Z(n12380) );
  AND U18570 ( .A(p_input[442]), .B(p_input[30442]), .Z(n12379) );
  AND U18571 ( .A(n12381), .B(n12382), .Z(o[4429]) );
  AND U18572 ( .A(p_input[24429]), .B(p_input[14429]), .Z(n12382) );
  AND U18573 ( .A(p_input[4429]), .B(p_input[34429]), .Z(n12381) );
  AND U18574 ( .A(n12383), .B(n12384), .Z(o[4428]) );
  AND U18575 ( .A(p_input[24428]), .B(p_input[14428]), .Z(n12384) );
  AND U18576 ( .A(p_input[4428]), .B(p_input[34428]), .Z(n12383) );
  AND U18577 ( .A(n12385), .B(n12386), .Z(o[4427]) );
  AND U18578 ( .A(p_input[24427]), .B(p_input[14427]), .Z(n12386) );
  AND U18579 ( .A(p_input[4427]), .B(p_input[34427]), .Z(n12385) );
  AND U18580 ( .A(n12387), .B(n12388), .Z(o[4426]) );
  AND U18581 ( .A(p_input[24426]), .B(p_input[14426]), .Z(n12388) );
  AND U18582 ( .A(p_input[4426]), .B(p_input[34426]), .Z(n12387) );
  AND U18583 ( .A(n12389), .B(n12390), .Z(o[4425]) );
  AND U18584 ( .A(p_input[24425]), .B(p_input[14425]), .Z(n12390) );
  AND U18585 ( .A(p_input[4425]), .B(p_input[34425]), .Z(n12389) );
  AND U18586 ( .A(n12391), .B(n12392), .Z(o[4424]) );
  AND U18587 ( .A(p_input[24424]), .B(p_input[14424]), .Z(n12392) );
  AND U18588 ( .A(p_input[4424]), .B(p_input[34424]), .Z(n12391) );
  AND U18589 ( .A(n12393), .B(n12394), .Z(o[4423]) );
  AND U18590 ( .A(p_input[24423]), .B(p_input[14423]), .Z(n12394) );
  AND U18591 ( .A(p_input[4423]), .B(p_input[34423]), .Z(n12393) );
  AND U18592 ( .A(n12395), .B(n12396), .Z(o[4422]) );
  AND U18593 ( .A(p_input[24422]), .B(p_input[14422]), .Z(n12396) );
  AND U18594 ( .A(p_input[4422]), .B(p_input[34422]), .Z(n12395) );
  AND U18595 ( .A(n12397), .B(n12398), .Z(o[4421]) );
  AND U18596 ( .A(p_input[24421]), .B(p_input[14421]), .Z(n12398) );
  AND U18597 ( .A(p_input[4421]), .B(p_input[34421]), .Z(n12397) );
  AND U18598 ( .A(n12399), .B(n12400), .Z(o[4420]) );
  AND U18599 ( .A(p_input[24420]), .B(p_input[14420]), .Z(n12400) );
  AND U18600 ( .A(p_input[4420]), .B(p_input[34420]), .Z(n12399) );
  AND U18601 ( .A(n12401), .B(n12402), .Z(o[441]) );
  AND U18602 ( .A(p_input[20441]), .B(p_input[10441]), .Z(n12402) );
  AND U18603 ( .A(p_input[441]), .B(p_input[30441]), .Z(n12401) );
  AND U18604 ( .A(n12403), .B(n12404), .Z(o[4419]) );
  AND U18605 ( .A(p_input[24419]), .B(p_input[14419]), .Z(n12404) );
  AND U18606 ( .A(p_input[4419]), .B(p_input[34419]), .Z(n12403) );
  AND U18607 ( .A(n12405), .B(n12406), .Z(o[4418]) );
  AND U18608 ( .A(p_input[24418]), .B(p_input[14418]), .Z(n12406) );
  AND U18609 ( .A(p_input[4418]), .B(p_input[34418]), .Z(n12405) );
  AND U18610 ( .A(n12407), .B(n12408), .Z(o[4417]) );
  AND U18611 ( .A(p_input[24417]), .B(p_input[14417]), .Z(n12408) );
  AND U18612 ( .A(p_input[4417]), .B(p_input[34417]), .Z(n12407) );
  AND U18613 ( .A(n12409), .B(n12410), .Z(o[4416]) );
  AND U18614 ( .A(p_input[24416]), .B(p_input[14416]), .Z(n12410) );
  AND U18615 ( .A(p_input[4416]), .B(p_input[34416]), .Z(n12409) );
  AND U18616 ( .A(n12411), .B(n12412), .Z(o[4415]) );
  AND U18617 ( .A(p_input[24415]), .B(p_input[14415]), .Z(n12412) );
  AND U18618 ( .A(p_input[4415]), .B(p_input[34415]), .Z(n12411) );
  AND U18619 ( .A(n12413), .B(n12414), .Z(o[4414]) );
  AND U18620 ( .A(p_input[24414]), .B(p_input[14414]), .Z(n12414) );
  AND U18621 ( .A(p_input[4414]), .B(p_input[34414]), .Z(n12413) );
  AND U18622 ( .A(n12415), .B(n12416), .Z(o[4413]) );
  AND U18623 ( .A(p_input[24413]), .B(p_input[14413]), .Z(n12416) );
  AND U18624 ( .A(p_input[4413]), .B(p_input[34413]), .Z(n12415) );
  AND U18625 ( .A(n12417), .B(n12418), .Z(o[4412]) );
  AND U18626 ( .A(p_input[24412]), .B(p_input[14412]), .Z(n12418) );
  AND U18627 ( .A(p_input[4412]), .B(p_input[34412]), .Z(n12417) );
  AND U18628 ( .A(n12419), .B(n12420), .Z(o[4411]) );
  AND U18629 ( .A(p_input[24411]), .B(p_input[14411]), .Z(n12420) );
  AND U18630 ( .A(p_input[4411]), .B(p_input[34411]), .Z(n12419) );
  AND U18631 ( .A(n12421), .B(n12422), .Z(o[4410]) );
  AND U18632 ( .A(p_input[24410]), .B(p_input[14410]), .Z(n12422) );
  AND U18633 ( .A(p_input[4410]), .B(p_input[34410]), .Z(n12421) );
  AND U18634 ( .A(n12423), .B(n12424), .Z(o[440]) );
  AND U18635 ( .A(p_input[20440]), .B(p_input[10440]), .Z(n12424) );
  AND U18636 ( .A(p_input[440]), .B(p_input[30440]), .Z(n12423) );
  AND U18637 ( .A(n12425), .B(n12426), .Z(o[4409]) );
  AND U18638 ( .A(p_input[24409]), .B(p_input[14409]), .Z(n12426) );
  AND U18639 ( .A(p_input[4409]), .B(p_input[34409]), .Z(n12425) );
  AND U18640 ( .A(n12427), .B(n12428), .Z(o[4408]) );
  AND U18641 ( .A(p_input[24408]), .B(p_input[14408]), .Z(n12428) );
  AND U18642 ( .A(p_input[4408]), .B(p_input[34408]), .Z(n12427) );
  AND U18643 ( .A(n12429), .B(n12430), .Z(o[4407]) );
  AND U18644 ( .A(p_input[24407]), .B(p_input[14407]), .Z(n12430) );
  AND U18645 ( .A(p_input[4407]), .B(p_input[34407]), .Z(n12429) );
  AND U18646 ( .A(n12431), .B(n12432), .Z(o[4406]) );
  AND U18647 ( .A(p_input[24406]), .B(p_input[14406]), .Z(n12432) );
  AND U18648 ( .A(p_input[4406]), .B(p_input[34406]), .Z(n12431) );
  AND U18649 ( .A(n12433), .B(n12434), .Z(o[4405]) );
  AND U18650 ( .A(p_input[24405]), .B(p_input[14405]), .Z(n12434) );
  AND U18651 ( .A(p_input[4405]), .B(p_input[34405]), .Z(n12433) );
  AND U18652 ( .A(n12435), .B(n12436), .Z(o[4404]) );
  AND U18653 ( .A(p_input[24404]), .B(p_input[14404]), .Z(n12436) );
  AND U18654 ( .A(p_input[4404]), .B(p_input[34404]), .Z(n12435) );
  AND U18655 ( .A(n12437), .B(n12438), .Z(o[4403]) );
  AND U18656 ( .A(p_input[24403]), .B(p_input[14403]), .Z(n12438) );
  AND U18657 ( .A(p_input[4403]), .B(p_input[34403]), .Z(n12437) );
  AND U18658 ( .A(n12439), .B(n12440), .Z(o[4402]) );
  AND U18659 ( .A(p_input[24402]), .B(p_input[14402]), .Z(n12440) );
  AND U18660 ( .A(p_input[4402]), .B(p_input[34402]), .Z(n12439) );
  AND U18661 ( .A(n12441), .B(n12442), .Z(o[4401]) );
  AND U18662 ( .A(p_input[24401]), .B(p_input[14401]), .Z(n12442) );
  AND U18663 ( .A(p_input[4401]), .B(p_input[34401]), .Z(n12441) );
  AND U18664 ( .A(n12443), .B(n12444), .Z(o[4400]) );
  AND U18665 ( .A(p_input[24400]), .B(p_input[14400]), .Z(n12444) );
  AND U18666 ( .A(p_input[4400]), .B(p_input[34400]), .Z(n12443) );
  AND U18667 ( .A(n12445), .B(n12446), .Z(o[43]) );
  AND U18668 ( .A(p_input[20043]), .B(p_input[10043]), .Z(n12446) );
  AND U18669 ( .A(p_input[43]), .B(p_input[30043]), .Z(n12445) );
  AND U18670 ( .A(n12447), .B(n12448), .Z(o[439]) );
  AND U18671 ( .A(p_input[20439]), .B(p_input[10439]), .Z(n12448) );
  AND U18672 ( .A(p_input[439]), .B(p_input[30439]), .Z(n12447) );
  AND U18673 ( .A(n12449), .B(n12450), .Z(o[4399]) );
  AND U18674 ( .A(p_input[24399]), .B(p_input[14399]), .Z(n12450) );
  AND U18675 ( .A(p_input[4399]), .B(p_input[34399]), .Z(n12449) );
  AND U18676 ( .A(n12451), .B(n12452), .Z(o[4398]) );
  AND U18677 ( .A(p_input[24398]), .B(p_input[14398]), .Z(n12452) );
  AND U18678 ( .A(p_input[4398]), .B(p_input[34398]), .Z(n12451) );
  AND U18679 ( .A(n12453), .B(n12454), .Z(o[4397]) );
  AND U18680 ( .A(p_input[24397]), .B(p_input[14397]), .Z(n12454) );
  AND U18681 ( .A(p_input[4397]), .B(p_input[34397]), .Z(n12453) );
  AND U18682 ( .A(n12455), .B(n12456), .Z(o[4396]) );
  AND U18683 ( .A(p_input[24396]), .B(p_input[14396]), .Z(n12456) );
  AND U18684 ( .A(p_input[4396]), .B(p_input[34396]), .Z(n12455) );
  AND U18685 ( .A(n12457), .B(n12458), .Z(o[4395]) );
  AND U18686 ( .A(p_input[24395]), .B(p_input[14395]), .Z(n12458) );
  AND U18687 ( .A(p_input[4395]), .B(p_input[34395]), .Z(n12457) );
  AND U18688 ( .A(n12459), .B(n12460), .Z(o[4394]) );
  AND U18689 ( .A(p_input[24394]), .B(p_input[14394]), .Z(n12460) );
  AND U18690 ( .A(p_input[4394]), .B(p_input[34394]), .Z(n12459) );
  AND U18691 ( .A(n12461), .B(n12462), .Z(o[4393]) );
  AND U18692 ( .A(p_input[24393]), .B(p_input[14393]), .Z(n12462) );
  AND U18693 ( .A(p_input[4393]), .B(p_input[34393]), .Z(n12461) );
  AND U18694 ( .A(n12463), .B(n12464), .Z(o[4392]) );
  AND U18695 ( .A(p_input[24392]), .B(p_input[14392]), .Z(n12464) );
  AND U18696 ( .A(p_input[4392]), .B(p_input[34392]), .Z(n12463) );
  AND U18697 ( .A(n12465), .B(n12466), .Z(o[4391]) );
  AND U18698 ( .A(p_input[24391]), .B(p_input[14391]), .Z(n12466) );
  AND U18699 ( .A(p_input[4391]), .B(p_input[34391]), .Z(n12465) );
  AND U18700 ( .A(n12467), .B(n12468), .Z(o[4390]) );
  AND U18701 ( .A(p_input[24390]), .B(p_input[14390]), .Z(n12468) );
  AND U18702 ( .A(p_input[4390]), .B(p_input[34390]), .Z(n12467) );
  AND U18703 ( .A(n12469), .B(n12470), .Z(o[438]) );
  AND U18704 ( .A(p_input[20438]), .B(p_input[10438]), .Z(n12470) );
  AND U18705 ( .A(p_input[438]), .B(p_input[30438]), .Z(n12469) );
  AND U18706 ( .A(n12471), .B(n12472), .Z(o[4389]) );
  AND U18707 ( .A(p_input[24389]), .B(p_input[14389]), .Z(n12472) );
  AND U18708 ( .A(p_input[4389]), .B(p_input[34389]), .Z(n12471) );
  AND U18709 ( .A(n12473), .B(n12474), .Z(o[4388]) );
  AND U18710 ( .A(p_input[24388]), .B(p_input[14388]), .Z(n12474) );
  AND U18711 ( .A(p_input[4388]), .B(p_input[34388]), .Z(n12473) );
  AND U18712 ( .A(n12475), .B(n12476), .Z(o[4387]) );
  AND U18713 ( .A(p_input[24387]), .B(p_input[14387]), .Z(n12476) );
  AND U18714 ( .A(p_input[4387]), .B(p_input[34387]), .Z(n12475) );
  AND U18715 ( .A(n12477), .B(n12478), .Z(o[4386]) );
  AND U18716 ( .A(p_input[24386]), .B(p_input[14386]), .Z(n12478) );
  AND U18717 ( .A(p_input[4386]), .B(p_input[34386]), .Z(n12477) );
  AND U18718 ( .A(n12479), .B(n12480), .Z(o[4385]) );
  AND U18719 ( .A(p_input[24385]), .B(p_input[14385]), .Z(n12480) );
  AND U18720 ( .A(p_input[4385]), .B(p_input[34385]), .Z(n12479) );
  AND U18721 ( .A(n12481), .B(n12482), .Z(o[4384]) );
  AND U18722 ( .A(p_input[24384]), .B(p_input[14384]), .Z(n12482) );
  AND U18723 ( .A(p_input[4384]), .B(p_input[34384]), .Z(n12481) );
  AND U18724 ( .A(n12483), .B(n12484), .Z(o[4383]) );
  AND U18725 ( .A(p_input[24383]), .B(p_input[14383]), .Z(n12484) );
  AND U18726 ( .A(p_input[4383]), .B(p_input[34383]), .Z(n12483) );
  AND U18727 ( .A(n12485), .B(n12486), .Z(o[4382]) );
  AND U18728 ( .A(p_input[24382]), .B(p_input[14382]), .Z(n12486) );
  AND U18729 ( .A(p_input[4382]), .B(p_input[34382]), .Z(n12485) );
  AND U18730 ( .A(n12487), .B(n12488), .Z(o[4381]) );
  AND U18731 ( .A(p_input[24381]), .B(p_input[14381]), .Z(n12488) );
  AND U18732 ( .A(p_input[4381]), .B(p_input[34381]), .Z(n12487) );
  AND U18733 ( .A(n12489), .B(n12490), .Z(o[4380]) );
  AND U18734 ( .A(p_input[24380]), .B(p_input[14380]), .Z(n12490) );
  AND U18735 ( .A(p_input[4380]), .B(p_input[34380]), .Z(n12489) );
  AND U18736 ( .A(n12491), .B(n12492), .Z(o[437]) );
  AND U18737 ( .A(p_input[20437]), .B(p_input[10437]), .Z(n12492) );
  AND U18738 ( .A(p_input[437]), .B(p_input[30437]), .Z(n12491) );
  AND U18739 ( .A(n12493), .B(n12494), .Z(o[4379]) );
  AND U18740 ( .A(p_input[24379]), .B(p_input[14379]), .Z(n12494) );
  AND U18741 ( .A(p_input[4379]), .B(p_input[34379]), .Z(n12493) );
  AND U18742 ( .A(n12495), .B(n12496), .Z(o[4378]) );
  AND U18743 ( .A(p_input[24378]), .B(p_input[14378]), .Z(n12496) );
  AND U18744 ( .A(p_input[4378]), .B(p_input[34378]), .Z(n12495) );
  AND U18745 ( .A(n12497), .B(n12498), .Z(o[4377]) );
  AND U18746 ( .A(p_input[24377]), .B(p_input[14377]), .Z(n12498) );
  AND U18747 ( .A(p_input[4377]), .B(p_input[34377]), .Z(n12497) );
  AND U18748 ( .A(n12499), .B(n12500), .Z(o[4376]) );
  AND U18749 ( .A(p_input[24376]), .B(p_input[14376]), .Z(n12500) );
  AND U18750 ( .A(p_input[4376]), .B(p_input[34376]), .Z(n12499) );
  AND U18751 ( .A(n12501), .B(n12502), .Z(o[4375]) );
  AND U18752 ( .A(p_input[24375]), .B(p_input[14375]), .Z(n12502) );
  AND U18753 ( .A(p_input[4375]), .B(p_input[34375]), .Z(n12501) );
  AND U18754 ( .A(n12503), .B(n12504), .Z(o[4374]) );
  AND U18755 ( .A(p_input[24374]), .B(p_input[14374]), .Z(n12504) );
  AND U18756 ( .A(p_input[4374]), .B(p_input[34374]), .Z(n12503) );
  AND U18757 ( .A(n12505), .B(n12506), .Z(o[4373]) );
  AND U18758 ( .A(p_input[24373]), .B(p_input[14373]), .Z(n12506) );
  AND U18759 ( .A(p_input[4373]), .B(p_input[34373]), .Z(n12505) );
  AND U18760 ( .A(n12507), .B(n12508), .Z(o[4372]) );
  AND U18761 ( .A(p_input[24372]), .B(p_input[14372]), .Z(n12508) );
  AND U18762 ( .A(p_input[4372]), .B(p_input[34372]), .Z(n12507) );
  AND U18763 ( .A(n12509), .B(n12510), .Z(o[4371]) );
  AND U18764 ( .A(p_input[24371]), .B(p_input[14371]), .Z(n12510) );
  AND U18765 ( .A(p_input[4371]), .B(p_input[34371]), .Z(n12509) );
  AND U18766 ( .A(n12511), .B(n12512), .Z(o[4370]) );
  AND U18767 ( .A(p_input[24370]), .B(p_input[14370]), .Z(n12512) );
  AND U18768 ( .A(p_input[4370]), .B(p_input[34370]), .Z(n12511) );
  AND U18769 ( .A(n12513), .B(n12514), .Z(o[436]) );
  AND U18770 ( .A(p_input[20436]), .B(p_input[10436]), .Z(n12514) );
  AND U18771 ( .A(p_input[436]), .B(p_input[30436]), .Z(n12513) );
  AND U18772 ( .A(n12515), .B(n12516), .Z(o[4369]) );
  AND U18773 ( .A(p_input[24369]), .B(p_input[14369]), .Z(n12516) );
  AND U18774 ( .A(p_input[4369]), .B(p_input[34369]), .Z(n12515) );
  AND U18775 ( .A(n12517), .B(n12518), .Z(o[4368]) );
  AND U18776 ( .A(p_input[24368]), .B(p_input[14368]), .Z(n12518) );
  AND U18777 ( .A(p_input[4368]), .B(p_input[34368]), .Z(n12517) );
  AND U18778 ( .A(n12519), .B(n12520), .Z(o[4367]) );
  AND U18779 ( .A(p_input[24367]), .B(p_input[14367]), .Z(n12520) );
  AND U18780 ( .A(p_input[4367]), .B(p_input[34367]), .Z(n12519) );
  AND U18781 ( .A(n12521), .B(n12522), .Z(o[4366]) );
  AND U18782 ( .A(p_input[24366]), .B(p_input[14366]), .Z(n12522) );
  AND U18783 ( .A(p_input[4366]), .B(p_input[34366]), .Z(n12521) );
  AND U18784 ( .A(n12523), .B(n12524), .Z(o[4365]) );
  AND U18785 ( .A(p_input[24365]), .B(p_input[14365]), .Z(n12524) );
  AND U18786 ( .A(p_input[4365]), .B(p_input[34365]), .Z(n12523) );
  AND U18787 ( .A(n12525), .B(n12526), .Z(o[4364]) );
  AND U18788 ( .A(p_input[24364]), .B(p_input[14364]), .Z(n12526) );
  AND U18789 ( .A(p_input[4364]), .B(p_input[34364]), .Z(n12525) );
  AND U18790 ( .A(n12527), .B(n12528), .Z(o[4363]) );
  AND U18791 ( .A(p_input[24363]), .B(p_input[14363]), .Z(n12528) );
  AND U18792 ( .A(p_input[4363]), .B(p_input[34363]), .Z(n12527) );
  AND U18793 ( .A(n12529), .B(n12530), .Z(o[4362]) );
  AND U18794 ( .A(p_input[24362]), .B(p_input[14362]), .Z(n12530) );
  AND U18795 ( .A(p_input[4362]), .B(p_input[34362]), .Z(n12529) );
  AND U18796 ( .A(n12531), .B(n12532), .Z(o[4361]) );
  AND U18797 ( .A(p_input[24361]), .B(p_input[14361]), .Z(n12532) );
  AND U18798 ( .A(p_input[4361]), .B(p_input[34361]), .Z(n12531) );
  AND U18799 ( .A(n12533), .B(n12534), .Z(o[4360]) );
  AND U18800 ( .A(p_input[24360]), .B(p_input[14360]), .Z(n12534) );
  AND U18801 ( .A(p_input[4360]), .B(p_input[34360]), .Z(n12533) );
  AND U18802 ( .A(n12535), .B(n12536), .Z(o[435]) );
  AND U18803 ( .A(p_input[20435]), .B(p_input[10435]), .Z(n12536) );
  AND U18804 ( .A(p_input[435]), .B(p_input[30435]), .Z(n12535) );
  AND U18805 ( .A(n12537), .B(n12538), .Z(o[4359]) );
  AND U18806 ( .A(p_input[24359]), .B(p_input[14359]), .Z(n12538) );
  AND U18807 ( .A(p_input[4359]), .B(p_input[34359]), .Z(n12537) );
  AND U18808 ( .A(n12539), .B(n12540), .Z(o[4358]) );
  AND U18809 ( .A(p_input[24358]), .B(p_input[14358]), .Z(n12540) );
  AND U18810 ( .A(p_input[4358]), .B(p_input[34358]), .Z(n12539) );
  AND U18811 ( .A(n12541), .B(n12542), .Z(o[4357]) );
  AND U18812 ( .A(p_input[24357]), .B(p_input[14357]), .Z(n12542) );
  AND U18813 ( .A(p_input[4357]), .B(p_input[34357]), .Z(n12541) );
  AND U18814 ( .A(n12543), .B(n12544), .Z(o[4356]) );
  AND U18815 ( .A(p_input[24356]), .B(p_input[14356]), .Z(n12544) );
  AND U18816 ( .A(p_input[4356]), .B(p_input[34356]), .Z(n12543) );
  AND U18817 ( .A(n12545), .B(n12546), .Z(o[4355]) );
  AND U18818 ( .A(p_input[24355]), .B(p_input[14355]), .Z(n12546) );
  AND U18819 ( .A(p_input[4355]), .B(p_input[34355]), .Z(n12545) );
  AND U18820 ( .A(n12547), .B(n12548), .Z(o[4354]) );
  AND U18821 ( .A(p_input[24354]), .B(p_input[14354]), .Z(n12548) );
  AND U18822 ( .A(p_input[4354]), .B(p_input[34354]), .Z(n12547) );
  AND U18823 ( .A(n12549), .B(n12550), .Z(o[4353]) );
  AND U18824 ( .A(p_input[24353]), .B(p_input[14353]), .Z(n12550) );
  AND U18825 ( .A(p_input[4353]), .B(p_input[34353]), .Z(n12549) );
  AND U18826 ( .A(n12551), .B(n12552), .Z(o[4352]) );
  AND U18827 ( .A(p_input[24352]), .B(p_input[14352]), .Z(n12552) );
  AND U18828 ( .A(p_input[4352]), .B(p_input[34352]), .Z(n12551) );
  AND U18829 ( .A(n12553), .B(n12554), .Z(o[4351]) );
  AND U18830 ( .A(p_input[24351]), .B(p_input[14351]), .Z(n12554) );
  AND U18831 ( .A(p_input[4351]), .B(p_input[34351]), .Z(n12553) );
  AND U18832 ( .A(n12555), .B(n12556), .Z(o[4350]) );
  AND U18833 ( .A(p_input[24350]), .B(p_input[14350]), .Z(n12556) );
  AND U18834 ( .A(p_input[4350]), .B(p_input[34350]), .Z(n12555) );
  AND U18835 ( .A(n12557), .B(n12558), .Z(o[434]) );
  AND U18836 ( .A(p_input[20434]), .B(p_input[10434]), .Z(n12558) );
  AND U18837 ( .A(p_input[434]), .B(p_input[30434]), .Z(n12557) );
  AND U18838 ( .A(n12559), .B(n12560), .Z(o[4349]) );
  AND U18839 ( .A(p_input[24349]), .B(p_input[14349]), .Z(n12560) );
  AND U18840 ( .A(p_input[4349]), .B(p_input[34349]), .Z(n12559) );
  AND U18841 ( .A(n12561), .B(n12562), .Z(o[4348]) );
  AND U18842 ( .A(p_input[24348]), .B(p_input[14348]), .Z(n12562) );
  AND U18843 ( .A(p_input[4348]), .B(p_input[34348]), .Z(n12561) );
  AND U18844 ( .A(n12563), .B(n12564), .Z(o[4347]) );
  AND U18845 ( .A(p_input[24347]), .B(p_input[14347]), .Z(n12564) );
  AND U18846 ( .A(p_input[4347]), .B(p_input[34347]), .Z(n12563) );
  AND U18847 ( .A(n12565), .B(n12566), .Z(o[4346]) );
  AND U18848 ( .A(p_input[24346]), .B(p_input[14346]), .Z(n12566) );
  AND U18849 ( .A(p_input[4346]), .B(p_input[34346]), .Z(n12565) );
  AND U18850 ( .A(n12567), .B(n12568), .Z(o[4345]) );
  AND U18851 ( .A(p_input[24345]), .B(p_input[14345]), .Z(n12568) );
  AND U18852 ( .A(p_input[4345]), .B(p_input[34345]), .Z(n12567) );
  AND U18853 ( .A(n12569), .B(n12570), .Z(o[4344]) );
  AND U18854 ( .A(p_input[24344]), .B(p_input[14344]), .Z(n12570) );
  AND U18855 ( .A(p_input[4344]), .B(p_input[34344]), .Z(n12569) );
  AND U18856 ( .A(n12571), .B(n12572), .Z(o[4343]) );
  AND U18857 ( .A(p_input[24343]), .B(p_input[14343]), .Z(n12572) );
  AND U18858 ( .A(p_input[4343]), .B(p_input[34343]), .Z(n12571) );
  AND U18859 ( .A(n12573), .B(n12574), .Z(o[4342]) );
  AND U18860 ( .A(p_input[24342]), .B(p_input[14342]), .Z(n12574) );
  AND U18861 ( .A(p_input[4342]), .B(p_input[34342]), .Z(n12573) );
  AND U18862 ( .A(n12575), .B(n12576), .Z(o[4341]) );
  AND U18863 ( .A(p_input[24341]), .B(p_input[14341]), .Z(n12576) );
  AND U18864 ( .A(p_input[4341]), .B(p_input[34341]), .Z(n12575) );
  AND U18865 ( .A(n12577), .B(n12578), .Z(o[4340]) );
  AND U18866 ( .A(p_input[24340]), .B(p_input[14340]), .Z(n12578) );
  AND U18867 ( .A(p_input[4340]), .B(p_input[34340]), .Z(n12577) );
  AND U18868 ( .A(n12579), .B(n12580), .Z(o[433]) );
  AND U18869 ( .A(p_input[20433]), .B(p_input[10433]), .Z(n12580) );
  AND U18870 ( .A(p_input[433]), .B(p_input[30433]), .Z(n12579) );
  AND U18871 ( .A(n12581), .B(n12582), .Z(o[4339]) );
  AND U18872 ( .A(p_input[24339]), .B(p_input[14339]), .Z(n12582) );
  AND U18873 ( .A(p_input[4339]), .B(p_input[34339]), .Z(n12581) );
  AND U18874 ( .A(n12583), .B(n12584), .Z(o[4338]) );
  AND U18875 ( .A(p_input[24338]), .B(p_input[14338]), .Z(n12584) );
  AND U18876 ( .A(p_input[4338]), .B(p_input[34338]), .Z(n12583) );
  AND U18877 ( .A(n12585), .B(n12586), .Z(o[4337]) );
  AND U18878 ( .A(p_input[24337]), .B(p_input[14337]), .Z(n12586) );
  AND U18879 ( .A(p_input[4337]), .B(p_input[34337]), .Z(n12585) );
  AND U18880 ( .A(n12587), .B(n12588), .Z(o[4336]) );
  AND U18881 ( .A(p_input[24336]), .B(p_input[14336]), .Z(n12588) );
  AND U18882 ( .A(p_input[4336]), .B(p_input[34336]), .Z(n12587) );
  AND U18883 ( .A(n12589), .B(n12590), .Z(o[4335]) );
  AND U18884 ( .A(p_input[24335]), .B(p_input[14335]), .Z(n12590) );
  AND U18885 ( .A(p_input[4335]), .B(p_input[34335]), .Z(n12589) );
  AND U18886 ( .A(n12591), .B(n12592), .Z(o[4334]) );
  AND U18887 ( .A(p_input[24334]), .B(p_input[14334]), .Z(n12592) );
  AND U18888 ( .A(p_input[4334]), .B(p_input[34334]), .Z(n12591) );
  AND U18889 ( .A(n12593), .B(n12594), .Z(o[4333]) );
  AND U18890 ( .A(p_input[24333]), .B(p_input[14333]), .Z(n12594) );
  AND U18891 ( .A(p_input[4333]), .B(p_input[34333]), .Z(n12593) );
  AND U18892 ( .A(n12595), .B(n12596), .Z(o[4332]) );
  AND U18893 ( .A(p_input[24332]), .B(p_input[14332]), .Z(n12596) );
  AND U18894 ( .A(p_input[4332]), .B(p_input[34332]), .Z(n12595) );
  AND U18895 ( .A(n12597), .B(n12598), .Z(o[4331]) );
  AND U18896 ( .A(p_input[24331]), .B(p_input[14331]), .Z(n12598) );
  AND U18897 ( .A(p_input[4331]), .B(p_input[34331]), .Z(n12597) );
  AND U18898 ( .A(n12599), .B(n12600), .Z(o[4330]) );
  AND U18899 ( .A(p_input[24330]), .B(p_input[14330]), .Z(n12600) );
  AND U18900 ( .A(p_input[4330]), .B(p_input[34330]), .Z(n12599) );
  AND U18901 ( .A(n12601), .B(n12602), .Z(o[432]) );
  AND U18902 ( .A(p_input[20432]), .B(p_input[10432]), .Z(n12602) );
  AND U18903 ( .A(p_input[432]), .B(p_input[30432]), .Z(n12601) );
  AND U18904 ( .A(n12603), .B(n12604), .Z(o[4329]) );
  AND U18905 ( .A(p_input[24329]), .B(p_input[14329]), .Z(n12604) );
  AND U18906 ( .A(p_input[4329]), .B(p_input[34329]), .Z(n12603) );
  AND U18907 ( .A(n12605), .B(n12606), .Z(o[4328]) );
  AND U18908 ( .A(p_input[24328]), .B(p_input[14328]), .Z(n12606) );
  AND U18909 ( .A(p_input[4328]), .B(p_input[34328]), .Z(n12605) );
  AND U18910 ( .A(n12607), .B(n12608), .Z(o[4327]) );
  AND U18911 ( .A(p_input[24327]), .B(p_input[14327]), .Z(n12608) );
  AND U18912 ( .A(p_input[4327]), .B(p_input[34327]), .Z(n12607) );
  AND U18913 ( .A(n12609), .B(n12610), .Z(o[4326]) );
  AND U18914 ( .A(p_input[24326]), .B(p_input[14326]), .Z(n12610) );
  AND U18915 ( .A(p_input[4326]), .B(p_input[34326]), .Z(n12609) );
  AND U18916 ( .A(n12611), .B(n12612), .Z(o[4325]) );
  AND U18917 ( .A(p_input[24325]), .B(p_input[14325]), .Z(n12612) );
  AND U18918 ( .A(p_input[4325]), .B(p_input[34325]), .Z(n12611) );
  AND U18919 ( .A(n12613), .B(n12614), .Z(o[4324]) );
  AND U18920 ( .A(p_input[24324]), .B(p_input[14324]), .Z(n12614) );
  AND U18921 ( .A(p_input[4324]), .B(p_input[34324]), .Z(n12613) );
  AND U18922 ( .A(n12615), .B(n12616), .Z(o[4323]) );
  AND U18923 ( .A(p_input[24323]), .B(p_input[14323]), .Z(n12616) );
  AND U18924 ( .A(p_input[4323]), .B(p_input[34323]), .Z(n12615) );
  AND U18925 ( .A(n12617), .B(n12618), .Z(o[4322]) );
  AND U18926 ( .A(p_input[24322]), .B(p_input[14322]), .Z(n12618) );
  AND U18927 ( .A(p_input[4322]), .B(p_input[34322]), .Z(n12617) );
  AND U18928 ( .A(n12619), .B(n12620), .Z(o[4321]) );
  AND U18929 ( .A(p_input[24321]), .B(p_input[14321]), .Z(n12620) );
  AND U18930 ( .A(p_input[4321]), .B(p_input[34321]), .Z(n12619) );
  AND U18931 ( .A(n12621), .B(n12622), .Z(o[4320]) );
  AND U18932 ( .A(p_input[24320]), .B(p_input[14320]), .Z(n12622) );
  AND U18933 ( .A(p_input[4320]), .B(p_input[34320]), .Z(n12621) );
  AND U18934 ( .A(n12623), .B(n12624), .Z(o[431]) );
  AND U18935 ( .A(p_input[20431]), .B(p_input[10431]), .Z(n12624) );
  AND U18936 ( .A(p_input[431]), .B(p_input[30431]), .Z(n12623) );
  AND U18937 ( .A(n12625), .B(n12626), .Z(o[4319]) );
  AND U18938 ( .A(p_input[24319]), .B(p_input[14319]), .Z(n12626) );
  AND U18939 ( .A(p_input[4319]), .B(p_input[34319]), .Z(n12625) );
  AND U18940 ( .A(n12627), .B(n12628), .Z(o[4318]) );
  AND U18941 ( .A(p_input[24318]), .B(p_input[14318]), .Z(n12628) );
  AND U18942 ( .A(p_input[4318]), .B(p_input[34318]), .Z(n12627) );
  AND U18943 ( .A(n12629), .B(n12630), .Z(o[4317]) );
  AND U18944 ( .A(p_input[24317]), .B(p_input[14317]), .Z(n12630) );
  AND U18945 ( .A(p_input[4317]), .B(p_input[34317]), .Z(n12629) );
  AND U18946 ( .A(n12631), .B(n12632), .Z(o[4316]) );
  AND U18947 ( .A(p_input[24316]), .B(p_input[14316]), .Z(n12632) );
  AND U18948 ( .A(p_input[4316]), .B(p_input[34316]), .Z(n12631) );
  AND U18949 ( .A(n12633), .B(n12634), .Z(o[4315]) );
  AND U18950 ( .A(p_input[24315]), .B(p_input[14315]), .Z(n12634) );
  AND U18951 ( .A(p_input[4315]), .B(p_input[34315]), .Z(n12633) );
  AND U18952 ( .A(n12635), .B(n12636), .Z(o[4314]) );
  AND U18953 ( .A(p_input[24314]), .B(p_input[14314]), .Z(n12636) );
  AND U18954 ( .A(p_input[4314]), .B(p_input[34314]), .Z(n12635) );
  AND U18955 ( .A(n12637), .B(n12638), .Z(o[4313]) );
  AND U18956 ( .A(p_input[24313]), .B(p_input[14313]), .Z(n12638) );
  AND U18957 ( .A(p_input[4313]), .B(p_input[34313]), .Z(n12637) );
  AND U18958 ( .A(n12639), .B(n12640), .Z(o[4312]) );
  AND U18959 ( .A(p_input[24312]), .B(p_input[14312]), .Z(n12640) );
  AND U18960 ( .A(p_input[4312]), .B(p_input[34312]), .Z(n12639) );
  AND U18961 ( .A(n12641), .B(n12642), .Z(o[4311]) );
  AND U18962 ( .A(p_input[24311]), .B(p_input[14311]), .Z(n12642) );
  AND U18963 ( .A(p_input[4311]), .B(p_input[34311]), .Z(n12641) );
  AND U18964 ( .A(n12643), .B(n12644), .Z(o[4310]) );
  AND U18965 ( .A(p_input[24310]), .B(p_input[14310]), .Z(n12644) );
  AND U18966 ( .A(p_input[4310]), .B(p_input[34310]), .Z(n12643) );
  AND U18967 ( .A(n12645), .B(n12646), .Z(o[430]) );
  AND U18968 ( .A(p_input[20430]), .B(p_input[10430]), .Z(n12646) );
  AND U18969 ( .A(p_input[430]), .B(p_input[30430]), .Z(n12645) );
  AND U18970 ( .A(n12647), .B(n12648), .Z(o[4309]) );
  AND U18971 ( .A(p_input[24309]), .B(p_input[14309]), .Z(n12648) );
  AND U18972 ( .A(p_input[4309]), .B(p_input[34309]), .Z(n12647) );
  AND U18973 ( .A(n12649), .B(n12650), .Z(o[4308]) );
  AND U18974 ( .A(p_input[24308]), .B(p_input[14308]), .Z(n12650) );
  AND U18975 ( .A(p_input[4308]), .B(p_input[34308]), .Z(n12649) );
  AND U18976 ( .A(n12651), .B(n12652), .Z(o[4307]) );
  AND U18977 ( .A(p_input[24307]), .B(p_input[14307]), .Z(n12652) );
  AND U18978 ( .A(p_input[4307]), .B(p_input[34307]), .Z(n12651) );
  AND U18979 ( .A(n12653), .B(n12654), .Z(o[4306]) );
  AND U18980 ( .A(p_input[24306]), .B(p_input[14306]), .Z(n12654) );
  AND U18981 ( .A(p_input[4306]), .B(p_input[34306]), .Z(n12653) );
  AND U18982 ( .A(n12655), .B(n12656), .Z(o[4305]) );
  AND U18983 ( .A(p_input[24305]), .B(p_input[14305]), .Z(n12656) );
  AND U18984 ( .A(p_input[4305]), .B(p_input[34305]), .Z(n12655) );
  AND U18985 ( .A(n12657), .B(n12658), .Z(o[4304]) );
  AND U18986 ( .A(p_input[24304]), .B(p_input[14304]), .Z(n12658) );
  AND U18987 ( .A(p_input[4304]), .B(p_input[34304]), .Z(n12657) );
  AND U18988 ( .A(n12659), .B(n12660), .Z(o[4303]) );
  AND U18989 ( .A(p_input[24303]), .B(p_input[14303]), .Z(n12660) );
  AND U18990 ( .A(p_input[4303]), .B(p_input[34303]), .Z(n12659) );
  AND U18991 ( .A(n12661), .B(n12662), .Z(o[4302]) );
  AND U18992 ( .A(p_input[24302]), .B(p_input[14302]), .Z(n12662) );
  AND U18993 ( .A(p_input[4302]), .B(p_input[34302]), .Z(n12661) );
  AND U18994 ( .A(n12663), .B(n12664), .Z(o[4301]) );
  AND U18995 ( .A(p_input[24301]), .B(p_input[14301]), .Z(n12664) );
  AND U18996 ( .A(p_input[4301]), .B(p_input[34301]), .Z(n12663) );
  AND U18997 ( .A(n12665), .B(n12666), .Z(o[4300]) );
  AND U18998 ( .A(p_input[24300]), .B(p_input[14300]), .Z(n12666) );
  AND U18999 ( .A(p_input[4300]), .B(p_input[34300]), .Z(n12665) );
  AND U19000 ( .A(n12667), .B(n12668), .Z(o[42]) );
  AND U19001 ( .A(p_input[20042]), .B(p_input[10042]), .Z(n12668) );
  AND U19002 ( .A(p_input[42]), .B(p_input[30042]), .Z(n12667) );
  AND U19003 ( .A(n12669), .B(n12670), .Z(o[429]) );
  AND U19004 ( .A(p_input[20429]), .B(p_input[10429]), .Z(n12670) );
  AND U19005 ( .A(p_input[429]), .B(p_input[30429]), .Z(n12669) );
  AND U19006 ( .A(n12671), .B(n12672), .Z(o[4299]) );
  AND U19007 ( .A(p_input[24299]), .B(p_input[14299]), .Z(n12672) );
  AND U19008 ( .A(p_input[4299]), .B(p_input[34299]), .Z(n12671) );
  AND U19009 ( .A(n12673), .B(n12674), .Z(o[4298]) );
  AND U19010 ( .A(p_input[24298]), .B(p_input[14298]), .Z(n12674) );
  AND U19011 ( .A(p_input[4298]), .B(p_input[34298]), .Z(n12673) );
  AND U19012 ( .A(n12675), .B(n12676), .Z(o[4297]) );
  AND U19013 ( .A(p_input[24297]), .B(p_input[14297]), .Z(n12676) );
  AND U19014 ( .A(p_input[4297]), .B(p_input[34297]), .Z(n12675) );
  AND U19015 ( .A(n12677), .B(n12678), .Z(o[4296]) );
  AND U19016 ( .A(p_input[24296]), .B(p_input[14296]), .Z(n12678) );
  AND U19017 ( .A(p_input[4296]), .B(p_input[34296]), .Z(n12677) );
  AND U19018 ( .A(n12679), .B(n12680), .Z(o[4295]) );
  AND U19019 ( .A(p_input[24295]), .B(p_input[14295]), .Z(n12680) );
  AND U19020 ( .A(p_input[4295]), .B(p_input[34295]), .Z(n12679) );
  AND U19021 ( .A(n12681), .B(n12682), .Z(o[4294]) );
  AND U19022 ( .A(p_input[24294]), .B(p_input[14294]), .Z(n12682) );
  AND U19023 ( .A(p_input[4294]), .B(p_input[34294]), .Z(n12681) );
  AND U19024 ( .A(n12683), .B(n12684), .Z(o[4293]) );
  AND U19025 ( .A(p_input[24293]), .B(p_input[14293]), .Z(n12684) );
  AND U19026 ( .A(p_input[4293]), .B(p_input[34293]), .Z(n12683) );
  AND U19027 ( .A(n12685), .B(n12686), .Z(o[4292]) );
  AND U19028 ( .A(p_input[24292]), .B(p_input[14292]), .Z(n12686) );
  AND U19029 ( .A(p_input[4292]), .B(p_input[34292]), .Z(n12685) );
  AND U19030 ( .A(n12687), .B(n12688), .Z(o[4291]) );
  AND U19031 ( .A(p_input[24291]), .B(p_input[14291]), .Z(n12688) );
  AND U19032 ( .A(p_input[4291]), .B(p_input[34291]), .Z(n12687) );
  AND U19033 ( .A(n12689), .B(n12690), .Z(o[4290]) );
  AND U19034 ( .A(p_input[24290]), .B(p_input[14290]), .Z(n12690) );
  AND U19035 ( .A(p_input[4290]), .B(p_input[34290]), .Z(n12689) );
  AND U19036 ( .A(n12691), .B(n12692), .Z(o[428]) );
  AND U19037 ( .A(p_input[20428]), .B(p_input[10428]), .Z(n12692) );
  AND U19038 ( .A(p_input[428]), .B(p_input[30428]), .Z(n12691) );
  AND U19039 ( .A(n12693), .B(n12694), .Z(o[4289]) );
  AND U19040 ( .A(p_input[24289]), .B(p_input[14289]), .Z(n12694) );
  AND U19041 ( .A(p_input[4289]), .B(p_input[34289]), .Z(n12693) );
  AND U19042 ( .A(n12695), .B(n12696), .Z(o[4288]) );
  AND U19043 ( .A(p_input[24288]), .B(p_input[14288]), .Z(n12696) );
  AND U19044 ( .A(p_input[4288]), .B(p_input[34288]), .Z(n12695) );
  AND U19045 ( .A(n12697), .B(n12698), .Z(o[4287]) );
  AND U19046 ( .A(p_input[24287]), .B(p_input[14287]), .Z(n12698) );
  AND U19047 ( .A(p_input[4287]), .B(p_input[34287]), .Z(n12697) );
  AND U19048 ( .A(n12699), .B(n12700), .Z(o[4286]) );
  AND U19049 ( .A(p_input[24286]), .B(p_input[14286]), .Z(n12700) );
  AND U19050 ( .A(p_input[4286]), .B(p_input[34286]), .Z(n12699) );
  AND U19051 ( .A(n12701), .B(n12702), .Z(o[4285]) );
  AND U19052 ( .A(p_input[24285]), .B(p_input[14285]), .Z(n12702) );
  AND U19053 ( .A(p_input[4285]), .B(p_input[34285]), .Z(n12701) );
  AND U19054 ( .A(n12703), .B(n12704), .Z(o[4284]) );
  AND U19055 ( .A(p_input[24284]), .B(p_input[14284]), .Z(n12704) );
  AND U19056 ( .A(p_input[4284]), .B(p_input[34284]), .Z(n12703) );
  AND U19057 ( .A(n12705), .B(n12706), .Z(o[4283]) );
  AND U19058 ( .A(p_input[24283]), .B(p_input[14283]), .Z(n12706) );
  AND U19059 ( .A(p_input[4283]), .B(p_input[34283]), .Z(n12705) );
  AND U19060 ( .A(n12707), .B(n12708), .Z(o[4282]) );
  AND U19061 ( .A(p_input[24282]), .B(p_input[14282]), .Z(n12708) );
  AND U19062 ( .A(p_input[4282]), .B(p_input[34282]), .Z(n12707) );
  AND U19063 ( .A(n12709), .B(n12710), .Z(o[4281]) );
  AND U19064 ( .A(p_input[24281]), .B(p_input[14281]), .Z(n12710) );
  AND U19065 ( .A(p_input[4281]), .B(p_input[34281]), .Z(n12709) );
  AND U19066 ( .A(n12711), .B(n12712), .Z(o[4280]) );
  AND U19067 ( .A(p_input[24280]), .B(p_input[14280]), .Z(n12712) );
  AND U19068 ( .A(p_input[4280]), .B(p_input[34280]), .Z(n12711) );
  AND U19069 ( .A(n12713), .B(n12714), .Z(o[427]) );
  AND U19070 ( .A(p_input[20427]), .B(p_input[10427]), .Z(n12714) );
  AND U19071 ( .A(p_input[427]), .B(p_input[30427]), .Z(n12713) );
  AND U19072 ( .A(n12715), .B(n12716), .Z(o[4279]) );
  AND U19073 ( .A(p_input[24279]), .B(p_input[14279]), .Z(n12716) );
  AND U19074 ( .A(p_input[4279]), .B(p_input[34279]), .Z(n12715) );
  AND U19075 ( .A(n12717), .B(n12718), .Z(o[4278]) );
  AND U19076 ( .A(p_input[24278]), .B(p_input[14278]), .Z(n12718) );
  AND U19077 ( .A(p_input[4278]), .B(p_input[34278]), .Z(n12717) );
  AND U19078 ( .A(n12719), .B(n12720), .Z(o[4277]) );
  AND U19079 ( .A(p_input[24277]), .B(p_input[14277]), .Z(n12720) );
  AND U19080 ( .A(p_input[4277]), .B(p_input[34277]), .Z(n12719) );
  AND U19081 ( .A(n12721), .B(n12722), .Z(o[4276]) );
  AND U19082 ( .A(p_input[24276]), .B(p_input[14276]), .Z(n12722) );
  AND U19083 ( .A(p_input[4276]), .B(p_input[34276]), .Z(n12721) );
  AND U19084 ( .A(n12723), .B(n12724), .Z(o[4275]) );
  AND U19085 ( .A(p_input[24275]), .B(p_input[14275]), .Z(n12724) );
  AND U19086 ( .A(p_input[4275]), .B(p_input[34275]), .Z(n12723) );
  AND U19087 ( .A(n12725), .B(n12726), .Z(o[4274]) );
  AND U19088 ( .A(p_input[24274]), .B(p_input[14274]), .Z(n12726) );
  AND U19089 ( .A(p_input[4274]), .B(p_input[34274]), .Z(n12725) );
  AND U19090 ( .A(n12727), .B(n12728), .Z(o[4273]) );
  AND U19091 ( .A(p_input[24273]), .B(p_input[14273]), .Z(n12728) );
  AND U19092 ( .A(p_input[4273]), .B(p_input[34273]), .Z(n12727) );
  AND U19093 ( .A(n12729), .B(n12730), .Z(o[4272]) );
  AND U19094 ( .A(p_input[24272]), .B(p_input[14272]), .Z(n12730) );
  AND U19095 ( .A(p_input[4272]), .B(p_input[34272]), .Z(n12729) );
  AND U19096 ( .A(n12731), .B(n12732), .Z(o[4271]) );
  AND U19097 ( .A(p_input[24271]), .B(p_input[14271]), .Z(n12732) );
  AND U19098 ( .A(p_input[4271]), .B(p_input[34271]), .Z(n12731) );
  AND U19099 ( .A(n12733), .B(n12734), .Z(o[4270]) );
  AND U19100 ( .A(p_input[24270]), .B(p_input[14270]), .Z(n12734) );
  AND U19101 ( .A(p_input[4270]), .B(p_input[34270]), .Z(n12733) );
  AND U19102 ( .A(n12735), .B(n12736), .Z(o[426]) );
  AND U19103 ( .A(p_input[20426]), .B(p_input[10426]), .Z(n12736) );
  AND U19104 ( .A(p_input[426]), .B(p_input[30426]), .Z(n12735) );
  AND U19105 ( .A(n12737), .B(n12738), .Z(o[4269]) );
  AND U19106 ( .A(p_input[24269]), .B(p_input[14269]), .Z(n12738) );
  AND U19107 ( .A(p_input[4269]), .B(p_input[34269]), .Z(n12737) );
  AND U19108 ( .A(n12739), .B(n12740), .Z(o[4268]) );
  AND U19109 ( .A(p_input[24268]), .B(p_input[14268]), .Z(n12740) );
  AND U19110 ( .A(p_input[4268]), .B(p_input[34268]), .Z(n12739) );
  AND U19111 ( .A(n12741), .B(n12742), .Z(o[4267]) );
  AND U19112 ( .A(p_input[24267]), .B(p_input[14267]), .Z(n12742) );
  AND U19113 ( .A(p_input[4267]), .B(p_input[34267]), .Z(n12741) );
  AND U19114 ( .A(n12743), .B(n12744), .Z(o[4266]) );
  AND U19115 ( .A(p_input[24266]), .B(p_input[14266]), .Z(n12744) );
  AND U19116 ( .A(p_input[4266]), .B(p_input[34266]), .Z(n12743) );
  AND U19117 ( .A(n12745), .B(n12746), .Z(o[4265]) );
  AND U19118 ( .A(p_input[24265]), .B(p_input[14265]), .Z(n12746) );
  AND U19119 ( .A(p_input[4265]), .B(p_input[34265]), .Z(n12745) );
  AND U19120 ( .A(n12747), .B(n12748), .Z(o[4264]) );
  AND U19121 ( .A(p_input[24264]), .B(p_input[14264]), .Z(n12748) );
  AND U19122 ( .A(p_input[4264]), .B(p_input[34264]), .Z(n12747) );
  AND U19123 ( .A(n12749), .B(n12750), .Z(o[4263]) );
  AND U19124 ( .A(p_input[24263]), .B(p_input[14263]), .Z(n12750) );
  AND U19125 ( .A(p_input[4263]), .B(p_input[34263]), .Z(n12749) );
  AND U19126 ( .A(n12751), .B(n12752), .Z(o[4262]) );
  AND U19127 ( .A(p_input[24262]), .B(p_input[14262]), .Z(n12752) );
  AND U19128 ( .A(p_input[4262]), .B(p_input[34262]), .Z(n12751) );
  AND U19129 ( .A(n12753), .B(n12754), .Z(o[4261]) );
  AND U19130 ( .A(p_input[24261]), .B(p_input[14261]), .Z(n12754) );
  AND U19131 ( .A(p_input[4261]), .B(p_input[34261]), .Z(n12753) );
  AND U19132 ( .A(n12755), .B(n12756), .Z(o[4260]) );
  AND U19133 ( .A(p_input[24260]), .B(p_input[14260]), .Z(n12756) );
  AND U19134 ( .A(p_input[4260]), .B(p_input[34260]), .Z(n12755) );
  AND U19135 ( .A(n12757), .B(n12758), .Z(o[425]) );
  AND U19136 ( .A(p_input[20425]), .B(p_input[10425]), .Z(n12758) );
  AND U19137 ( .A(p_input[425]), .B(p_input[30425]), .Z(n12757) );
  AND U19138 ( .A(n12759), .B(n12760), .Z(o[4259]) );
  AND U19139 ( .A(p_input[24259]), .B(p_input[14259]), .Z(n12760) );
  AND U19140 ( .A(p_input[4259]), .B(p_input[34259]), .Z(n12759) );
  AND U19141 ( .A(n12761), .B(n12762), .Z(o[4258]) );
  AND U19142 ( .A(p_input[24258]), .B(p_input[14258]), .Z(n12762) );
  AND U19143 ( .A(p_input[4258]), .B(p_input[34258]), .Z(n12761) );
  AND U19144 ( .A(n12763), .B(n12764), .Z(o[4257]) );
  AND U19145 ( .A(p_input[24257]), .B(p_input[14257]), .Z(n12764) );
  AND U19146 ( .A(p_input[4257]), .B(p_input[34257]), .Z(n12763) );
  AND U19147 ( .A(n12765), .B(n12766), .Z(o[4256]) );
  AND U19148 ( .A(p_input[24256]), .B(p_input[14256]), .Z(n12766) );
  AND U19149 ( .A(p_input[4256]), .B(p_input[34256]), .Z(n12765) );
  AND U19150 ( .A(n12767), .B(n12768), .Z(o[4255]) );
  AND U19151 ( .A(p_input[24255]), .B(p_input[14255]), .Z(n12768) );
  AND U19152 ( .A(p_input[4255]), .B(p_input[34255]), .Z(n12767) );
  AND U19153 ( .A(n12769), .B(n12770), .Z(o[4254]) );
  AND U19154 ( .A(p_input[24254]), .B(p_input[14254]), .Z(n12770) );
  AND U19155 ( .A(p_input[4254]), .B(p_input[34254]), .Z(n12769) );
  AND U19156 ( .A(n12771), .B(n12772), .Z(o[4253]) );
  AND U19157 ( .A(p_input[24253]), .B(p_input[14253]), .Z(n12772) );
  AND U19158 ( .A(p_input[4253]), .B(p_input[34253]), .Z(n12771) );
  AND U19159 ( .A(n12773), .B(n12774), .Z(o[4252]) );
  AND U19160 ( .A(p_input[24252]), .B(p_input[14252]), .Z(n12774) );
  AND U19161 ( .A(p_input[4252]), .B(p_input[34252]), .Z(n12773) );
  AND U19162 ( .A(n12775), .B(n12776), .Z(o[4251]) );
  AND U19163 ( .A(p_input[24251]), .B(p_input[14251]), .Z(n12776) );
  AND U19164 ( .A(p_input[4251]), .B(p_input[34251]), .Z(n12775) );
  AND U19165 ( .A(n12777), .B(n12778), .Z(o[4250]) );
  AND U19166 ( .A(p_input[24250]), .B(p_input[14250]), .Z(n12778) );
  AND U19167 ( .A(p_input[4250]), .B(p_input[34250]), .Z(n12777) );
  AND U19168 ( .A(n12779), .B(n12780), .Z(o[424]) );
  AND U19169 ( .A(p_input[20424]), .B(p_input[10424]), .Z(n12780) );
  AND U19170 ( .A(p_input[424]), .B(p_input[30424]), .Z(n12779) );
  AND U19171 ( .A(n12781), .B(n12782), .Z(o[4249]) );
  AND U19172 ( .A(p_input[24249]), .B(p_input[14249]), .Z(n12782) );
  AND U19173 ( .A(p_input[4249]), .B(p_input[34249]), .Z(n12781) );
  AND U19174 ( .A(n12783), .B(n12784), .Z(o[4248]) );
  AND U19175 ( .A(p_input[24248]), .B(p_input[14248]), .Z(n12784) );
  AND U19176 ( .A(p_input[4248]), .B(p_input[34248]), .Z(n12783) );
  AND U19177 ( .A(n12785), .B(n12786), .Z(o[4247]) );
  AND U19178 ( .A(p_input[24247]), .B(p_input[14247]), .Z(n12786) );
  AND U19179 ( .A(p_input[4247]), .B(p_input[34247]), .Z(n12785) );
  AND U19180 ( .A(n12787), .B(n12788), .Z(o[4246]) );
  AND U19181 ( .A(p_input[24246]), .B(p_input[14246]), .Z(n12788) );
  AND U19182 ( .A(p_input[4246]), .B(p_input[34246]), .Z(n12787) );
  AND U19183 ( .A(n12789), .B(n12790), .Z(o[4245]) );
  AND U19184 ( .A(p_input[24245]), .B(p_input[14245]), .Z(n12790) );
  AND U19185 ( .A(p_input[4245]), .B(p_input[34245]), .Z(n12789) );
  AND U19186 ( .A(n12791), .B(n12792), .Z(o[4244]) );
  AND U19187 ( .A(p_input[24244]), .B(p_input[14244]), .Z(n12792) );
  AND U19188 ( .A(p_input[4244]), .B(p_input[34244]), .Z(n12791) );
  AND U19189 ( .A(n12793), .B(n12794), .Z(o[4243]) );
  AND U19190 ( .A(p_input[24243]), .B(p_input[14243]), .Z(n12794) );
  AND U19191 ( .A(p_input[4243]), .B(p_input[34243]), .Z(n12793) );
  AND U19192 ( .A(n12795), .B(n12796), .Z(o[4242]) );
  AND U19193 ( .A(p_input[24242]), .B(p_input[14242]), .Z(n12796) );
  AND U19194 ( .A(p_input[4242]), .B(p_input[34242]), .Z(n12795) );
  AND U19195 ( .A(n12797), .B(n12798), .Z(o[4241]) );
  AND U19196 ( .A(p_input[24241]), .B(p_input[14241]), .Z(n12798) );
  AND U19197 ( .A(p_input[4241]), .B(p_input[34241]), .Z(n12797) );
  AND U19198 ( .A(n12799), .B(n12800), .Z(o[4240]) );
  AND U19199 ( .A(p_input[24240]), .B(p_input[14240]), .Z(n12800) );
  AND U19200 ( .A(p_input[4240]), .B(p_input[34240]), .Z(n12799) );
  AND U19201 ( .A(n12801), .B(n12802), .Z(o[423]) );
  AND U19202 ( .A(p_input[20423]), .B(p_input[10423]), .Z(n12802) );
  AND U19203 ( .A(p_input[423]), .B(p_input[30423]), .Z(n12801) );
  AND U19204 ( .A(n12803), .B(n12804), .Z(o[4239]) );
  AND U19205 ( .A(p_input[24239]), .B(p_input[14239]), .Z(n12804) );
  AND U19206 ( .A(p_input[4239]), .B(p_input[34239]), .Z(n12803) );
  AND U19207 ( .A(n12805), .B(n12806), .Z(o[4238]) );
  AND U19208 ( .A(p_input[24238]), .B(p_input[14238]), .Z(n12806) );
  AND U19209 ( .A(p_input[4238]), .B(p_input[34238]), .Z(n12805) );
  AND U19210 ( .A(n12807), .B(n12808), .Z(o[4237]) );
  AND U19211 ( .A(p_input[24237]), .B(p_input[14237]), .Z(n12808) );
  AND U19212 ( .A(p_input[4237]), .B(p_input[34237]), .Z(n12807) );
  AND U19213 ( .A(n12809), .B(n12810), .Z(o[4236]) );
  AND U19214 ( .A(p_input[24236]), .B(p_input[14236]), .Z(n12810) );
  AND U19215 ( .A(p_input[4236]), .B(p_input[34236]), .Z(n12809) );
  AND U19216 ( .A(n12811), .B(n12812), .Z(o[4235]) );
  AND U19217 ( .A(p_input[24235]), .B(p_input[14235]), .Z(n12812) );
  AND U19218 ( .A(p_input[4235]), .B(p_input[34235]), .Z(n12811) );
  AND U19219 ( .A(n12813), .B(n12814), .Z(o[4234]) );
  AND U19220 ( .A(p_input[24234]), .B(p_input[14234]), .Z(n12814) );
  AND U19221 ( .A(p_input[4234]), .B(p_input[34234]), .Z(n12813) );
  AND U19222 ( .A(n12815), .B(n12816), .Z(o[4233]) );
  AND U19223 ( .A(p_input[24233]), .B(p_input[14233]), .Z(n12816) );
  AND U19224 ( .A(p_input[4233]), .B(p_input[34233]), .Z(n12815) );
  AND U19225 ( .A(n12817), .B(n12818), .Z(o[4232]) );
  AND U19226 ( .A(p_input[24232]), .B(p_input[14232]), .Z(n12818) );
  AND U19227 ( .A(p_input[4232]), .B(p_input[34232]), .Z(n12817) );
  AND U19228 ( .A(n12819), .B(n12820), .Z(o[4231]) );
  AND U19229 ( .A(p_input[24231]), .B(p_input[14231]), .Z(n12820) );
  AND U19230 ( .A(p_input[4231]), .B(p_input[34231]), .Z(n12819) );
  AND U19231 ( .A(n12821), .B(n12822), .Z(o[4230]) );
  AND U19232 ( .A(p_input[24230]), .B(p_input[14230]), .Z(n12822) );
  AND U19233 ( .A(p_input[4230]), .B(p_input[34230]), .Z(n12821) );
  AND U19234 ( .A(n12823), .B(n12824), .Z(o[422]) );
  AND U19235 ( .A(p_input[20422]), .B(p_input[10422]), .Z(n12824) );
  AND U19236 ( .A(p_input[422]), .B(p_input[30422]), .Z(n12823) );
  AND U19237 ( .A(n12825), .B(n12826), .Z(o[4229]) );
  AND U19238 ( .A(p_input[24229]), .B(p_input[14229]), .Z(n12826) );
  AND U19239 ( .A(p_input[4229]), .B(p_input[34229]), .Z(n12825) );
  AND U19240 ( .A(n12827), .B(n12828), .Z(o[4228]) );
  AND U19241 ( .A(p_input[24228]), .B(p_input[14228]), .Z(n12828) );
  AND U19242 ( .A(p_input[4228]), .B(p_input[34228]), .Z(n12827) );
  AND U19243 ( .A(n12829), .B(n12830), .Z(o[4227]) );
  AND U19244 ( .A(p_input[24227]), .B(p_input[14227]), .Z(n12830) );
  AND U19245 ( .A(p_input[4227]), .B(p_input[34227]), .Z(n12829) );
  AND U19246 ( .A(n12831), .B(n12832), .Z(o[4226]) );
  AND U19247 ( .A(p_input[24226]), .B(p_input[14226]), .Z(n12832) );
  AND U19248 ( .A(p_input[4226]), .B(p_input[34226]), .Z(n12831) );
  AND U19249 ( .A(n12833), .B(n12834), .Z(o[4225]) );
  AND U19250 ( .A(p_input[24225]), .B(p_input[14225]), .Z(n12834) );
  AND U19251 ( .A(p_input[4225]), .B(p_input[34225]), .Z(n12833) );
  AND U19252 ( .A(n12835), .B(n12836), .Z(o[4224]) );
  AND U19253 ( .A(p_input[24224]), .B(p_input[14224]), .Z(n12836) );
  AND U19254 ( .A(p_input[4224]), .B(p_input[34224]), .Z(n12835) );
  AND U19255 ( .A(n12837), .B(n12838), .Z(o[4223]) );
  AND U19256 ( .A(p_input[24223]), .B(p_input[14223]), .Z(n12838) );
  AND U19257 ( .A(p_input[4223]), .B(p_input[34223]), .Z(n12837) );
  AND U19258 ( .A(n12839), .B(n12840), .Z(o[4222]) );
  AND U19259 ( .A(p_input[24222]), .B(p_input[14222]), .Z(n12840) );
  AND U19260 ( .A(p_input[4222]), .B(p_input[34222]), .Z(n12839) );
  AND U19261 ( .A(n12841), .B(n12842), .Z(o[4221]) );
  AND U19262 ( .A(p_input[24221]), .B(p_input[14221]), .Z(n12842) );
  AND U19263 ( .A(p_input[4221]), .B(p_input[34221]), .Z(n12841) );
  AND U19264 ( .A(n12843), .B(n12844), .Z(o[4220]) );
  AND U19265 ( .A(p_input[24220]), .B(p_input[14220]), .Z(n12844) );
  AND U19266 ( .A(p_input[4220]), .B(p_input[34220]), .Z(n12843) );
  AND U19267 ( .A(n12845), .B(n12846), .Z(o[421]) );
  AND U19268 ( .A(p_input[20421]), .B(p_input[10421]), .Z(n12846) );
  AND U19269 ( .A(p_input[421]), .B(p_input[30421]), .Z(n12845) );
  AND U19270 ( .A(n12847), .B(n12848), .Z(o[4219]) );
  AND U19271 ( .A(p_input[24219]), .B(p_input[14219]), .Z(n12848) );
  AND U19272 ( .A(p_input[4219]), .B(p_input[34219]), .Z(n12847) );
  AND U19273 ( .A(n12849), .B(n12850), .Z(o[4218]) );
  AND U19274 ( .A(p_input[24218]), .B(p_input[14218]), .Z(n12850) );
  AND U19275 ( .A(p_input[4218]), .B(p_input[34218]), .Z(n12849) );
  AND U19276 ( .A(n12851), .B(n12852), .Z(o[4217]) );
  AND U19277 ( .A(p_input[24217]), .B(p_input[14217]), .Z(n12852) );
  AND U19278 ( .A(p_input[4217]), .B(p_input[34217]), .Z(n12851) );
  AND U19279 ( .A(n12853), .B(n12854), .Z(o[4216]) );
  AND U19280 ( .A(p_input[24216]), .B(p_input[14216]), .Z(n12854) );
  AND U19281 ( .A(p_input[4216]), .B(p_input[34216]), .Z(n12853) );
  AND U19282 ( .A(n12855), .B(n12856), .Z(o[4215]) );
  AND U19283 ( .A(p_input[24215]), .B(p_input[14215]), .Z(n12856) );
  AND U19284 ( .A(p_input[4215]), .B(p_input[34215]), .Z(n12855) );
  AND U19285 ( .A(n12857), .B(n12858), .Z(o[4214]) );
  AND U19286 ( .A(p_input[24214]), .B(p_input[14214]), .Z(n12858) );
  AND U19287 ( .A(p_input[4214]), .B(p_input[34214]), .Z(n12857) );
  AND U19288 ( .A(n12859), .B(n12860), .Z(o[4213]) );
  AND U19289 ( .A(p_input[24213]), .B(p_input[14213]), .Z(n12860) );
  AND U19290 ( .A(p_input[4213]), .B(p_input[34213]), .Z(n12859) );
  AND U19291 ( .A(n12861), .B(n12862), .Z(o[4212]) );
  AND U19292 ( .A(p_input[24212]), .B(p_input[14212]), .Z(n12862) );
  AND U19293 ( .A(p_input[4212]), .B(p_input[34212]), .Z(n12861) );
  AND U19294 ( .A(n12863), .B(n12864), .Z(o[4211]) );
  AND U19295 ( .A(p_input[24211]), .B(p_input[14211]), .Z(n12864) );
  AND U19296 ( .A(p_input[4211]), .B(p_input[34211]), .Z(n12863) );
  AND U19297 ( .A(n12865), .B(n12866), .Z(o[4210]) );
  AND U19298 ( .A(p_input[24210]), .B(p_input[14210]), .Z(n12866) );
  AND U19299 ( .A(p_input[4210]), .B(p_input[34210]), .Z(n12865) );
  AND U19300 ( .A(n12867), .B(n12868), .Z(o[420]) );
  AND U19301 ( .A(p_input[20420]), .B(p_input[10420]), .Z(n12868) );
  AND U19302 ( .A(p_input[420]), .B(p_input[30420]), .Z(n12867) );
  AND U19303 ( .A(n12869), .B(n12870), .Z(o[4209]) );
  AND U19304 ( .A(p_input[24209]), .B(p_input[14209]), .Z(n12870) );
  AND U19305 ( .A(p_input[4209]), .B(p_input[34209]), .Z(n12869) );
  AND U19306 ( .A(n12871), .B(n12872), .Z(o[4208]) );
  AND U19307 ( .A(p_input[24208]), .B(p_input[14208]), .Z(n12872) );
  AND U19308 ( .A(p_input[4208]), .B(p_input[34208]), .Z(n12871) );
  AND U19309 ( .A(n12873), .B(n12874), .Z(o[4207]) );
  AND U19310 ( .A(p_input[24207]), .B(p_input[14207]), .Z(n12874) );
  AND U19311 ( .A(p_input[4207]), .B(p_input[34207]), .Z(n12873) );
  AND U19312 ( .A(n12875), .B(n12876), .Z(o[4206]) );
  AND U19313 ( .A(p_input[24206]), .B(p_input[14206]), .Z(n12876) );
  AND U19314 ( .A(p_input[4206]), .B(p_input[34206]), .Z(n12875) );
  AND U19315 ( .A(n12877), .B(n12878), .Z(o[4205]) );
  AND U19316 ( .A(p_input[24205]), .B(p_input[14205]), .Z(n12878) );
  AND U19317 ( .A(p_input[4205]), .B(p_input[34205]), .Z(n12877) );
  AND U19318 ( .A(n12879), .B(n12880), .Z(o[4204]) );
  AND U19319 ( .A(p_input[24204]), .B(p_input[14204]), .Z(n12880) );
  AND U19320 ( .A(p_input[4204]), .B(p_input[34204]), .Z(n12879) );
  AND U19321 ( .A(n12881), .B(n12882), .Z(o[4203]) );
  AND U19322 ( .A(p_input[24203]), .B(p_input[14203]), .Z(n12882) );
  AND U19323 ( .A(p_input[4203]), .B(p_input[34203]), .Z(n12881) );
  AND U19324 ( .A(n12883), .B(n12884), .Z(o[4202]) );
  AND U19325 ( .A(p_input[24202]), .B(p_input[14202]), .Z(n12884) );
  AND U19326 ( .A(p_input[4202]), .B(p_input[34202]), .Z(n12883) );
  AND U19327 ( .A(n12885), .B(n12886), .Z(o[4201]) );
  AND U19328 ( .A(p_input[24201]), .B(p_input[14201]), .Z(n12886) );
  AND U19329 ( .A(p_input[4201]), .B(p_input[34201]), .Z(n12885) );
  AND U19330 ( .A(n12887), .B(n12888), .Z(o[4200]) );
  AND U19331 ( .A(p_input[24200]), .B(p_input[14200]), .Z(n12888) );
  AND U19332 ( .A(p_input[4200]), .B(p_input[34200]), .Z(n12887) );
  AND U19333 ( .A(n12889), .B(n12890), .Z(o[41]) );
  AND U19334 ( .A(p_input[20041]), .B(p_input[10041]), .Z(n12890) );
  AND U19335 ( .A(p_input[41]), .B(p_input[30041]), .Z(n12889) );
  AND U19336 ( .A(n12891), .B(n12892), .Z(o[419]) );
  AND U19337 ( .A(p_input[20419]), .B(p_input[10419]), .Z(n12892) );
  AND U19338 ( .A(p_input[419]), .B(p_input[30419]), .Z(n12891) );
  AND U19339 ( .A(n12893), .B(n12894), .Z(o[4199]) );
  AND U19340 ( .A(p_input[24199]), .B(p_input[14199]), .Z(n12894) );
  AND U19341 ( .A(p_input[4199]), .B(p_input[34199]), .Z(n12893) );
  AND U19342 ( .A(n12895), .B(n12896), .Z(o[4198]) );
  AND U19343 ( .A(p_input[24198]), .B(p_input[14198]), .Z(n12896) );
  AND U19344 ( .A(p_input[4198]), .B(p_input[34198]), .Z(n12895) );
  AND U19345 ( .A(n12897), .B(n12898), .Z(o[4197]) );
  AND U19346 ( .A(p_input[24197]), .B(p_input[14197]), .Z(n12898) );
  AND U19347 ( .A(p_input[4197]), .B(p_input[34197]), .Z(n12897) );
  AND U19348 ( .A(n12899), .B(n12900), .Z(o[4196]) );
  AND U19349 ( .A(p_input[24196]), .B(p_input[14196]), .Z(n12900) );
  AND U19350 ( .A(p_input[4196]), .B(p_input[34196]), .Z(n12899) );
  AND U19351 ( .A(n12901), .B(n12902), .Z(o[4195]) );
  AND U19352 ( .A(p_input[24195]), .B(p_input[14195]), .Z(n12902) );
  AND U19353 ( .A(p_input[4195]), .B(p_input[34195]), .Z(n12901) );
  AND U19354 ( .A(n12903), .B(n12904), .Z(o[4194]) );
  AND U19355 ( .A(p_input[24194]), .B(p_input[14194]), .Z(n12904) );
  AND U19356 ( .A(p_input[4194]), .B(p_input[34194]), .Z(n12903) );
  AND U19357 ( .A(n12905), .B(n12906), .Z(o[4193]) );
  AND U19358 ( .A(p_input[24193]), .B(p_input[14193]), .Z(n12906) );
  AND U19359 ( .A(p_input[4193]), .B(p_input[34193]), .Z(n12905) );
  AND U19360 ( .A(n12907), .B(n12908), .Z(o[4192]) );
  AND U19361 ( .A(p_input[24192]), .B(p_input[14192]), .Z(n12908) );
  AND U19362 ( .A(p_input[4192]), .B(p_input[34192]), .Z(n12907) );
  AND U19363 ( .A(n12909), .B(n12910), .Z(o[4191]) );
  AND U19364 ( .A(p_input[24191]), .B(p_input[14191]), .Z(n12910) );
  AND U19365 ( .A(p_input[4191]), .B(p_input[34191]), .Z(n12909) );
  AND U19366 ( .A(n12911), .B(n12912), .Z(o[4190]) );
  AND U19367 ( .A(p_input[24190]), .B(p_input[14190]), .Z(n12912) );
  AND U19368 ( .A(p_input[4190]), .B(p_input[34190]), .Z(n12911) );
  AND U19369 ( .A(n12913), .B(n12914), .Z(o[418]) );
  AND U19370 ( .A(p_input[20418]), .B(p_input[10418]), .Z(n12914) );
  AND U19371 ( .A(p_input[418]), .B(p_input[30418]), .Z(n12913) );
  AND U19372 ( .A(n12915), .B(n12916), .Z(o[4189]) );
  AND U19373 ( .A(p_input[24189]), .B(p_input[14189]), .Z(n12916) );
  AND U19374 ( .A(p_input[4189]), .B(p_input[34189]), .Z(n12915) );
  AND U19375 ( .A(n12917), .B(n12918), .Z(o[4188]) );
  AND U19376 ( .A(p_input[24188]), .B(p_input[14188]), .Z(n12918) );
  AND U19377 ( .A(p_input[4188]), .B(p_input[34188]), .Z(n12917) );
  AND U19378 ( .A(n12919), .B(n12920), .Z(o[4187]) );
  AND U19379 ( .A(p_input[24187]), .B(p_input[14187]), .Z(n12920) );
  AND U19380 ( .A(p_input[4187]), .B(p_input[34187]), .Z(n12919) );
  AND U19381 ( .A(n12921), .B(n12922), .Z(o[4186]) );
  AND U19382 ( .A(p_input[24186]), .B(p_input[14186]), .Z(n12922) );
  AND U19383 ( .A(p_input[4186]), .B(p_input[34186]), .Z(n12921) );
  AND U19384 ( .A(n12923), .B(n12924), .Z(o[4185]) );
  AND U19385 ( .A(p_input[24185]), .B(p_input[14185]), .Z(n12924) );
  AND U19386 ( .A(p_input[4185]), .B(p_input[34185]), .Z(n12923) );
  AND U19387 ( .A(n12925), .B(n12926), .Z(o[4184]) );
  AND U19388 ( .A(p_input[24184]), .B(p_input[14184]), .Z(n12926) );
  AND U19389 ( .A(p_input[4184]), .B(p_input[34184]), .Z(n12925) );
  AND U19390 ( .A(n12927), .B(n12928), .Z(o[4183]) );
  AND U19391 ( .A(p_input[24183]), .B(p_input[14183]), .Z(n12928) );
  AND U19392 ( .A(p_input[4183]), .B(p_input[34183]), .Z(n12927) );
  AND U19393 ( .A(n12929), .B(n12930), .Z(o[4182]) );
  AND U19394 ( .A(p_input[24182]), .B(p_input[14182]), .Z(n12930) );
  AND U19395 ( .A(p_input[4182]), .B(p_input[34182]), .Z(n12929) );
  AND U19396 ( .A(n12931), .B(n12932), .Z(o[4181]) );
  AND U19397 ( .A(p_input[24181]), .B(p_input[14181]), .Z(n12932) );
  AND U19398 ( .A(p_input[4181]), .B(p_input[34181]), .Z(n12931) );
  AND U19399 ( .A(n12933), .B(n12934), .Z(o[4180]) );
  AND U19400 ( .A(p_input[24180]), .B(p_input[14180]), .Z(n12934) );
  AND U19401 ( .A(p_input[4180]), .B(p_input[34180]), .Z(n12933) );
  AND U19402 ( .A(n12935), .B(n12936), .Z(o[417]) );
  AND U19403 ( .A(p_input[20417]), .B(p_input[10417]), .Z(n12936) );
  AND U19404 ( .A(p_input[417]), .B(p_input[30417]), .Z(n12935) );
  AND U19405 ( .A(n12937), .B(n12938), .Z(o[4179]) );
  AND U19406 ( .A(p_input[24179]), .B(p_input[14179]), .Z(n12938) );
  AND U19407 ( .A(p_input[4179]), .B(p_input[34179]), .Z(n12937) );
  AND U19408 ( .A(n12939), .B(n12940), .Z(o[4178]) );
  AND U19409 ( .A(p_input[24178]), .B(p_input[14178]), .Z(n12940) );
  AND U19410 ( .A(p_input[4178]), .B(p_input[34178]), .Z(n12939) );
  AND U19411 ( .A(n12941), .B(n12942), .Z(o[4177]) );
  AND U19412 ( .A(p_input[24177]), .B(p_input[14177]), .Z(n12942) );
  AND U19413 ( .A(p_input[4177]), .B(p_input[34177]), .Z(n12941) );
  AND U19414 ( .A(n12943), .B(n12944), .Z(o[4176]) );
  AND U19415 ( .A(p_input[24176]), .B(p_input[14176]), .Z(n12944) );
  AND U19416 ( .A(p_input[4176]), .B(p_input[34176]), .Z(n12943) );
  AND U19417 ( .A(n12945), .B(n12946), .Z(o[4175]) );
  AND U19418 ( .A(p_input[24175]), .B(p_input[14175]), .Z(n12946) );
  AND U19419 ( .A(p_input[4175]), .B(p_input[34175]), .Z(n12945) );
  AND U19420 ( .A(n12947), .B(n12948), .Z(o[4174]) );
  AND U19421 ( .A(p_input[24174]), .B(p_input[14174]), .Z(n12948) );
  AND U19422 ( .A(p_input[4174]), .B(p_input[34174]), .Z(n12947) );
  AND U19423 ( .A(n12949), .B(n12950), .Z(o[4173]) );
  AND U19424 ( .A(p_input[24173]), .B(p_input[14173]), .Z(n12950) );
  AND U19425 ( .A(p_input[4173]), .B(p_input[34173]), .Z(n12949) );
  AND U19426 ( .A(n12951), .B(n12952), .Z(o[4172]) );
  AND U19427 ( .A(p_input[24172]), .B(p_input[14172]), .Z(n12952) );
  AND U19428 ( .A(p_input[4172]), .B(p_input[34172]), .Z(n12951) );
  AND U19429 ( .A(n12953), .B(n12954), .Z(o[4171]) );
  AND U19430 ( .A(p_input[24171]), .B(p_input[14171]), .Z(n12954) );
  AND U19431 ( .A(p_input[4171]), .B(p_input[34171]), .Z(n12953) );
  AND U19432 ( .A(n12955), .B(n12956), .Z(o[4170]) );
  AND U19433 ( .A(p_input[24170]), .B(p_input[14170]), .Z(n12956) );
  AND U19434 ( .A(p_input[4170]), .B(p_input[34170]), .Z(n12955) );
  AND U19435 ( .A(n12957), .B(n12958), .Z(o[416]) );
  AND U19436 ( .A(p_input[20416]), .B(p_input[10416]), .Z(n12958) );
  AND U19437 ( .A(p_input[416]), .B(p_input[30416]), .Z(n12957) );
  AND U19438 ( .A(n12959), .B(n12960), .Z(o[4169]) );
  AND U19439 ( .A(p_input[24169]), .B(p_input[14169]), .Z(n12960) );
  AND U19440 ( .A(p_input[4169]), .B(p_input[34169]), .Z(n12959) );
  AND U19441 ( .A(n12961), .B(n12962), .Z(o[4168]) );
  AND U19442 ( .A(p_input[24168]), .B(p_input[14168]), .Z(n12962) );
  AND U19443 ( .A(p_input[4168]), .B(p_input[34168]), .Z(n12961) );
  AND U19444 ( .A(n12963), .B(n12964), .Z(o[4167]) );
  AND U19445 ( .A(p_input[24167]), .B(p_input[14167]), .Z(n12964) );
  AND U19446 ( .A(p_input[4167]), .B(p_input[34167]), .Z(n12963) );
  AND U19447 ( .A(n12965), .B(n12966), .Z(o[4166]) );
  AND U19448 ( .A(p_input[24166]), .B(p_input[14166]), .Z(n12966) );
  AND U19449 ( .A(p_input[4166]), .B(p_input[34166]), .Z(n12965) );
  AND U19450 ( .A(n12967), .B(n12968), .Z(o[4165]) );
  AND U19451 ( .A(p_input[24165]), .B(p_input[14165]), .Z(n12968) );
  AND U19452 ( .A(p_input[4165]), .B(p_input[34165]), .Z(n12967) );
  AND U19453 ( .A(n12969), .B(n12970), .Z(o[4164]) );
  AND U19454 ( .A(p_input[24164]), .B(p_input[14164]), .Z(n12970) );
  AND U19455 ( .A(p_input[4164]), .B(p_input[34164]), .Z(n12969) );
  AND U19456 ( .A(n12971), .B(n12972), .Z(o[4163]) );
  AND U19457 ( .A(p_input[24163]), .B(p_input[14163]), .Z(n12972) );
  AND U19458 ( .A(p_input[4163]), .B(p_input[34163]), .Z(n12971) );
  AND U19459 ( .A(n12973), .B(n12974), .Z(o[4162]) );
  AND U19460 ( .A(p_input[24162]), .B(p_input[14162]), .Z(n12974) );
  AND U19461 ( .A(p_input[4162]), .B(p_input[34162]), .Z(n12973) );
  AND U19462 ( .A(n12975), .B(n12976), .Z(o[4161]) );
  AND U19463 ( .A(p_input[24161]), .B(p_input[14161]), .Z(n12976) );
  AND U19464 ( .A(p_input[4161]), .B(p_input[34161]), .Z(n12975) );
  AND U19465 ( .A(n12977), .B(n12978), .Z(o[4160]) );
  AND U19466 ( .A(p_input[24160]), .B(p_input[14160]), .Z(n12978) );
  AND U19467 ( .A(p_input[4160]), .B(p_input[34160]), .Z(n12977) );
  AND U19468 ( .A(n12979), .B(n12980), .Z(o[415]) );
  AND U19469 ( .A(p_input[20415]), .B(p_input[10415]), .Z(n12980) );
  AND U19470 ( .A(p_input[415]), .B(p_input[30415]), .Z(n12979) );
  AND U19471 ( .A(n12981), .B(n12982), .Z(o[4159]) );
  AND U19472 ( .A(p_input[24159]), .B(p_input[14159]), .Z(n12982) );
  AND U19473 ( .A(p_input[4159]), .B(p_input[34159]), .Z(n12981) );
  AND U19474 ( .A(n12983), .B(n12984), .Z(o[4158]) );
  AND U19475 ( .A(p_input[24158]), .B(p_input[14158]), .Z(n12984) );
  AND U19476 ( .A(p_input[4158]), .B(p_input[34158]), .Z(n12983) );
  AND U19477 ( .A(n12985), .B(n12986), .Z(o[4157]) );
  AND U19478 ( .A(p_input[24157]), .B(p_input[14157]), .Z(n12986) );
  AND U19479 ( .A(p_input[4157]), .B(p_input[34157]), .Z(n12985) );
  AND U19480 ( .A(n12987), .B(n12988), .Z(o[4156]) );
  AND U19481 ( .A(p_input[24156]), .B(p_input[14156]), .Z(n12988) );
  AND U19482 ( .A(p_input[4156]), .B(p_input[34156]), .Z(n12987) );
  AND U19483 ( .A(n12989), .B(n12990), .Z(o[4155]) );
  AND U19484 ( .A(p_input[24155]), .B(p_input[14155]), .Z(n12990) );
  AND U19485 ( .A(p_input[4155]), .B(p_input[34155]), .Z(n12989) );
  AND U19486 ( .A(n12991), .B(n12992), .Z(o[4154]) );
  AND U19487 ( .A(p_input[24154]), .B(p_input[14154]), .Z(n12992) );
  AND U19488 ( .A(p_input[4154]), .B(p_input[34154]), .Z(n12991) );
  AND U19489 ( .A(n12993), .B(n12994), .Z(o[4153]) );
  AND U19490 ( .A(p_input[24153]), .B(p_input[14153]), .Z(n12994) );
  AND U19491 ( .A(p_input[4153]), .B(p_input[34153]), .Z(n12993) );
  AND U19492 ( .A(n12995), .B(n12996), .Z(o[4152]) );
  AND U19493 ( .A(p_input[24152]), .B(p_input[14152]), .Z(n12996) );
  AND U19494 ( .A(p_input[4152]), .B(p_input[34152]), .Z(n12995) );
  AND U19495 ( .A(n12997), .B(n12998), .Z(o[4151]) );
  AND U19496 ( .A(p_input[24151]), .B(p_input[14151]), .Z(n12998) );
  AND U19497 ( .A(p_input[4151]), .B(p_input[34151]), .Z(n12997) );
  AND U19498 ( .A(n12999), .B(n13000), .Z(o[4150]) );
  AND U19499 ( .A(p_input[24150]), .B(p_input[14150]), .Z(n13000) );
  AND U19500 ( .A(p_input[4150]), .B(p_input[34150]), .Z(n12999) );
  AND U19501 ( .A(n13001), .B(n13002), .Z(o[414]) );
  AND U19502 ( .A(p_input[20414]), .B(p_input[10414]), .Z(n13002) );
  AND U19503 ( .A(p_input[414]), .B(p_input[30414]), .Z(n13001) );
  AND U19504 ( .A(n13003), .B(n13004), .Z(o[4149]) );
  AND U19505 ( .A(p_input[24149]), .B(p_input[14149]), .Z(n13004) );
  AND U19506 ( .A(p_input[4149]), .B(p_input[34149]), .Z(n13003) );
  AND U19507 ( .A(n13005), .B(n13006), .Z(o[4148]) );
  AND U19508 ( .A(p_input[24148]), .B(p_input[14148]), .Z(n13006) );
  AND U19509 ( .A(p_input[4148]), .B(p_input[34148]), .Z(n13005) );
  AND U19510 ( .A(n13007), .B(n13008), .Z(o[4147]) );
  AND U19511 ( .A(p_input[24147]), .B(p_input[14147]), .Z(n13008) );
  AND U19512 ( .A(p_input[4147]), .B(p_input[34147]), .Z(n13007) );
  AND U19513 ( .A(n13009), .B(n13010), .Z(o[4146]) );
  AND U19514 ( .A(p_input[24146]), .B(p_input[14146]), .Z(n13010) );
  AND U19515 ( .A(p_input[4146]), .B(p_input[34146]), .Z(n13009) );
  AND U19516 ( .A(n13011), .B(n13012), .Z(o[4145]) );
  AND U19517 ( .A(p_input[24145]), .B(p_input[14145]), .Z(n13012) );
  AND U19518 ( .A(p_input[4145]), .B(p_input[34145]), .Z(n13011) );
  AND U19519 ( .A(n13013), .B(n13014), .Z(o[4144]) );
  AND U19520 ( .A(p_input[24144]), .B(p_input[14144]), .Z(n13014) );
  AND U19521 ( .A(p_input[4144]), .B(p_input[34144]), .Z(n13013) );
  AND U19522 ( .A(n13015), .B(n13016), .Z(o[4143]) );
  AND U19523 ( .A(p_input[24143]), .B(p_input[14143]), .Z(n13016) );
  AND U19524 ( .A(p_input[4143]), .B(p_input[34143]), .Z(n13015) );
  AND U19525 ( .A(n13017), .B(n13018), .Z(o[4142]) );
  AND U19526 ( .A(p_input[24142]), .B(p_input[14142]), .Z(n13018) );
  AND U19527 ( .A(p_input[4142]), .B(p_input[34142]), .Z(n13017) );
  AND U19528 ( .A(n13019), .B(n13020), .Z(o[4141]) );
  AND U19529 ( .A(p_input[24141]), .B(p_input[14141]), .Z(n13020) );
  AND U19530 ( .A(p_input[4141]), .B(p_input[34141]), .Z(n13019) );
  AND U19531 ( .A(n13021), .B(n13022), .Z(o[4140]) );
  AND U19532 ( .A(p_input[24140]), .B(p_input[14140]), .Z(n13022) );
  AND U19533 ( .A(p_input[4140]), .B(p_input[34140]), .Z(n13021) );
  AND U19534 ( .A(n13023), .B(n13024), .Z(o[413]) );
  AND U19535 ( .A(p_input[20413]), .B(p_input[10413]), .Z(n13024) );
  AND U19536 ( .A(p_input[413]), .B(p_input[30413]), .Z(n13023) );
  AND U19537 ( .A(n13025), .B(n13026), .Z(o[4139]) );
  AND U19538 ( .A(p_input[24139]), .B(p_input[14139]), .Z(n13026) );
  AND U19539 ( .A(p_input[4139]), .B(p_input[34139]), .Z(n13025) );
  AND U19540 ( .A(n13027), .B(n13028), .Z(o[4138]) );
  AND U19541 ( .A(p_input[24138]), .B(p_input[14138]), .Z(n13028) );
  AND U19542 ( .A(p_input[4138]), .B(p_input[34138]), .Z(n13027) );
  AND U19543 ( .A(n13029), .B(n13030), .Z(o[4137]) );
  AND U19544 ( .A(p_input[24137]), .B(p_input[14137]), .Z(n13030) );
  AND U19545 ( .A(p_input[4137]), .B(p_input[34137]), .Z(n13029) );
  AND U19546 ( .A(n13031), .B(n13032), .Z(o[4136]) );
  AND U19547 ( .A(p_input[24136]), .B(p_input[14136]), .Z(n13032) );
  AND U19548 ( .A(p_input[4136]), .B(p_input[34136]), .Z(n13031) );
  AND U19549 ( .A(n13033), .B(n13034), .Z(o[4135]) );
  AND U19550 ( .A(p_input[24135]), .B(p_input[14135]), .Z(n13034) );
  AND U19551 ( .A(p_input[4135]), .B(p_input[34135]), .Z(n13033) );
  AND U19552 ( .A(n13035), .B(n13036), .Z(o[4134]) );
  AND U19553 ( .A(p_input[24134]), .B(p_input[14134]), .Z(n13036) );
  AND U19554 ( .A(p_input[4134]), .B(p_input[34134]), .Z(n13035) );
  AND U19555 ( .A(n13037), .B(n13038), .Z(o[4133]) );
  AND U19556 ( .A(p_input[24133]), .B(p_input[14133]), .Z(n13038) );
  AND U19557 ( .A(p_input[4133]), .B(p_input[34133]), .Z(n13037) );
  AND U19558 ( .A(n13039), .B(n13040), .Z(o[4132]) );
  AND U19559 ( .A(p_input[24132]), .B(p_input[14132]), .Z(n13040) );
  AND U19560 ( .A(p_input[4132]), .B(p_input[34132]), .Z(n13039) );
  AND U19561 ( .A(n13041), .B(n13042), .Z(o[4131]) );
  AND U19562 ( .A(p_input[24131]), .B(p_input[14131]), .Z(n13042) );
  AND U19563 ( .A(p_input[4131]), .B(p_input[34131]), .Z(n13041) );
  AND U19564 ( .A(n13043), .B(n13044), .Z(o[4130]) );
  AND U19565 ( .A(p_input[24130]), .B(p_input[14130]), .Z(n13044) );
  AND U19566 ( .A(p_input[4130]), .B(p_input[34130]), .Z(n13043) );
  AND U19567 ( .A(n13045), .B(n13046), .Z(o[412]) );
  AND U19568 ( .A(p_input[20412]), .B(p_input[10412]), .Z(n13046) );
  AND U19569 ( .A(p_input[412]), .B(p_input[30412]), .Z(n13045) );
  AND U19570 ( .A(n13047), .B(n13048), .Z(o[4129]) );
  AND U19571 ( .A(p_input[24129]), .B(p_input[14129]), .Z(n13048) );
  AND U19572 ( .A(p_input[4129]), .B(p_input[34129]), .Z(n13047) );
  AND U19573 ( .A(n13049), .B(n13050), .Z(o[4128]) );
  AND U19574 ( .A(p_input[24128]), .B(p_input[14128]), .Z(n13050) );
  AND U19575 ( .A(p_input[4128]), .B(p_input[34128]), .Z(n13049) );
  AND U19576 ( .A(n13051), .B(n13052), .Z(o[4127]) );
  AND U19577 ( .A(p_input[24127]), .B(p_input[14127]), .Z(n13052) );
  AND U19578 ( .A(p_input[4127]), .B(p_input[34127]), .Z(n13051) );
  AND U19579 ( .A(n13053), .B(n13054), .Z(o[4126]) );
  AND U19580 ( .A(p_input[24126]), .B(p_input[14126]), .Z(n13054) );
  AND U19581 ( .A(p_input[4126]), .B(p_input[34126]), .Z(n13053) );
  AND U19582 ( .A(n13055), .B(n13056), .Z(o[4125]) );
  AND U19583 ( .A(p_input[24125]), .B(p_input[14125]), .Z(n13056) );
  AND U19584 ( .A(p_input[4125]), .B(p_input[34125]), .Z(n13055) );
  AND U19585 ( .A(n13057), .B(n13058), .Z(o[4124]) );
  AND U19586 ( .A(p_input[24124]), .B(p_input[14124]), .Z(n13058) );
  AND U19587 ( .A(p_input[4124]), .B(p_input[34124]), .Z(n13057) );
  AND U19588 ( .A(n13059), .B(n13060), .Z(o[4123]) );
  AND U19589 ( .A(p_input[24123]), .B(p_input[14123]), .Z(n13060) );
  AND U19590 ( .A(p_input[4123]), .B(p_input[34123]), .Z(n13059) );
  AND U19591 ( .A(n13061), .B(n13062), .Z(o[4122]) );
  AND U19592 ( .A(p_input[24122]), .B(p_input[14122]), .Z(n13062) );
  AND U19593 ( .A(p_input[4122]), .B(p_input[34122]), .Z(n13061) );
  AND U19594 ( .A(n13063), .B(n13064), .Z(o[4121]) );
  AND U19595 ( .A(p_input[24121]), .B(p_input[14121]), .Z(n13064) );
  AND U19596 ( .A(p_input[4121]), .B(p_input[34121]), .Z(n13063) );
  AND U19597 ( .A(n13065), .B(n13066), .Z(o[4120]) );
  AND U19598 ( .A(p_input[24120]), .B(p_input[14120]), .Z(n13066) );
  AND U19599 ( .A(p_input[4120]), .B(p_input[34120]), .Z(n13065) );
  AND U19600 ( .A(n13067), .B(n13068), .Z(o[411]) );
  AND U19601 ( .A(p_input[20411]), .B(p_input[10411]), .Z(n13068) );
  AND U19602 ( .A(p_input[411]), .B(p_input[30411]), .Z(n13067) );
  AND U19603 ( .A(n13069), .B(n13070), .Z(o[4119]) );
  AND U19604 ( .A(p_input[24119]), .B(p_input[14119]), .Z(n13070) );
  AND U19605 ( .A(p_input[4119]), .B(p_input[34119]), .Z(n13069) );
  AND U19606 ( .A(n13071), .B(n13072), .Z(o[4118]) );
  AND U19607 ( .A(p_input[24118]), .B(p_input[14118]), .Z(n13072) );
  AND U19608 ( .A(p_input[4118]), .B(p_input[34118]), .Z(n13071) );
  AND U19609 ( .A(n13073), .B(n13074), .Z(o[4117]) );
  AND U19610 ( .A(p_input[24117]), .B(p_input[14117]), .Z(n13074) );
  AND U19611 ( .A(p_input[4117]), .B(p_input[34117]), .Z(n13073) );
  AND U19612 ( .A(n13075), .B(n13076), .Z(o[4116]) );
  AND U19613 ( .A(p_input[24116]), .B(p_input[14116]), .Z(n13076) );
  AND U19614 ( .A(p_input[4116]), .B(p_input[34116]), .Z(n13075) );
  AND U19615 ( .A(n13077), .B(n13078), .Z(o[4115]) );
  AND U19616 ( .A(p_input[24115]), .B(p_input[14115]), .Z(n13078) );
  AND U19617 ( .A(p_input[4115]), .B(p_input[34115]), .Z(n13077) );
  AND U19618 ( .A(n13079), .B(n13080), .Z(o[4114]) );
  AND U19619 ( .A(p_input[24114]), .B(p_input[14114]), .Z(n13080) );
  AND U19620 ( .A(p_input[4114]), .B(p_input[34114]), .Z(n13079) );
  AND U19621 ( .A(n13081), .B(n13082), .Z(o[4113]) );
  AND U19622 ( .A(p_input[24113]), .B(p_input[14113]), .Z(n13082) );
  AND U19623 ( .A(p_input[4113]), .B(p_input[34113]), .Z(n13081) );
  AND U19624 ( .A(n13083), .B(n13084), .Z(o[4112]) );
  AND U19625 ( .A(p_input[24112]), .B(p_input[14112]), .Z(n13084) );
  AND U19626 ( .A(p_input[4112]), .B(p_input[34112]), .Z(n13083) );
  AND U19627 ( .A(n13085), .B(n13086), .Z(o[4111]) );
  AND U19628 ( .A(p_input[24111]), .B(p_input[14111]), .Z(n13086) );
  AND U19629 ( .A(p_input[4111]), .B(p_input[34111]), .Z(n13085) );
  AND U19630 ( .A(n13087), .B(n13088), .Z(o[4110]) );
  AND U19631 ( .A(p_input[24110]), .B(p_input[14110]), .Z(n13088) );
  AND U19632 ( .A(p_input[4110]), .B(p_input[34110]), .Z(n13087) );
  AND U19633 ( .A(n13089), .B(n13090), .Z(o[410]) );
  AND U19634 ( .A(p_input[20410]), .B(p_input[10410]), .Z(n13090) );
  AND U19635 ( .A(p_input[410]), .B(p_input[30410]), .Z(n13089) );
  AND U19636 ( .A(n13091), .B(n13092), .Z(o[4109]) );
  AND U19637 ( .A(p_input[24109]), .B(p_input[14109]), .Z(n13092) );
  AND U19638 ( .A(p_input[4109]), .B(p_input[34109]), .Z(n13091) );
  AND U19639 ( .A(n13093), .B(n13094), .Z(o[4108]) );
  AND U19640 ( .A(p_input[24108]), .B(p_input[14108]), .Z(n13094) );
  AND U19641 ( .A(p_input[4108]), .B(p_input[34108]), .Z(n13093) );
  AND U19642 ( .A(n13095), .B(n13096), .Z(o[4107]) );
  AND U19643 ( .A(p_input[24107]), .B(p_input[14107]), .Z(n13096) );
  AND U19644 ( .A(p_input[4107]), .B(p_input[34107]), .Z(n13095) );
  AND U19645 ( .A(n13097), .B(n13098), .Z(o[4106]) );
  AND U19646 ( .A(p_input[24106]), .B(p_input[14106]), .Z(n13098) );
  AND U19647 ( .A(p_input[4106]), .B(p_input[34106]), .Z(n13097) );
  AND U19648 ( .A(n13099), .B(n13100), .Z(o[4105]) );
  AND U19649 ( .A(p_input[24105]), .B(p_input[14105]), .Z(n13100) );
  AND U19650 ( .A(p_input[4105]), .B(p_input[34105]), .Z(n13099) );
  AND U19651 ( .A(n13101), .B(n13102), .Z(o[4104]) );
  AND U19652 ( .A(p_input[24104]), .B(p_input[14104]), .Z(n13102) );
  AND U19653 ( .A(p_input[4104]), .B(p_input[34104]), .Z(n13101) );
  AND U19654 ( .A(n13103), .B(n13104), .Z(o[4103]) );
  AND U19655 ( .A(p_input[24103]), .B(p_input[14103]), .Z(n13104) );
  AND U19656 ( .A(p_input[4103]), .B(p_input[34103]), .Z(n13103) );
  AND U19657 ( .A(n13105), .B(n13106), .Z(o[4102]) );
  AND U19658 ( .A(p_input[24102]), .B(p_input[14102]), .Z(n13106) );
  AND U19659 ( .A(p_input[4102]), .B(p_input[34102]), .Z(n13105) );
  AND U19660 ( .A(n13107), .B(n13108), .Z(o[4101]) );
  AND U19661 ( .A(p_input[24101]), .B(p_input[14101]), .Z(n13108) );
  AND U19662 ( .A(p_input[4101]), .B(p_input[34101]), .Z(n13107) );
  AND U19663 ( .A(n13109), .B(n13110), .Z(o[4100]) );
  AND U19664 ( .A(p_input[24100]), .B(p_input[14100]), .Z(n13110) );
  AND U19665 ( .A(p_input[4100]), .B(p_input[34100]), .Z(n13109) );
  AND U19666 ( .A(n13111), .B(n13112), .Z(o[40]) );
  AND U19667 ( .A(p_input[20040]), .B(p_input[10040]), .Z(n13112) );
  AND U19668 ( .A(p_input[40]), .B(p_input[30040]), .Z(n13111) );
  AND U19669 ( .A(n13113), .B(n13114), .Z(o[409]) );
  AND U19670 ( .A(p_input[20409]), .B(p_input[10409]), .Z(n13114) );
  AND U19671 ( .A(p_input[409]), .B(p_input[30409]), .Z(n13113) );
  AND U19672 ( .A(n13115), .B(n13116), .Z(o[4099]) );
  AND U19673 ( .A(p_input[24099]), .B(p_input[14099]), .Z(n13116) );
  AND U19674 ( .A(p_input[4099]), .B(p_input[34099]), .Z(n13115) );
  AND U19675 ( .A(n13117), .B(n13118), .Z(o[4098]) );
  AND U19676 ( .A(p_input[24098]), .B(p_input[14098]), .Z(n13118) );
  AND U19677 ( .A(p_input[4098]), .B(p_input[34098]), .Z(n13117) );
  AND U19678 ( .A(n13119), .B(n13120), .Z(o[4097]) );
  AND U19679 ( .A(p_input[24097]), .B(p_input[14097]), .Z(n13120) );
  AND U19680 ( .A(p_input[4097]), .B(p_input[34097]), .Z(n13119) );
  AND U19681 ( .A(n13121), .B(n13122), .Z(o[4096]) );
  AND U19682 ( .A(p_input[24096]), .B(p_input[14096]), .Z(n13122) );
  AND U19683 ( .A(p_input[4096]), .B(p_input[34096]), .Z(n13121) );
  AND U19684 ( .A(n13123), .B(n13124), .Z(o[4095]) );
  AND U19685 ( .A(p_input[24095]), .B(p_input[14095]), .Z(n13124) );
  AND U19686 ( .A(p_input[4095]), .B(p_input[34095]), .Z(n13123) );
  AND U19687 ( .A(n13125), .B(n13126), .Z(o[4094]) );
  AND U19688 ( .A(p_input[24094]), .B(p_input[14094]), .Z(n13126) );
  AND U19689 ( .A(p_input[4094]), .B(p_input[34094]), .Z(n13125) );
  AND U19690 ( .A(n13127), .B(n13128), .Z(o[4093]) );
  AND U19691 ( .A(p_input[24093]), .B(p_input[14093]), .Z(n13128) );
  AND U19692 ( .A(p_input[4093]), .B(p_input[34093]), .Z(n13127) );
  AND U19693 ( .A(n13129), .B(n13130), .Z(o[4092]) );
  AND U19694 ( .A(p_input[24092]), .B(p_input[14092]), .Z(n13130) );
  AND U19695 ( .A(p_input[4092]), .B(p_input[34092]), .Z(n13129) );
  AND U19696 ( .A(n13131), .B(n13132), .Z(o[4091]) );
  AND U19697 ( .A(p_input[24091]), .B(p_input[14091]), .Z(n13132) );
  AND U19698 ( .A(p_input[4091]), .B(p_input[34091]), .Z(n13131) );
  AND U19699 ( .A(n13133), .B(n13134), .Z(o[4090]) );
  AND U19700 ( .A(p_input[24090]), .B(p_input[14090]), .Z(n13134) );
  AND U19701 ( .A(p_input[4090]), .B(p_input[34090]), .Z(n13133) );
  AND U19702 ( .A(n13135), .B(n13136), .Z(o[408]) );
  AND U19703 ( .A(p_input[20408]), .B(p_input[10408]), .Z(n13136) );
  AND U19704 ( .A(p_input[408]), .B(p_input[30408]), .Z(n13135) );
  AND U19705 ( .A(n13137), .B(n13138), .Z(o[4089]) );
  AND U19706 ( .A(p_input[24089]), .B(p_input[14089]), .Z(n13138) );
  AND U19707 ( .A(p_input[4089]), .B(p_input[34089]), .Z(n13137) );
  AND U19708 ( .A(n13139), .B(n13140), .Z(o[4088]) );
  AND U19709 ( .A(p_input[24088]), .B(p_input[14088]), .Z(n13140) );
  AND U19710 ( .A(p_input[4088]), .B(p_input[34088]), .Z(n13139) );
  AND U19711 ( .A(n13141), .B(n13142), .Z(o[4087]) );
  AND U19712 ( .A(p_input[24087]), .B(p_input[14087]), .Z(n13142) );
  AND U19713 ( .A(p_input[4087]), .B(p_input[34087]), .Z(n13141) );
  AND U19714 ( .A(n13143), .B(n13144), .Z(o[4086]) );
  AND U19715 ( .A(p_input[24086]), .B(p_input[14086]), .Z(n13144) );
  AND U19716 ( .A(p_input[4086]), .B(p_input[34086]), .Z(n13143) );
  AND U19717 ( .A(n13145), .B(n13146), .Z(o[4085]) );
  AND U19718 ( .A(p_input[24085]), .B(p_input[14085]), .Z(n13146) );
  AND U19719 ( .A(p_input[4085]), .B(p_input[34085]), .Z(n13145) );
  AND U19720 ( .A(n13147), .B(n13148), .Z(o[4084]) );
  AND U19721 ( .A(p_input[24084]), .B(p_input[14084]), .Z(n13148) );
  AND U19722 ( .A(p_input[4084]), .B(p_input[34084]), .Z(n13147) );
  AND U19723 ( .A(n13149), .B(n13150), .Z(o[4083]) );
  AND U19724 ( .A(p_input[24083]), .B(p_input[14083]), .Z(n13150) );
  AND U19725 ( .A(p_input[4083]), .B(p_input[34083]), .Z(n13149) );
  AND U19726 ( .A(n13151), .B(n13152), .Z(o[4082]) );
  AND U19727 ( .A(p_input[24082]), .B(p_input[14082]), .Z(n13152) );
  AND U19728 ( .A(p_input[4082]), .B(p_input[34082]), .Z(n13151) );
  AND U19729 ( .A(n13153), .B(n13154), .Z(o[4081]) );
  AND U19730 ( .A(p_input[24081]), .B(p_input[14081]), .Z(n13154) );
  AND U19731 ( .A(p_input[4081]), .B(p_input[34081]), .Z(n13153) );
  AND U19732 ( .A(n13155), .B(n13156), .Z(o[4080]) );
  AND U19733 ( .A(p_input[24080]), .B(p_input[14080]), .Z(n13156) );
  AND U19734 ( .A(p_input[4080]), .B(p_input[34080]), .Z(n13155) );
  AND U19735 ( .A(n13157), .B(n13158), .Z(o[407]) );
  AND U19736 ( .A(p_input[20407]), .B(p_input[10407]), .Z(n13158) );
  AND U19737 ( .A(p_input[407]), .B(p_input[30407]), .Z(n13157) );
  AND U19738 ( .A(n13159), .B(n13160), .Z(o[4079]) );
  AND U19739 ( .A(p_input[24079]), .B(p_input[14079]), .Z(n13160) );
  AND U19740 ( .A(p_input[4079]), .B(p_input[34079]), .Z(n13159) );
  AND U19741 ( .A(n13161), .B(n13162), .Z(o[4078]) );
  AND U19742 ( .A(p_input[24078]), .B(p_input[14078]), .Z(n13162) );
  AND U19743 ( .A(p_input[4078]), .B(p_input[34078]), .Z(n13161) );
  AND U19744 ( .A(n13163), .B(n13164), .Z(o[4077]) );
  AND U19745 ( .A(p_input[24077]), .B(p_input[14077]), .Z(n13164) );
  AND U19746 ( .A(p_input[4077]), .B(p_input[34077]), .Z(n13163) );
  AND U19747 ( .A(n13165), .B(n13166), .Z(o[4076]) );
  AND U19748 ( .A(p_input[24076]), .B(p_input[14076]), .Z(n13166) );
  AND U19749 ( .A(p_input[4076]), .B(p_input[34076]), .Z(n13165) );
  AND U19750 ( .A(n13167), .B(n13168), .Z(o[4075]) );
  AND U19751 ( .A(p_input[24075]), .B(p_input[14075]), .Z(n13168) );
  AND U19752 ( .A(p_input[4075]), .B(p_input[34075]), .Z(n13167) );
  AND U19753 ( .A(n13169), .B(n13170), .Z(o[4074]) );
  AND U19754 ( .A(p_input[24074]), .B(p_input[14074]), .Z(n13170) );
  AND U19755 ( .A(p_input[4074]), .B(p_input[34074]), .Z(n13169) );
  AND U19756 ( .A(n13171), .B(n13172), .Z(o[4073]) );
  AND U19757 ( .A(p_input[24073]), .B(p_input[14073]), .Z(n13172) );
  AND U19758 ( .A(p_input[4073]), .B(p_input[34073]), .Z(n13171) );
  AND U19759 ( .A(n13173), .B(n13174), .Z(o[4072]) );
  AND U19760 ( .A(p_input[24072]), .B(p_input[14072]), .Z(n13174) );
  AND U19761 ( .A(p_input[4072]), .B(p_input[34072]), .Z(n13173) );
  AND U19762 ( .A(n13175), .B(n13176), .Z(o[4071]) );
  AND U19763 ( .A(p_input[24071]), .B(p_input[14071]), .Z(n13176) );
  AND U19764 ( .A(p_input[4071]), .B(p_input[34071]), .Z(n13175) );
  AND U19765 ( .A(n13177), .B(n13178), .Z(o[4070]) );
  AND U19766 ( .A(p_input[24070]), .B(p_input[14070]), .Z(n13178) );
  AND U19767 ( .A(p_input[4070]), .B(p_input[34070]), .Z(n13177) );
  AND U19768 ( .A(n13179), .B(n13180), .Z(o[406]) );
  AND U19769 ( .A(p_input[20406]), .B(p_input[10406]), .Z(n13180) );
  AND U19770 ( .A(p_input[406]), .B(p_input[30406]), .Z(n13179) );
  AND U19771 ( .A(n13181), .B(n13182), .Z(o[4069]) );
  AND U19772 ( .A(p_input[24069]), .B(p_input[14069]), .Z(n13182) );
  AND U19773 ( .A(p_input[4069]), .B(p_input[34069]), .Z(n13181) );
  AND U19774 ( .A(n13183), .B(n13184), .Z(o[4068]) );
  AND U19775 ( .A(p_input[24068]), .B(p_input[14068]), .Z(n13184) );
  AND U19776 ( .A(p_input[4068]), .B(p_input[34068]), .Z(n13183) );
  AND U19777 ( .A(n13185), .B(n13186), .Z(o[4067]) );
  AND U19778 ( .A(p_input[24067]), .B(p_input[14067]), .Z(n13186) );
  AND U19779 ( .A(p_input[4067]), .B(p_input[34067]), .Z(n13185) );
  AND U19780 ( .A(n13187), .B(n13188), .Z(o[4066]) );
  AND U19781 ( .A(p_input[24066]), .B(p_input[14066]), .Z(n13188) );
  AND U19782 ( .A(p_input[4066]), .B(p_input[34066]), .Z(n13187) );
  AND U19783 ( .A(n13189), .B(n13190), .Z(o[4065]) );
  AND U19784 ( .A(p_input[24065]), .B(p_input[14065]), .Z(n13190) );
  AND U19785 ( .A(p_input[4065]), .B(p_input[34065]), .Z(n13189) );
  AND U19786 ( .A(n13191), .B(n13192), .Z(o[4064]) );
  AND U19787 ( .A(p_input[24064]), .B(p_input[14064]), .Z(n13192) );
  AND U19788 ( .A(p_input[4064]), .B(p_input[34064]), .Z(n13191) );
  AND U19789 ( .A(n13193), .B(n13194), .Z(o[4063]) );
  AND U19790 ( .A(p_input[24063]), .B(p_input[14063]), .Z(n13194) );
  AND U19791 ( .A(p_input[4063]), .B(p_input[34063]), .Z(n13193) );
  AND U19792 ( .A(n13195), .B(n13196), .Z(o[4062]) );
  AND U19793 ( .A(p_input[24062]), .B(p_input[14062]), .Z(n13196) );
  AND U19794 ( .A(p_input[4062]), .B(p_input[34062]), .Z(n13195) );
  AND U19795 ( .A(n13197), .B(n13198), .Z(o[4061]) );
  AND U19796 ( .A(p_input[24061]), .B(p_input[14061]), .Z(n13198) );
  AND U19797 ( .A(p_input[4061]), .B(p_input[34061]), .Z(n13197) );
  AND U19798 ( .A(n13199), .B(n13200), .Z(o[4060]) );
  AND U19799 ( .A(p_input[24060]), .B(p_input[14060]), .Z(n13200) );
  AND U19800 ( .A(p_input[4060]), .B(p_input[34060]), .Z(n13199) );
  AND U19801 ( .A(n13201), .B(n13202), .Z(o[405]) );
  AND U19802 ( .A(p_input[20405]), .B(p_input[10405]), .Z(n13202) );
  AND U19803 ( .A(p_input[405]), .B(p_input[30405]), .Z(n13201) );
  AND U19804 ( .A(n13203), .B(n13204), .Z(o[4059]) );
  AND U19805 ( .A(p_input[24059]), .B(p_input[14059]), .Z(n13204) );
  AND U19806 ( .A(p_input[4059]), .B(p_input[34059]), .Z(n13203) );
  AND U19807 ( .A(n13205), .B(n13206), .Z(o[4058]) );
  AND U19808 ( .A(p_input[24058]), .B(p_input[14058]), .Z(n13206) );
  AND U19809 ( .A(p_input[4058]), .B(p_input[34058]), .Z(n13205) );
  AND U19810 ( .A(n13207), .B(n13208), .Z(o[4057]) );
  AND U19811 ( .A(p_input[24057]), .B(p_input[14057]), .Z(n13208) );
  AND U19812 ( .A(p_input[4057]), .B(p_input[34057]), .Z(n13207) );
  AND U19813 ( .A(n13209), .B(n13210), .Z(o[4056]) );
  AND U19814 ( .A(p_input[24056]), .B(p_input[14056]), .Z(n13210) );
  AND U19815 ( .A(p_input[4056]), .B(p_input[34056]), .Z(n13209) );
  AND U19816 ( .A(n13211), .B(n13212), .Z(o[4055]) );
  AND U19817 ( .A(p_input[24055]), .B(p_input[14055]), .Z(n13212) );
  AND U19818 ( .A(p_input[4055]), .B(p_input[34055]), .Z(n13211) );
  AND U19819 ( .A(n13213), .B(n13214), .Z(o[4054]) );
  AND U19820 ( .A(p_input[24054]), .B(p_input[14054]), .Z(n13214) );
  AND U19821 ( .A(p_input[4054]), .B(p_input[34054]), .Z(n13213) );
  AND U19822 ( .A(n13215), .B(n13216), .Z(o[4053]) );
  AND U19823 ( .A(p_input[24053]), .B(p_input[14053]), .Z(n13216) );
  AND U19824 ( .A(p_input[4053]), .B(p_input[34053]), .Z(n13215) );
  AND U19825 ( .A(n13217), .B(n13218), .Z(o[4052]) );
  AND U19826 ( .A(p_input[24052]), .B(p_input[14052]), .Z(n13218) );
  AND U19827 ( .A(p_input[4052]), .B(p_input[34052]), .Z(n13217) );
  AND U19828 ( .A(n13219), .B(n13220), .Z(o[4051]) );
  AND U19829 ( .A(p_input[24051]), .B(p_input[14051]), .Z(n13220) );
  AND U19830 ( .A(p_input[4051]), .B(p_input[34051]), .Z(n13219) );
  AND U19831 ( .A(n13221), .B(n13222), .Z(o[4050]) );
  AND U19832 ( .A(p_input[24050]), .B(p_input[14050]), .Z(n13222) );
  AND U19833 ( .A(p_input[4050]), .B(p_input[34050]), .Z(n13221) );
  AND U19834 ( .A(n13223), .B(n13224), .Z(o[404]) );
  AND U19835 ( .A(p_input[20404]), .B(p_input[10404]), .Z(n13224) );
  AND U19836 ( .A(p_input[404]), .B(p_input[30404]), .Z(n13223) );
  AND U19837 ( .A(n13225), .B(n13226), .Z(o[4049]) );
  AND U19838 ( .A(p_input[24049]), .B(p_input[14049]), .Z(n13226) );
  AND U19839 ( .A(p_input[4049]), .B(p_input[34049]), .Z(n13225) );
  AND U19840 ( .A(n13227), .B(n13228), .Z(o[4048]) );
  AND U19841 ( .A(p_input[24048]), .B(p_input[14048]), .Z(n13228) );
  AND U19842 ( .A(p_input[4048]), .B(p_input[34048]), .Z(n13227) );
  AND U19843 ( .A(n13229), .B(n13230), .Z(o[4047]) );
  AND U19844 ( .A(p_input[24047]), .B(p_input[14047]), .Z(n13230) );
  AND U19845 ( .A(p_input[4047]), .B(p_input[34047]), .Z(n13229) );
  AND U19846 ( .A(n13231), .B(n13232), .Z(o[4046]) );
  AND U19847 ( .A(p_input[24046]), .B(p_input[14046]), .Z(n13232) );
  AND U19848 ( .A(p_input[4046]), .B(p_input[34046]), .Z(n13231) );
  AND U19849 ( .A(n13233), .B(n13234), .Z(o[4045]) );
  AND U19850 ( .A(p_input[24045]), .B(p_input[14045]), .Z(n13234) );
  AND U19851 ( .A(p_input[4045]), .B(p_input[34045]), .Z(n13233) );
  AND U19852 ( .A(n13235), .B(n13236), .Z(o[4044]) );
  AND U19853 ( .A(p_input[24044]), .B(p_input[14044]), .Z(n13236) );
  AND U19854 ( .A(p_input[4044]), .B(p_input[34044]), .Z(n13235) );
  AND U19855 ( .A(n13237), .B(n13238), .Z(o[4043]) );
  AND U19856 ( .A(p_input[24043]), .B(p_input[14043]), .Z(n13238) );
  AND U19857 ( .A(p_input[4043]), .B(p_input[34043]), .Z(n13237) );
  AND U19858 ( .A(n13239), .B(n13240), .Z(o[4042]) );
  AND U19859 ( .A(p_input[24042]), .B(p_input[14042]), .Z(n13240) );
  AND U19860 ( .A(p_input[4042]), .B(p_input[34042]), .Z(n13239) );
  AND U19861 ( .A(n13241), .B(n13242), .Z(o[4041]) );
  AND U19862 ( .A(p_input[24041]), .B(p_input[14041]), .Z(n13242) );
  AND U19863 ( .A(p_input[4041]), .B(p_input[34041]), .Z(n13241) );
  AND U19864 ( .A(n13243), .B(n13244), .Z(o[4040]) );
  AND U19865 ( .A(p_input[24040]), .B(p_input[14040]), .Z(n13244) );
  AND U19866 ( .A(p_input[4040]), .B(p_input[34040]), .Z(n13243) );
  AND U19867 ( .A(n13245), .B(n13246), .Z(o[403]) );
  AND U19868 ( .A(p_input[20403]), .B(p_input[10403]), .Z(n13246) );
  AND U19869 ( .A(p_input[403]), .B(p_input[30403]), .Z(n13245) );
  AND U19870 ( .A(n13247), .B(n13248), .Z(o[4039]) );
  AND U19871 ( .A(p_input[24039]), .B(p_input[14039]), .Z(n13248) );
  AND U19872 ( .A(p_input[4039]), .B(p_input[34039]), .Z(n13247) );
  AND U19873 ( .A(n13249), .B(n13250), .Z(o[4038]) );
  AND U19874 ( .A(p_input[24038]), .B(p_input[14038]), .Z(n13250) );
  AND U19875 ( .A(p_input[4038]), .B(p_input[34038]), .Z(n13249) );
  AND U19876 ( .A(n13251), .B(n13252), .Z(o[4037]) );
  AND U19877 ( .A(p_input[24037]), .B(p_input[14037]), .Z(n13252) );
  AND U19878 ( .A(p_input[4037]), .B(p_input[34037]), .Z(n13251) );
  AND U19879 ( .A(n13253), .B(n13254), .Z(o[4036]) );
  AND U19880 ( .A(p_input[24036]), .B(p_input[14036]), .Z(n13254) );
  AND U19881 ( .A(p_input[4036]), .B(p_input[34036]), .Z(n13253) );
  AND U19882 ( .A(n13255), .B(n13256), .Z(o[4035]) );
  AND U19883 ( .A(p_input[24035]), .B(p_input[14035]), .Z(n13256) );
  AND U19884 ( .A(p_input[4035]), .B(p_input[34035]), .Z(n13255) );
  AND U19885 ( .A(n13257), .B(n13258), .Z(o[4034]) );
  AND U19886 ( .A(p_input[24034]), .B(p_input[14034]), .Z(n13258) );
  AND U19887 ( .A(p_input[4034]), .B(p_input[34034]), .Z(n13257) );
  AND U19888 ( .A(n13259), .B(n13260), .Z(o[4033]) );
  AND U19889 ( .A(p_input[24033]), .B(p_input[14033]), .Z(n13260) );
  AND U19890 ( .A(p_input[4033]), .B(p_input[34033]), .Z(n13259) );
  AND U19891 ( .A(n13261), .B(n13262), .Z(o[4032]) );
  AND U19892 ( .A(p_input[24032]), .B(p_input[14032]), .Z(n13262) );
  AND U19893 ( .A(p_input[4032]), .B(p_input[34032]), .Z(n13261) );
  AND U19894 ( .A(n13263), .B(n13264), .Z(o[4031]) );
  AND U19895 ( .A(p_input[24031]), .B(p_input[14031]), .Z(n13264) );
  AND U19896 ( .A(p_input[4031]), .B(p_input[34031]), .Z(n13263) );
  AND U19897 ( .A(n13265), .B(n13266), .Z(o[4030]) );
  AND U19898 ( .A(p_input[24030]), .B(p_input[14030]), .Z(n13266) );
  AND U19899 ( .A(p_input[4030]), .B(p_input[34030]), .Z(n13265) );
  AND U19900 ( .A(n13267), .B(n13268), .Z(o[402]) );
  AND U19901 ( .A(p_input[20402]), .B(p_input[10402]), .Z(n13268) );
  AND U19902 ( .A(p_input[402]), .B(p_input[30402]), .Z(n13267) );
  AND U19903 ( .A(n13269), .B(n13270), .Z(o[4029]) );
  AND U19904 ( .A(p_input[24029]), .B(p_input[14029]), .Z(n13270) );
  AND U19905 ( .A(p_input[4029]), .B(p_input[34029]), .Z(n13269) );
  AND U19906 ( .A(n13271), .B(n13272), .Z(o[4028]) );
  AND U19907 ( .A(p_input[24028]), .B(p_input[14028]), .Z(n13272) );
  AND U19908 ( .A(p_input[4028]), .B(p_input[34028]), .Z(n13271) );
  AND U19909 ( .A(n13273), .B(n13274), .Z(o[4027]) );
  AND U19910 ( .A(p_input[24027]), .B(p_input[14027]), .Z(n13274) );
  AND U19911 ( .A(p_input[4027]), .B(p_input[34027]), .Z(n13273) );
  AND U19912 ( .A(n13275), .B(n13276), .Z(o[4026]) );
  AND U19913 ( .A(p_input[24026]), .B(p_input[14026]), .Z(n13276) );
  AND U19914 ( .A(p_input[4026]), .B(p_input[34026]), .Z(n13275) );
  AND U19915 ( .A(n13277), .B(n13278), .Z(o[4025]) );
  AND U19916 ( .A(p_input[24025]), .B(p_input[14025]), .Z(n13278) );
  AND U19917 ( .A(p_input[4025]), .B(p_input[34025]), .Z(n13277) );
  AND U19918 ( .A(n13279), .B(n13280), .Z(o[4024]) );
  AND U19919 ( .A(p_input[24024]), .B(p_input[14024]), .Z(n13280) );
  AND U19920 ( .A(p_input[4024]), .B(p_input[34024]), .Z(n13279) );
  AND U19921 ( .A(n13281), .B(n13282), .Z(o[4023]) );
  AND U19922 ( .A(p_input[24023]), .B(p_input[14023]), .Z(n13282) );
  AND U19923 ( .A(p_input[4023]), .B(p_input[34023]), .Z(n13281) );
  AND U19924 ( .A(n13283), .B(n13284), .Z(o[4022]) );
  AND U19925 ( .A(p_input[24022]), .B(p_input[14022]), .Z(n13284) );
  AND U19926 ( .A(p_input[4022]), .B(p_input[34022]), .Z(n13283) );
  AND U19927 ( .A(n13285), .B(n13286), .Z(o[4021]) );
  AND U19928 ( .A(p_input[24021]), .B(p_input[14021]), .Z(n13286) );
  AND U19929 ( .A(p_input[4021]), .B(p_input[34021]), .Z(n13285) );
  AND U19930 ( .A(n13287), .B(n13288), .Z(o[4020]) );
  AND U19931 ( .A(p_input[24020]), .B(p_input[14020]), .Z(n13288) );
  AND U19932 ( .A(p_input[4020]), .B(p_input[34020]), .Z(n13287) );
  AND U19933 ( .A(n13289), .B(n13290), .Z(o[401]) );
  AND U19934 ( .A(p_input[20401]), .B(p_input[10401]), .Z(n13290) );
  AND U19935 ( .A(p_input[401]), .B(p_input[30401]), .Z(n13289) );
  AND U19936 ( .A(n13291), .B(n13292), .Z(o[4019]) );
  AND U19937 ( .A(p_input[24019]), .B(p_input[14019]), .Z(n13292) );
  AND U19938 ( .A(p_input[4019]), .B(p_input[34019]), .Z(n13291) );
  AND U19939 ( .A(n13293), .B(n13294), .Z(o[4018]) );
  AND U19940 ( .A(p_input[24018]), .B(p_input[14018]), .Z(n13294) );
  AND U19941 ( .A(p_input[4018]), .B(p_input[34018]), .Z(n13293) );
  AND U19942 ( .A(n13295), .B(n13296), .Z(o[4017]) );
  AND U19943 ( .A(p_input[24017]), .B(p_input[14017]), .Z(n13296) );
  AND U19944 ( .A(p_input[4017]), .B(p_input[34017]), .Z(n13295) );
  AND U19945 ( .A(n13297), .B(n13298), .Z(o[4016]) );
  AND U19946 ( .A(p_input[24016]), .B(p_input[14016]), .Z(n13298) );
  AND U19947 ( .A(p_input[4016]), .B(p_input[34016]), .Z(n13297) );
  AND U19948 ( .A(n13299), .B(n13300), .Z(o[4015]) );
  AND U19949 ( .A(p_input[24015]), .B(p_input[14015]), .Z(n13300) );
  AND U19950 ( .A(p_input[4015]), .B(p_input[34015]), .Z(n13299) );
  AND U19951 ( .A(n13301), .B(n13302), .Z(o[4014]) );
  AND U19952 ( .A(p_input[24014]), .B(p_input[14014]), .Z(n13302) );
  AND U19953 ( .A(p_input[4014]), .B(p_input[34014]), .Z(n13301) );
  AND U19954 ( .A(n13303), .B(n13304), .Z(o[4013]) );
  AND U19955 ( .A(p_input[24013]), .B(p_input[14013]), .Z(n13304) );
  AND U19956 ( .A(p_input[4013]), .B(p_input[34013]), .Z(n13303) );
  AND U19957 ( .A(n13305), .B(n13306), .Z(o[4012]) );
  AND U19958 ( .A(p_input[24012]), .B(p_input[14012]), .Z(n13306) );
  AND U19959 ( .A(p_input[4012]), .B(p_input[34012]), .Z(n13305) );
  AND U19960 ( .A(n13307), .B(n13308), .Z(o[4011]) );
  AND U19961 ( .A(p_input[24011]), .B(p_input[14011]), .Z(n13308) );
  AND U19962 ( .A(p_input[4011]), .B(p_input[34011]), .Z(n13307) );
  AND U19963 ( .A(n13309), .B(n13310), .Z(o[4010]) );
  AND U19964 ( .A(p_input[24010]), .B(p_input[14010]), .Z(n13310) );
  AND U19965 ( .A(p_input[4010]), .B(p_input[34010]), .Z(n13309) );
  AND U19966 ( .A(n13311), .B(n13312), .Z(o[400]) );
  AND U19967 ( .A(p_input[20400]), .B(p_input[10400]), .Z(n13312) );
  AND U19968 ( .A(p_input[400]), .B(p_input[30400]), .Z(n13311) );
  AND U19969 ( .A(n13313), .B(n13314), .Z(o[4009]) );
  AND U19970 ( .A(p_input[24009]), .B(p_input[14009]), .Z(n13314) );
  AND U19971 ( .A(p_input[4009]), .B(p_input[34009]), .Z(n13313) );
  AND U19972 ( .A(n13315), .B(n13316), .Z(o[4008]) );
  AND U19973 ( .A(p_input[24008]), .B(p_input[14008]), .Z(n13316) );
  AND U19974 ( .A(p_input[4008]), .B(p_input[34008]), .Z(n13315) );
  AND U19975 ( .A(n13317), .B(n13318), .Z(o[4007]) );
  AND U19976 ( .A(p_input[24007]), .B(p_input[14007]), .Z(n13318) );
  AND U19977 ( .A(p_input[4007]), .B(p_input[34007]), .Z(n13317) );
  AND U19978 ( .A(n13319), .B(n13320), .Z(o[4006]) );
  AND U19979 ( .A(p_input[24006]), .B(p_input[14006]), .Z(n13320) );
  AND U19980 ( .A(p_input[4006]), .B(p_input[34006]), .Z(n13319) );
  AND U19981 ( .A(n13321), .B(n13322), .Z(o[4005]) );
  AND U19982 ( .A(p_input[24005]), .B(p_input[14005]), .Z(n13322) );
  AND U19983 ( .A(p_input[4005]), .B(p_input[34005]), .Z(n13321) );
  AND U19984 ( .A(n13323), .B(n13324), .Z(o[4004]) );
  AND U19985 ( .A(p_input[24004]), .B(p_input[14004]), .Z(n13324) );
  AND U19986 ( .A(p_input[4004]), .B(p_input[34004]), .Z(n13323) );
  AND U19987 ( .A(n13325), .B(n13326), .Z(o[4003]) );
  AND U19988 ( .A(p_input[24003]), .B(p_input[14003]), .Z(n13326) );
  AND U19989 ( .A(p_input[4003]), .B(p_input[34003]), .Z(n13325) );
  AND U19990 ( .A(n13327), .B(n13328), .Z(o[4002]) );
  AND U19991 ( .A(p_input[24002]), .B(p_input[14002]), .Z(n13328) );
  AND U19992 ( .A(p_input[4002]), .B(p_input[34002]), .Z(n13327) );
  AND U19993 ( .A(n13329), .B(n13330), .Z(o[4001]) );
  AND U19994 ( .A(p_input[24001]), .B(p_input[14001]), .Z(n13330) );
  AND U19995 ( .A(p_input[4001]), .B(p_input[34001]), .Z(n13329) );
  AND U19996 ( .A(n13331), .B(n13332), .Z(o[4000]) );
  AND U19997 ( .A(p_input[24000]), .B(p_input[14000]), .Z(n13332) );
  AND U19998 ( .A(p_input[4000]), .B(p_input[34000]), .Z(n13331) );
  AND U19999 ( .A(n13333), .B(n13334), .Z(o[3]) );
  AND U20000 ( .A(p_input[20003]), .B(p_input[10003]), .Z(n13334) );
  AND U20001 ( .A(p_input[3]), .B(p_input[30003]), .Z(n13333) );
  AND U20002 ( .A(n13335), .B(n13336), .Z(o[39]) );
  AND U20003 ( .A(p_input[20039]), .B(p_input[10039]), .Z(n13336) );
  AND U20004 ( .A(p_input[39]), .B(p_input[30039]), .Z(n13335) );
  AND U20005 ( .A(n13337), .B(n13338), .Z(o[399]) );
  AND U20006 ( .A(p_input[20399]), .B(p_input[10399]), .Z(n13338) );
  AND U20007 ( .A(p_input[399]), .B(p_input[30399]), .Z(n13337) );
  AND U20008 ( .A(n13339), .B(n13340), .Z(o[3999]) );
  AND U20009 ( .A(p_input[23999]), .B(p_input[13999]), .Z(n13340) );
  AND U20010 ( .A(p_input[3999]), .B(p_input[33999]), .Z(n13339) );
  AND U20011 ( .A(n13341), .B(n13342), .Z(o[3998]) );
  AND U20012 ( .A(p_input[23998]), .B(p_input[13998]), .Z(n13342) );
  AND U20013 ( .A(p_input[3998]), .B(p_input[33998]), .Z(n13341) );
  AND U20014 ( .A(n13343), .B(n13344), .Z(o[3997]) );
  AND U20015 ( .A(p_input[23997]), .B(p_input[13997]), .Z(n13344) );
  AND U20016 ( .A(p_input[3997]), .B(p_input[33997]), .Z(n13343) );
  AND U20017 ( .A(n13345), .B(n13346), .Z(o[3996]) );
  AND U20018 ( .A(p_input[23996]), .B(p_input[13996]), .Z(n13346) );
  AND U20019 ( .A(p_input[3996]), .B(p_input[33996]), .Z(n13345) );
  AND U20020 ( .A(n13347), .B(n13348), .Z(o[3995]) );
  AND U20021 ( .A(p_input[23995]), .B(p_input[13995]), .Z(n13348) );
  AND U20022 ( .A(p_input[3995]), .B(p_input[33995]), .Z(n13347) );
  AND U20023 ( .A(n13349), .B(n13350), .Z(o[3994]) );
  AND U20024 ( .A(p_input[23994]), .B(p_input[13994]), .Z(n13350) );
  AND U20025 ( .A(p_input[3994]), .B(p_input[33994]), .Z(n13349) );
  AND U20026 ( .A(n13351), .B(n13352), .Z(o[3993]) );
  AND U20027 ( .A(p_input[23993]), .B(p_input[13993]), .Z(n13352) );
  AND U20028 ( .A(p_input[3993]), .B(p_input[33993]), .Z(n13351) );
  AND U20029 ( .A(n13353), .B(n13354), .Z(o[3992]) );
  AND U20030 ( .A(p_input[23992]), .B(p_input[13992]), .Z(n13354) );
  AND U20031 ( .A(p_input[3992]), .B(p_input[33992]), .Z(n13353) );
  AND U20032 ( .A(n13355), .B(n13356), .Z(o[3991]) );
  AND U20033 ( .A(p_input[23991]), .B(p_input[13991]), .Z(n13356) );
  AND U20034 ( .A(p_input[3991]), .B(p_input[33991]), .Z(n13355) );
  AND U20035 ( .A(n13357), .B(n13358), .Z(o[3990]) );
  AND U20036 ( .A(p_input[23990]), .B(p_input[13990]), .Z(n13358) );
  AND U20037 ( .A(p_input[3990]), .B(p_input[33990]), .Z(n13357) );
  AND U20038 ( .A(n13359), .B(n13360), .Z(o[398]) );
  AND U20039 ( .A(p_input[20398]), .B(p_input[10398]), .Z(n13360) );
  AND U20040 ( .A(p_input[398]), .B(p_input[30398]), .Z(n13359) );
  AND U20041 ( .A(n13361), .B(n13362), .Z(o[3989]) );
  AND U20042 ( .A(p_input[23989]), .B(p_input[13989]), .Z(n13362) );
  AND U20043 ( .A(p_input[3989]), .B(p_input[33989]), .Z(n13361) );
  AND U20044 ( .A(n13363), .B(n13364), .Z(o[3988]) );
  AND U20045 ( .A(p_input[23988]), .B(p_input[13988]), .Z(n13364) );
  AND U20046 ( .A(p_input[3988]), .B(p_input[33988]), .Z(n13363) );
  AND U20047 ( .A(n13365), .B(n13366), .Z(o[3987]) );
  AND U20048 ( .A(p_input[23987]), .B(p_input[13987]), .Z(n13366) );
  AND U20049 ( .A(p_input[3987]), .B(p_input[33987]), .Z(n13365) );
  AND U20050 ( .A(n13367), .B(n13368), .Z(o[3986]) );
  AND U20051 ( .A(p_input[23986]), .B(p_input[13986]), .Z(n13368) );
  AND U20052 ( .A(p_input[3986]), .B(p_input[33986]), .Z(n13367) );
  AND U20053 ( .A(n13369), .B(n13370), .Z(o[3985]) );
  AND U20054 ( .A(p_input[23985]), .B(p_input[13985]), .Z(n13370) );
  AND U20055 ( .A(p_input[3985]), .B(p_input[33985]), .Z(n13369) );
  AND U20056 ( .A(n13371), .B(n13372), .Z(o[3984]) );
  AND U20057 ( .A(p_input[23984]), .B(p_input[13984]), .Z(n13372) );
  AND U20058 ( .A(p_input[3984]), .B(p_input[33984]), .Z(n13371) );
  AND U20059 ( .A(n13373), .B(n13374), .Z(o[3983]) );
  AND U20060 ( .A(p_input[23983]), .B(p_input[13983]), .Z(n13374) );
  AND U20061 ( .A(p_input[3983]), .B(p_input[33983]), .Z(n13373) );
  AND U20062 ( .A(n13375), .B(n13376), .Z(o[3982]) );
  AND U20063 ( .A(p_input[23982]), .B(p_input[13982]), .Z(n13376) );
  AND U20064 ( .A(p_input[3982]), .B(p_input[33982]), .Z(n13375) );
  AND U20065 ( .A(n13377), .B(n13378), .Z(o[3981]) );
  AND U20066 ( .A(p_input[23981]), .B(p_input[13981]), .Z(n13378) );
  AND U20067 ( .A(p_input[3981]), .B(p_input[33981]), .Z(n13377) );
  AND U20068 ( .A(n13379), .B(n13380), .Z(o[3980]) );
  AND U20069 ( .A(p_input[23980]), .B(p_input[13980]), .Z(n13380) );
  AND U20070 ( .A(p_input[3980]), .B(p_input[33980]), .Z(n13379) );
  AND U20071 ( .A(n13381), .B(n13382), .Z(o[397]) );
  AND U20072 ( .A(p_input[20397]), .B(p_input[10397]), .Z(n13382) );
  AND U20073 ( .A(p_input[397]), .B(p_input[30397]), .Z(n13381) );
  AND U20074 ( .A(n13383), .B(n13384), .Z(o[3979]) );
  AND U20075 ( .A(p_input[23979]), .B(p_input[13979]), .Z(n13384) );
  AND U20076 ( .A(p_input[3979]), .B(p_input[33979]), .Z(n13383) );
  AND U20077 ( .A(n13385), .B(n13386), .Z(o[3978]) );
  AND U20078 ( .A(p_input[23978]), .B(p_input[13978]), .Z(n13386) );
  AND U20079 ( .A(p_input[3978]), .B(p_input[33978]), .Z(n13385) );
  AND U20080 ( .A(n13387), .B(n13388), .Z(o[3977]) );
  AND U20081 ( .A(p_input[23977]), .B(p_input[13977]), .Z(n13388) );
  AND U20082 ( .A(p_input[3977]), .B(p_input[33977]), .Z(n13387) );
  AND U20083 ( .A(n13389), .B(n13390), .Z(o[3976]) );
  AND U20084 ( .A(p_input[23976]), .B(p_input[13976]), .Z(n13390) );
  AND U20085 ( .A(p_input[3976]), .B(p_input[33976]), .Z(n13389) );
  AND U20086 ( .A(n13391), .B(n13392), .Z(o[3975]) );
  AND U20087 ( .A(p_input[23975]), .B(p_input[13975]), .Z(n13392) );
  AND U20088 ( .A(p_input[3975]), .B(p_input[33975]), .Z(n13391) );
  AND U20089 ( .A(n13393), .B(n13394), .Z(o[3974]) );
  AND U20090 ( .A(p_input[23974]), .B(p_input[13974]), .Z(n13394) );
  AND U20091 ( .A(p_input[3974]), .B(p_input[33974]), .Z(n13393) );
  AND U20092 ( .A(n13395), .B(n13396), .Z(o[3973]) );
  AND U20093 ( .A(p_input[23973]), .B(p_input[13973]), .Z(n13396) );
  AND U20094 ( .A(p_input[3973]), .B(p_input[33973]), .Z(n13395) );
  AND U20095 ( .A(n13397), .B(n13398), .Z(o[3972]) );
  AND U20096 ( .A(p_input[23972]), .B(p_input[13972]), .Z(n13398) );
  AND U20097 ( .A(p_input[3972]), .B(p_input[33972]), .Z(n13397) );
  AND U20098 ( .A(n13399), .B(n13400), .Z(o[3971]) );
  AND U20099 ( .A(p_input[23971]), .B(p_input[13971]), .Z(n13400) );
  AND U20100 ( .A(p_input[3971]), .B(p_input[33971]), .Z(n13399) );
  AND U20101 ( .A(n13401), .B(n13402), .Z(o[3970]) );
  AND U20102 ( .A(p_input[23970]), .B(p_input[13970]), .Z(n13402) );
  AND U20103 ( .A(p_input[3970]), .B(p_input[33970]), .Z(n13401) );
  AND U20104 ( .A(n13403), .B(n13404), .Z(o[396]) );
  AND U20105 ( .A(p_input[20396]), .B(p_input[10396]), .Z(n13404) );
  AND U20106 ( .A(p_input[396]), .B(p_input[30396]), .Z(n13403) );
  AND U20107 ( .A(n13405), .B(n13406), .Z(o[3969]) );
  AND U20108 ( .A(p_input[23969]), .B(p_input[13969]), .Z(n13406) );
  AND U20109 ( .A(p_input[3969]), .B(p_input[33969]), .Z(n13405) );
  AND U20110 ( .A(n13407), .B(n13408), .Z(o[3968]) );
  AND U20111 ( .A(p_input[23968]), .B(p_input[13968]), .Z(n13408) );
  AND U20112 ( .A(p_input[3968]), .B(p_input[33968]), .Z(n13407) );
  AND U20113 ( .A(n13409), .B(n13410), .Z(o[3967]) );
  AND U20114 ( .A(p_input[23967]), .B(p_input[13967]), .Z(n13410) );
  AND U20115 ( .A(p_input[3967]), .B(p_input[33967]), .Z(n13409) );
  AND U20116 ( .A(n13411), .B(n13412), .Z(o[3966]) );
  AND U20117 ( .A(p_input[23966]), .B(p_input[13966]), .Z(n13412) );
  AND U20118 ( .A(p_input[3966]), .B(p_input[33966]), .Z(n13411) );
  AND U20119 ( .A(n13413), .B(n13414), .Z(o[3965]) );
  AND U20120 ( .A(p_input[23965]), .B(p_input[13965]), .Z(n13414) );
  AND U20121 ( .A(p_input[3965]), .B(p_input[33965]), .Z(n13413) );
  AND U20122 ( .A(n13415), .B(n13416), .Z(o[3964]) );
  AND U20123 ( .A(p_input[23964]), .B(p_input[13964]), .Z(n13416) );
  AND U20124 ( .A(p_input[3964]), .B(p_input[33964]), .Z(n13415) );
  AND U20125 ( .A(n13417), .B(n13418), .Z(o[3963]) );
  AND U20126 ( .A(p_input[23963]), .B(p_input[13963]), .Z(n13418) );
  AND U20127 ( .A(p_input[3963]), .B(p_input[33963]), .Z(n13417) );
  AND U20128 ( .A(n13419), .B(n13420), .Z(o[3962]) );
  AND U20129 ( .A(p_input[23962]), .B(p_input[13962]), .Z(n13420) );
  AND U20130 ( .A(p_input[3962]), .B(p_input[33962]), .Z(n13419) );
  AND U20131 ( .A(n13421), .B(n13422), .Z(o[3961]) );
  AND U20132 ( .A(p_input[23961]), .B(p_input[13961]), .Z(n13422) );
  AND U20133 ( .A(p_input[3961]), .B(p_input[33961]), .Z(n13421) );
  AND U20134 ( .A(n13423), .B(n13424), .Z(o[3960]) );
  AND U20135 ( .A(p_input[23960]), .B(p_input[13960]), .Z(n13424) );
  AND U20136 ( .A(p_input[3960]), .B(p_input[33960]), .Z(n13423) );
  AND U20137 ( .A(n13425), .B(n13426), .Z(o[395]) );
  AND U20138 ( .A(p_input[20395]), .B(p_input[10395]), .Z(n13426) );
  AND U20139 ( .A(p_input[395]), .B(p_input[30395]), .Z(n13425) );
  AND U20140 ( .A(n13427), .B(n13428), .Z(o[3959]) );
  AND U20141 ( .A(p_input[23959]), .B(p_input[13959]), .Z(n13428) );
  AND U20142 ( .A(p_input[3959]), .B(p_input[33959]), .Z(n13427) );
  AND U20143 ( .A(n13429), .B(n13430), .Z(o[3958]) );
  AND U20144 ( .A(p_input[23958]), .B(p_input[13958]), .Z(n13430) );
  AND U20145 ( .A(p_input[3958]), .B(p_input[33958]), .Z(n13429) );
  AND U20146 ( .A(n13431), .B(n13432), .Z(o[3957]) );
  AND U20147 ( .A(p_input[23957]), .B(p_input[13957]), .Z(n13432) );
  AND U20148 ( .A(p_input[3957]), .B(p_input[33957]), .Z(n13431) );
  AND U20149 ( .A(n13433), .B(n13434), .Z(o[3956]) );
  AND U20150 ( .A(p_input[23956]), .B(p_input[13956]), .Z(n13434) );
  AND U20151 ( .A(p_input[3956]), .B(p_input[33956]), .Z(n13433) );
  AND U20152 ( .A(n13435), .B(n13436), .Z(o[3955]) );
  AND U20153 ( .A(p_input[23955]), .B(p_input[13955]), .Z(n13436) );
  AND U20154 ( .A(p_input[3955]), .B(p_input[33955]), .Z(n13435) );
  AND U20155 ( .A(n13437), .B(n13438), .Z(o[3954]) );
  AND U20156 ( .A(p_input[23954]), .B(p_input[13954]), .Z(n13438) );
  AND U20157 ( .A(p_input[3954]), .B(p_input[33954]), .Z(n13437) );
  AND U20158 ( .A(n13439), .B(n13440), .Z(o[3953]) );
  AND U20159 ( .A(p_input[23953]), .B(p_input[13953]), .Z(n13440) );
  AND U20160 ( .A(p_input[3953]), .B(p_input[33953]), .Z(n13439) );
  AND U20161 ( .A(n13441), .B(n13442), .Z(o[3952]) );
  AND U20162 ( .A(p_input[23952]), .B(p_input[13952]), .Z(n13442) );
  AND U20163 ( .A(p_input[3952]), .B(p_input[33952]), .Z(n13441) );
  AND U20164 ( .A(n13443), .B(n13444), .Z(o[3951]) );
  AND U20165 ( .A(p_input[23951]), .B(p_input[13951]), .Z(n13444) );
  AND U20166 ( .A(p_input[3951]), .B(p_input[33951]), .Z(n13443) );
  AND U20167 ( .A(n13445), .B(n13446), .Z(o[3950]) );
  AND U20168 ( .A(p_input[23950]), .B(p_input[13950]), .Z(n13446) );
  AND U20169 ( .A(p_input[3950]), .B(p_input[33950]), .Z(n13445) );
  AND U20170 ( .A(n13447), .B(n13448), .Z(o[394]) );
  AND U20171 ( .A(p_input[20394]), .B(p_input[10394]), .Z(n13448) );
  AND U20172 ( .A(p_input[394]), .B(p_input[30394]), .Z(n13447) );
  AND U20173 ( .A(n13449), .B(n13450), .Z(o[3949]) );
  AND U20174 ( .A(p_input[23949]), .B(p_input[13949]), .Z(n13450) );
  AND U20175 ( .A(p_input[3949]), .B(p_input[33949]), .Z(n13449) );
  AND U20176 ( .A(n13451), .B(n13452), .Z(o[3948]) );
  AND U20177 ( .A(p_input[23948]), .B(p_input[13948]), .Z(n13452) );
  AND U20178 ( .A(p_input[3948]), .B(p_input[33948]), .Z(n13451) );
  AND U20179 ( .A(n13453), .B(n13454), .Z(o[3947]) );
  AND U20180 ( .A(p_input[23947]), .B(p_input[13947]), .Z(n13454) );
  AND U20181 ( .A(p_input[3947]), .B(p_input[33947]), .Z(n13453) );
  AND U20182 ( .A(n13455), .B(n13456), .Z(o[3946]) );
  AND U20183 ( .A(p_input[23946]), .B(p_input[13946]), .Z(n13456) );
  AND U20184 ( .A(p_input[3946]), .B(p_input[33946]), .Z(n13455) );
  AND U20185 ( .A(n13457), .B(n13458), .Z(o[3945]) );
  AND U20186 ( .A(p_input[23945]), .B(p_input[13945]), .Z(n13458) );
  AND U20187 ( .A(p_input[3945]), .B(p_input[33945]), .Z(n13457) );
  AND U20188 ( .A(n13459), .B(n13460), .Z(o[3944]) );
  AND U20189 ( .A(p_input[23944]), .B(p_input[13944]), .Z(n13460) );
  AND U20190 ( .A(p_input[3944]), .B(p_input[33944]), .Z(n13459) );
  AND U20191 ( .A(n13461), .B(n13462), .Z(o[3943]) );
  AND U20192 ( .A(p_input[23943]), .B(p_input[13943]), .Z(n13462) );
  AND U20193 ( .A(p_input[3943]), .B(p_input[33943]), .Z(n13461) );
  AND U20194 ( .A(n13463), .B(n13464), .Z(o[3942]) );
  AND U20195 ( .A(p_input[23942]), .B(p_input[13942]), .Z(n13464) );
  AND U20196 ( .A(p_input[3942]), .B(p_input[33942]), .Z(n13463) );
  AND U20197 ( .A(n13465), .B(n13466), .Z(o[3941]) );
  AND U20198 ( .A(p_input[23941]), .B(p_input[13941]), .Z(n13466) );
  AND U20199 ( .A(p_input[3941]), .B(p_input[33941]), .Z(n13465) );
  AND U20200 ( .A(n13467), .B(n13468), .Z(o[3940]) );
  AND U20201 ( .A(p_input[23940]), .B(p_input[13940]), .Z(n13468) );
  AND U20202 ( .A(p_input[3940]), .B(p_input[33940]), .Z(n13467) );
  AND U20203 ( .A(n13469), .B(n13470), .Z(o[393]) );
  AND U20204 ( .A(p_input[20393]), .B(p_input[10393]), .Z(n13470) );
  AND U20205 ( .A(p_input[393]), .B(p_input[30393]), .Z(n13469) );
  AND U20206 ( .A(n13471), .B(n13472), .Z(o[3939]) );
  AND U20207 ( .A(p_input[23939]), .B(p_input[13939]), .Z(n13472) );
  AND U20208 ( .A(p_input[3939]), .B(p_input[33939]), .Z(n13471) );
  AND U20209 ( .A(n13473), .B(n13474), .Z(o[3938]) );
  AND U20210 ( .A(p_input[23938]), .B(p_input[13938]), .Z(n13474) );
  AND U20211 ( .A(p_input[3938]), .B(p_input[33938]), .Z(n13473) );
  AND U20212 ( .A(n13475), .B(n13476), .Z(o[3937]) );
  AND U20213 ( .A(p_input[23937]), .B(p_input[13937]), .Z(n13476) );
  AND U20214 ( .A(p_input[3937]), .B(p_input[33937]), .Z(n13475) );
  AND U20215 ( .A(n13477), .B(n13478), .Z(o[3936]) );
  AND U20216 ( .A(p_input[23936]), .B(p_input[13936]), .Z(n13478) );
  AND U20217 ( .A(p_input[3936]), .B(p_input[33936]), .Z(n13477) );
  AND U20218 ( .A(n13479), .B(n13480), .Z(o[3935]) );
  AND U20219 ( .A(p_input[23935]), .B(p_input[13935]), .Z(n13480) );
  AND U20220 ( .A(p_input[3935]), .B(p_input[33935]), .Z(n13479) );
  AND U20221 ( .A(n13481), .B(n13482), .Z(o[3934]) );
  AND U20222 ( .A(p_input[23934]), .B(p_input[13934]), .Z(n13482) );
  AND U20223 ( .A(p_input[3934]), .B(p_input[33934]), .Z(n13481) );
  AND U20224 ( .A(n13483), .B(n13484), .Z(o[3933]) );
  AND U20225 ( .A(p_input[23933]), .B(p_input[13933]), .Z(n13484) );
  AND U20226 ( .A(p_input[3933]), .B(p_input[33933]), .Z(n13483) );
  AND U20227 ( .A(n13485), .B(n13486), .Z(o[3932]) );
  AND U20228 ( .A(p_input[23932]), .B(p_input[13932]), .Z(n13486) );
  AND U20229 ( .A(p_input[3932]), .B(p_input[33932]), .Z(n13485) );
  AND U20230 ( .A(n13487), .B(n13488), .Z(o[3931]) );
  AND U20231 ( .A(p_input[23931]), .B(p_input[13931]), .Z(n13488) );
  AND U20232 ( .A(p_input[3931]), .B(p_input[33931]), .Z(n13487) );
  AND U20233 ( .A(n13489), .B(n13490), .Z(o[3930]) );
  AND U20234 ( .A(p_input[23930]), .B(p_input[13930]), .Z(n13490) );
  AND U20235 ( .A(p_input[3930]), .B(p_input[33930]), .Z(n13489) );
  AND U20236 ( .A(n13491), .B(n13492), .Z(o[392]) );
  AND U20237 ( .A(p_input[20392]), .B(p_input[10392]), .Z(n13492) );
  AND U20238 ( .A(p_input[392]), .B(p_input[30392]), .Z(n13491) );
  AND U20239 ( .A(n13493), .B(n13494), .Z(o[3929]) );
  AND U20240 ( .A(p_input[23929]), .B(p_input[13929]), .Z(n13494) );
  AND U20241 ( .A(p_input[3929]), .B(p_input[33929]), .Z(n13493) );
  AND U20242 ( .A(n13495), .B(n13496), .Z(o[3928]) );
  AND U20243 ( .A(p_input[23928]), .B(p_input[13928]), .Z(n13496) );
  AND U20244 ( .A(p_input[3928]), .B(p_input[33928]), .Z(n13495) );
  AND U20245 ( .A(n13497), .B(n13498), .Z(o[3927]) );
  AND U20246 ( .A(p_input[23927]), .B(p_input[13927]), .Z(n13498) );
  AND U20247 ( .A(p_input[3927]), .B(p_input[33927]), .Z(n13497) );
  AND U20248 ( .A(n13499), .B(n13500), .Z(o[3926]) );
  AND U20249 ( .A(p_input[23926]), .B(p_input[13926]), .Z(n13500) );
  AND U20250 ( .A(p_input[3926]), .B(p_input[33926]), .Z(n13499) );
  AND U20251 ( .A(n13501), .B(n13502), .Z(o[3925]) );
  AND U20252 ( .A(p_input[23925]), .B(p_input[13925]), .Z(n13502) );
  AND U20253 ( .A(p_input[3925]), .B(p_input[33925]), .Z(n13501) );
  AND U20254 ( .A(n13503), .B(n13504), .Z(o[3924]) );
  AND U20255 ( .A(p_input[23924]), .B(p_input[13924]), .Z(n13504) );
  AND U20256 ( .A(p_input[3924]), .B(p_input[33924]), .Z(n13503) );
  AND U20257 ( .A(n13505), .B(n13506), .Z(o[3923]) );
  AND U20258 ( .A(p_input[23923]), .B(p_input[13923]), .Z(n13506) );
  AND U20259 ( .A(p_input[3923]), .B(p_input[33923]), .Z(n13505) );
  AND U20260 ( .A(n13507), .B(n13508), .Z(o[3922]) );
  AND U20261 ( .A(p_input[23922]), .B(p_input[13922]), .Z(n13508) );
  AND U20262 ( .A(p_input[3922]), .B(p_input[33922]), .Z(n13507) );
  AND U20263 ( .A(n13509), .B(n13510), .Z(o[3921]) );
  AND U20264 ( .A(p_input[23921]), .B(p_input[13921]), .Z(n13510) );
  AND U20265 ( .A(p_input[3921]), .B(p_input[33921]), .Z(n13509) );
  AND U20266 ( .A(n13511), .B(n13512), .Z(o[3920]) );
  AND U20267 ( .A(p_input[23920]), .B(p_input[13920]), .Z(n13512) );
  AND U20268 ( .A(p_input[3920]), .B(p_input[33920]), .Z(n13511) );
  AND U20269 ( .A(n13513), .B(n13514), .Z(o[391]) );
  AND U20270 ( .A(p_input[20391]), .B(p_input[10391]), .Z(n13514) );
  AND U20271 ( .A(p_input[391]), .B(p_input[30391]), .Z(n13513) );
  AND U20272 ( .A(n13515), .B(n13516), .Z(o[3919]) );
  AND U20273 ( .A(p_input[23919]), .B(p_input[13919]), .Z(n13516) );
  AND U20274 ( .A(p_input[3919]), .B(p_input[33919]), .Z(n13515) );
  AND U20275 ( .A(n13517), .B(n13518), .Z(o[3918]) );
  AND U20276 ( .A(p_input[23918]), .B(p_input[13918]), .Z(n13518) );
  AND U20277 ( .A(p_input[3918]), .B(p_input[33918]), .Z(n13517) );
  AND U20278 ( .A(n13519), .B(n13520), .Z(o[3917]) );
  AND U20279 ( .A(p_input[23917]), .B(p_input[13917]), .Z(n13520) );
  AND U20280 ( .A(p_input[3917]), .B(p_input[33917]), .Z(n13519) );
  AND U20281 ( .A(n13521), .B(n13522), .Z(o[3916]) );
  AND U20282 ( .A(p_input[23916]), .B(p_input[13916]), .Z(n13522) );
  AND U20283 ( .A(p_input[3916]), .B(p_input[33916]), .Z(n13521) );
  AND U20284 ( .A(n13523), .B(n13524), .Z(o[3915]) );
  AND U20285 ( .A(p_input[23915]), .B(p_input[13915]), .Z(n13524) );
  AND U20286 ( .A(p_input[3915]), .B(p_input[33915]), .Z(n13523) );
  AND U20287 ( .A(n13525), .B(n13526), .Z(o[3914]) );
  AND U20288 ( .A(p_input[23914]), .B(p_input[13914]), .Z(n13526) );
  AND U20289 ( .A(p_input[3914]), .B(p_input[33914]), .Z(n13525) );
  AND U20290 ( .A(n13527), .B(n13528), .Z(o[3913]) );
  AND U20291 ( .A(p_input[23913]), .B(p_input[13913]), .Z(n13528) );
  AND U20292 ( .A(p_input[3913]), .B(p_input[33913]), .Z(n13527) );
  AND U20293 ( .A(n13529), .B(n13530), .Z(o[3912]) );
  AND U20294 ( .A(p_input[23912]), .B(p_input[13912]), .Z(n13530) );
  AND U20295 ( .A(p_input[3912]), .B(p_input[33912]), .Z(n13529) );
  AND U20296 ( .A(n13531), .B(n13532), .Z(o[3911]) );
  AND U20297 ( .A(p_input[23911]), .B(p_input[13911]), .Z(n13532) );
  AND U20298 ( .A(p_input[3911]), .B(p_input[33911]), .Z(n13531) );
  AND U20299 ( .A(n13533), .B(n13534), .Z(o[3910]) );
  AND U20300 ( .A(p_input[23910]), .B(p_input[13910]), .Z(n13534) );
  AND U20301 ( .A(p_input[3910]), .B(p_input[33910]), .Z(n13533) );
  AND U20302 ( .A(n13535), .B(n13536), .Z(o[390]) );
  AND U20303 ( .A(p_input[20390]), .B(p_input[10390]), .Z(n13536) );
  AND U20304 ( .A(p_input[390]), .B(p_input[30390]), .Z(n13535) );
  AND U20305 ( .A(n13537), .B(n13538), .Z(o[3909]) );
  AND U20306 ( .A(p_input[23909]), .B(p_input[13909]), .Z(n13538) );
  AND U20307 ( .A(p_input[3909]), .B(p_input[33909]), .Z(n13537) );
  AND U20308 ( .A(n13539), .B(n13540), .Z(o[3908]) );
  AND U20309 ( .A(p_input[23908]), .B(p_input[13908]), .Z(n13540) );
  AND U20310 ( .A(p_input[3908]), .B(p_input[33908]), .Z(n13539) );
  AND U20311 ( .A(n13541), .B(n13542), .Z(o[3907]) );
  AND U20312 ( .A(p_input[23907]), .B(p_input[13907]), .Z(n13542) );
  AND U20313 ( .A(p_input[3907]), .B(p_input[33907]), .Z(n13541) );
  AND U20314 ( .A(n13543), .B(n13544), .Z(o[3906]) );
  AND U20315 ( .A(p_input[23906]), .B(p_input[13906]), .Z(n13544) );
  AND U20316 ( .A(p_input[3906]), .B(p_input[33906]), .Z(n13543) );
  AND U20317 ( .A(n13545), .B(n13546), .Z(o[3905]) );
  AND U20318 ( .A(p_input[23905]), .B(p_input[13905]), .Z(n13546) );
  AND U20319 ( .A(p_input[3905]), .B(p_input[33905]), .Z(n13545) );
  AND U20320 ( .A(n13547), .B(n13548), .Z(o[3904]) );
  AND U20321 ( .A(p_input[23904]), .B(p_input[13904]), .Z(n13548) );
  AND U20322 ( .A(p_input[3904]), .B(p_input[33904]), .Z(n13547) );
  AND U20323 ( .A(n13549), .B(n13550), .Z(o[3903]) );
  AND U20324 ( .A(p_input[23903]), .B(p_input[13903]), .Z(n13550) );
  AND U20325 ( .A(p_input[3903]), .B(p_input[33903]), .Z(n13549) );
  AND U20326 ( .A(n13551), .B(n13552), .Z(o[3902]) );
  AND U20327 ( .A(p_input[23902]), .B(p_input[13902]), .Z(n13552) );
  AND U20328 ( .A(p_input[3902]), .B(p_input[33902]), .Z(n13551) );
  AND U20329 ( .A(n13553), .B(n13554), .Z(o[3901]) );
  AND U20330 ( .A(p_input[23901]), .B(p_input[13901]), .Z(n13554) );
  AND U20331 ( .A(p_input[3901]), .B(p_input[33901]), .Z(n13553) );
  AND U20332 ( .A(n13555), .B(n13556), .Z(o[3900]) );
  AND U20333 ( .A(p_input[23900]), .B(p_input[13900]), .Z(n13556) );
  AND U20334 ( .A(p_input[3900]), .B(p_input[33900]), .Z(n13555) );
  AND U20335 ( .A(n13557), .B(n13558), .Z(o[38]) );
  AND U20336 ( .A(p_input[20038]), .B(p_input[10038]), .Z(n13558) );
  AND U20337 ( .A(p_input[38]), .B(p_input[30038]), .Z(n13557) );
  AND U20338 ( .A(n13559), .B(n13560), .Z(o[389]) );
  AND U20339 ( .A(p_input[20389]), .B(p_input[10389]), .Z(n13560) );
  AND U20340 ( .A(p_input[389]), .B(p_input[30389]), .Z(n13559) );
  AND U20341 ( .A(n13561), .B(n13562), .Z(o[3899]) );
  AND U20342 ( .A(p_input[23899]), .B(p_input[13899]), .Z(n13562) );
  AND U20343 ( .A(p_input[3899]), .B(p_input[33899]), .Z(n13561) );
  AND U20344 ( .A(n13563), .B(n13564), .Z(o[3898]) );
  AND U20345 ( .A(p_input[23898]), .B(p_input[13898]), .Z(n13564) );
  AND U20346 ( .A(p_input[3898]), .B(p_input[33898]), .Z(n13563) );
  AND U20347 ( .A(n13565), .B(n13566), .Z(o[3897]) );
  AND U20348 ( .A(p_input[23897]), .B(p_input[13897]), .Z(n13566) );
  AND U20349 ( .A(p_input[3897]), .B(p_input[33897]), .Z(n13565) );
  AND U20350 ( .A(n13567), .B(n13568), .Z(o[3896]) );
  AND U20351 ( .A(p_input[23896]), .B(p_input[13896]), .Z(n13568) );
  AND U20352 ( .A(p_input[3896]), .B(p_input[33896]), .Z(n13567) );
  AND U20353 ( .A(n13569), .B(n13570), .Z(o[3895]) );
  AND U20354 ( .A(p_input[23895]), .B(p_input[13895]), .Z(n13570) );
  AND U20355 ( .A(p_input[3895]), .B(p_input[33895]), .Z(n13569) );
  AND U20356 ( .A(n13571), .B(n13572), .Z(o[3894]) );
  AND U20357 ( .A(p_input[23894]), .B(p_input[13894]), .Z(n13572) );
  AND U20358 ( .A(p_input[3894]), .B(p_input[33894]), .Z(n13571) );
  AND U20359 ( .A(n13573), .B(n13574), .Z(o[3893]) );
  AND U20360 ( .A(p_input[23893]), .B(p_input[13893]), .Z(n13574) );
  AND U20361 ( .A(p_input[3893]), .B(p_input[33893]), .Z(n13573) );
  AND U20362 ( .A(n13575), .B(n13576), .Z(o[3892]) );
  AND U20363 ( .A(p_input[23892]), .B(p_input[13892]), .Z(n13576) );
  AND U20364 ( .A(p_input[3892]), .B(p_input[33892]), .Z(n13575) );
  AND U20365 ( .A(n13577), .B(n13578), .Z(o[3891]) );
  AND U20366 ( .A(p_input[23891]), .B(p_input[13891]), .Z(n13578) );
  AND U20367 ( .A(p_input[3891]), .B(p_input[33891]), .Z(n13577) );
  AND U20368 ( .A(n13579), .B(n13580), .Z(o[3890]) );
  AND U20369 ( .A(p_input[23890]), .B(p_input[13890]), .Z(n13580) );
  AND U20370 ( .A(p_input[3890]), .B(p_input[33890]), .Z(n13579) );
  AND U20371 ( .A(n13581), .B(n13582), .Z(o[388]) );
  AND U20372 ( .A(p_input[20388]), .B(p_input[10388]), .Z(n13582) );
  AND U20373 ( .A(p_input[388]), .B(p_input[30388]), .Z(n13581) );
  AND U20374 ( .A(n13583), .B(n13584), .Z(o[3889]) );
  AND U20375 ( .A(p_input[23889]), .B(p_input[13889]), .Z(n13584) );
  AND U20376 ( .A(p_input[3889]), .B(p_input[33889]), .Z(n13583) );
  AND U20377 ( .A(n13585), .B(n13586), .Z(o[3888]) );
  AND U20378 ( .A(p_input[23888]), .B(p_input[13888]), .Z(n13586) );
  AND U20379 ( .A(p_input[3888]), .B(p_input[33888]), .Z(n13585) );
  AND U20380 ( .A(n13587), .B(n13588), .Z(o[3887]) );
  AND U20381 ( .A(p_input[23887]), .B(p_input[13887]), .Z(n13588) );
  AND U20382 ( .A(p_input[3887]), .B(p_input[33887]), .Z(n13587) );
  AND U20383 ( .A(n13589), .B(n13590), .Z(o[3886]) );
  AND U20384 ( .A(p_input[23886]), .B(p_input[13886]), .Z(n13590) );
  AND U20385 ( .A(p_input[3886]), .B(p_input[33886]), .Z(n13589) );
  AND U20386 ( .A(n13591), .B(n13592), .Z(o[3885]) );
  AND U20387 ( .A(p_input[23885]), .B(p_input[13885]), .Z(n13592) );
  AND U20388 ( .A(p_input[3885]), .B(p_input[33885]), .Z(n13591) );
  AND U20389 ( .A(n13593), .B(n13594), .Z(o[3884]) );
  AND U20390 ( .A(p_input[23884]), .B(p_input[13884]), .Z(n13594) );
  AND U20391 ( .A(p_input[3884]), .B(p_input[33884]), .Z(n13593) );
  AND U20392 ( .A(n13595), .B(n13596), .Z(o[3883]) );
  AND U20393 ( .A(p_input[23883]), .B(p_input[13883]), .Z(n13596) );
  AND U20394 ( .A(p_input[3883]), .B(p_input[33883]), .Z(n13595) );
  AND U20395 ( .A(n13597), .B(n13598), .Z(o[3882]) );
  AND U20396 ( .A(p_input[23882]), .B(p_input[13882]), .Z(n13598) );
  AND U20397 ( .A(p_input[3882]), .B(p_input[33882]), .Z(n13597) );
  AND U20398 ( .A(n13599), .B(n13600), .Z(o[3881]) );
  AND U20399 ( .A(p_input[23881]), .B(p_input[13881]), .Z(n13600) );
  AND U20400 ( .A(p_input[3881]), .B(p_input[33881]), .Z(n13599) );
  AND U20401 ( .A(n13601), .B(n13602), .Z(o[3880]) );
  AND U20402 ( .A(p_input[23880]), .B(p_input[13880]), .Z(n13602) );
  AND U20403 ( .A(p_input[3880]), .B(p_input[33880]), .Z(n13601) );
  AND U20404 ( .A(n13603), .B(n13604), .Z(o[387]) );
  AND U20405 ( .A(p_input[20387]), .B(p_input[10387]), .Z(n13604) );
  AND U20406 ( .A(p_input[387]), .B(p_input[30387]), .Z(n13603) );
  AND U20407 ( .A(n13605), .B(n13606), .Z(o[3879]) );
  AND U20408 ( .A(p_input[23879]), .B(p_input[13879]), .Z(n13606) );
  AND U20409 ( .A(p_input[3879]), .B(p_input[33879]), .Z(n13605) );
  AND U20410 ( .A(n13607), .B(n13608), .Z(o[3878]) );
  AND U20411 ( .A(p_input[23878]), .B(p_input[13878]), .Z(n13608) );
  AND U20412 ( .A(p_input[3878]), .B(p_input[33878]), .Z(n13607) );
  AND U20413 ( .A(n13609), .B(n13610), .Z(o[3877]) );
  AND U20414 ( .A(p_input[23877]), .B(p_input[13877]), .Z(n13610) );
  AND U20415 ( .A(p_input[3877]), .B(p_input[33877]), .Z(n13609) );
  AND U20416 ( .A(n13611), .B(n13612), .Z(o[3876]) );
  AND U20417 ( .A(p_input[23876]), .B(p_input[13876]), .Z(n13612) );
  AND U20418 ( .A(p_input[3876]), .B(p_input[33876]), .Z(n13611) );
  AND U20419 ( .A(n13613), .B(n13614), .Z(o[3875]) );
  AND U20420 ( .A(p_input[23875]), .B(p_input[13875]), .Z(n13614) );
  AND U20421 ( .A(p_input[3875]), .B(p_input[33875]), .Z(n13613) );
  AND U20422 ( .A(n13615), .B(n13616), .Z(o[3874]) );
  AND U20423 ( .A(p_input[23874]), .B(p_input[13874]), .Z(n13616) );
  AND U20424 ( .A(p_input[3874]), .B(p_input[33874]), .Z(n13615) );
  AND U20425 ( .A(n13617), .B(n13618), .Z(o[3873]) );
  AND U20426 ( .A(p_input[23873]), .B(p_input[13873]), .Z(n13618) );
  AND U20427 ( .A(p_input[3873]), .B(p_input[33873]), .Z(n13617) );
  AND U20428 ( .A(n13619), .B(n13620), .Z(o[3872]) );
  AND U20429 ( .A(p_input[23872]), .B(p_input[13872]), .Z(n13620) );
  AND U20430 ( .A(p_input[3872]), .B(p_input[33872]), .Z(n13619) );
  AND U20431 ( .A(n13621), .B(n13622), .Z(o[3871]) );
  AND U20432 ( .A(p_input[23871]), .B(p_input[13871]), .Z(n13622) );
  AND U20433 ( .A(p_input[3871]), .B(p_input[33871]), .Z(n13621) );
  AND U20434 ( .A(n13623), .B(n13624), .Z(o[3870]) );
  AND U20435 ( .A(p_input[23870]), .B(p_input[13870]), .Z(n13624) );
  AND U20436 ( .A(p_input[3870]), .B(p_input[33870]), .Z(n13623) );
  AND U20437 ( .A(n13625), .B(n13626), .Z(o[386]) );
  AND U20438 ( .A(p_input[20386]), .B(p_input[10386]), .Z(n13626) );
  AND U20439 ( .A(p_input[386]), .B(p_input[30386]), .Z(n13625) );
  AND U20440 ( .A(n13627), .B(n13628), .Z(o[3869]) );
  AND U20441 ( .A(p_input[23869]), .B(p_input[13869]), .Z(n13628) );
  AND U20442 ( .A(p_input[3869]), .B(p_input[33869]), .Z(n13627) );
  AND U20443 ( .A(n13629), .B(n13630), .Z(o[3868]) );
  AND U20444 ( .A(p_input[23868]), .B(p_input[13868]), .Z(n13630) );
  AND U20445 ( .A(p_input[3868]), .B(p_input[33868]), .Z(n13629) );
  AND U20446 ( .A(n13631), .B(n13632), .Z(o[3867]) );
  AND U20447 ( .A(p_input[23867]), .B(p_input[13867]), .Z(n13632) );
  AND U20448 ( .A(p_input[3867]), .B(p_input[33867]), .Z(n13631) );
  AND U20449 ( .A(n13633), .B(n13634), .Z(o[3866]) );
  AND U20450 ( .A(p_input[23866]), .B(p_input[13866]), .Z(n13634) );
  AND U20451 ( .A(p_input[3866]), .B(p_input[33866]), .Z(n13633) );
  AND U20452 ( .A(n13635), .B(n13636), .Z(o[3865]) );
  AND U20453 ( .A(p_input[23865]), .B(p_input[13865]), .Z(n13636) );
  AND U20454 ( .A(p_input[3865]), .B(p_input[33865]), .Z(n13635) );
  AND U20455 ( .A(n13637), .B(n13638), .Z(o[3864]) );
  AND U20456 ( .A(p_input[23864]), .B(p_input[13864]), .Z(n13638) );
  AND U20457 ( .A(p_input[3864]), .B(p_input[33864]), .Z(n13637) );
  AND U20458 ( .A(n13639), .B(n13640), .Z(o[3863]) );
  AND U20459 ( .A(p_input[23863]), .B(p_input[13863]), .Z(n13640) );
  AND U20460 ( .A(p_input[3863]), .B(p_input[33863]), .Z(n13639) );
  AND U20461 ( .A(n13641), .B(n13642), .Z(o[3862]) );
  AND U20462 ( .A(p_input[23862]), .B(p_input[13862]), .Z(n13642) );
  AND U20463 ( .A(p_input[3862]), .B(p_input[33862]), .Z(n13641) );
  AND U20464 ( .A(n13643), .B(n13644), .Z(o[3861]) );
  AND U20465 ( .A(p_input[23861]), .B(p_input[13861]), .Z(n13644) );
  AND U20466 ( .A(p_input[3861]), .B(p_input[33861]), .Z(n13643) );
  AND U20467 ( .A(n13645), .B(n13646), .Z(o[3860]) );
  AND U20468 ( .A(p_input[23860]), .B(p_input[13860]), .Z(n13646) );
  AND U20469 ( .A(p_input[3860]), .B(p_input[33860]), .Z(n13645) );
  AND U20470 ( .A(n13647), .B(n13648), .Z(o[385]) );
  AND U20471 ( .A(p_input[20385]), .B(p_input[10385]), .Z(n13648) );
  AND U20472 ( .A(p_input[385]), .B(p_input[30385]), .Z(n13647) );
  AND U20473 ( .A(n13649), .B(n13650), .Z(o[3859]) );
  AND U20474 ( .A(p_input[23859]), .B(p_input[13859]), .Z(n13650) );
  AND U20475 ( .A(p_input[3859]), .B(p_input[33859]), .Z(n13649) );
  AND U20476 ( .A(n13651), .B(n13652), .Z(o[3858]) );
  AND U20477 ( .A(p_input[23858]), .B(p_input[13858]), .Z(n13652) );
  AND U20478 ( .A(p_input[3858]), .B(p_input[33858]), .Z(n13651) );
  AND U20479 ( .A(n13653), .B(n13654), .Z(o[3857]) );
  AND U20480 ( .A(p_input[23857]), .B(p_input[13857]), .Z(n13654) );
  AND U20481 ( .A(p_input[3857]), .B(p_input[33857]), .Z(n13653) );
  AND U20482 ( .A(n13655), .B(n13656), .Z(o[3856]) );
  AND U20483 ( .A(p_input[23856]), .B(p_input[13856]), .Z(n13656) );
  AND U20484 ( .A(p_input[3856]), .B(p_input[33856]), .Z(n13655) );
  AND U20485 ( .A(n13657), .B(n13658), .Z(o[3855]) );
  AND U20486 ( .A(p_input[23855]), .B(p_input[13855]), .Z(n13658) );
  AND U20487 ( .A(p_input[3855]), .B(p_input[33855]), .Z(n13657) );
  AND U20488 ( .A(n13659), .B(n13660), .Z(o[3854]) );
  AND U20489 ( .A(p_input[23854]), .B(p_input[13854]), .Z(n13660) );
  AND U20490 ( .A(p_input[3854]), .B(p_input[33854]), .Z(n13659) );
  AND U20491 ( .A(n13661), .B(n13662), .Z(o[3853]) );
  AND U20492 ( .A(p_input[23853]), .B(p_input[13853]), .Z(n13662) );
  AND U20493 ( .A(p_input[3853]), .B(p_input[33853]), .Z(n13661) );
  AND U20494 ( .A(n13663), .B(n13664), .Z(o[3852]) );
  AND U20495 ( .A(p_input[23852]), .B(p_input[13852]), .Z(n13664) );
  AND U20496 ( .A(p_input[3852]), .B(p_input[33852]), .Z(n13663) );
  AND U20497 ( .A(n13665), .B(n13666), .Z(o[3851]) );
  AND U20498 ( .A(p_input[23851]), .B(p_input[13851]), .Z(n13666) );
  AND U20499 ( .A(p_input[3851]), .B(p_input[33851]), .Z(n13665) );
  AND U20500 ( .A(n13667), .B(n13668), .Z(o[3850]) );
  AND U20501 ( .A(p_input[23850]), .B(p_input[13850]), .Z(n13668) );
  AND U20502 ( .A(p_input[3850]), .B(p_input[33850]), .Z(n13667) );
  AND U20503 ( .A(n13669), .B(n13670), .Z(o[384]) );
  AND U20504 ( .A(p_input[20384]), .B(p_input[10384]), .Z(n13670) );
  AND U20505 ( .A(p_input[384]), .B(p_input[30384]), .Z(n13669) );
  AND U20506 ( .A(n13671), .B(n13672), .Z(o[3849]) );
  AND U20507 ( .A(p_input[23849]), .B(p_input[13849]), .Z(n13672) );
  AND U20508 ( .A(p_input[3849]), .B(p_input[33849]), .Z(n13671) );
  AND U20509 ( .A(n13673), .B(n13674), .Z(o[3848]) );
  AND U20510 ( .A(p_input[23848]), .B(p_input[13848]), .Z(n13674) );
  AND U20511 ( .A(p_input[3848]), .B(p_input[33848]), .Z(n13673) );
  AND U20512 ( .A(n13675), .B(n13676), .Z(o[3847]) );
  AND U20513 ( .A(p_input[23847]), .B(p_input[13847]), .Z(n13676) );
  AND U20514 ( .A(p_input[3847]), .B(p_input[33847]), .Z(n13675) );
  AND U20515 ( .A(n13677), .B(n13678), .Z(o[3846]) );
  AND U20516 ( .A(p_input[23846]), .B(p_input[13846]), .Z(n13678) );
  AND U20517 ( .A(p_input[3846]), .B(p_input[33846]), .Z(n13677) );
  AND U20518 ( .A(n13679), .B(n13680), .Z(o[3845]) );
  AND U20519 ( .A(p_input[23845]), .B(p_input[13845]), .Z(n13680) );
  AND U20520 ( .A(p_input[3845]), .B(p_input[33845]), .Z(n13679) );
  AND U20521 ( .A(n13681), .B(n13682), .Z(o[3844]) );
  AND U20522 ( .A(p_input[23844]), .B(p_input[13844]), .Z(n13682) );
  AND U20523 ( .A(p_input[3844]), .B(p_input[33844]), .Z(n13681) );
  AND U20524 ( .A(n13683), .B(n13684), .Z(o[3843]) );
  AND U20525 ( .A(p_input[23843]), .B(p_input[13843]), .Z(n13684) );
  AND U20526 ( .A(p_input[3843]), .B(p_input[33843]), .Z(n13683) );
  AND U20527 ( .A(n13685), .B(n13686), .Z(o[3842]) );
  AND U20528 ( .A(p_input[23842]), .B(p_input[13842]), .Z(n13686) );
  AND U20529 ( .A(p_input[3842]), .B(p_input[33842]), .Z(n13685) );
  AND U20530 ( .A(n13687), .B(n13688), .Z(o[3841]) );
  AND U20531 ( .A(p_input[23841]), .B(p_input[13841]), .Z(n13688) );
  AND U20532 ( .A(p_input[3841]), .B(p_input[33841]), .Z(n13687) );
  AND U20533 ( .A(n13689), .B(n13690), .Z(o[3840]) );
  AND U20534 ( .A(p_input[23840]), .B(p_input[13840]), .Z(n13690) );
  AND U20535 ( .A(p_input[3840]), .B(p_input[33840]), .Z(n13689) );
  AND U20536 ( .A(n13691), .B(n13692), .Z(o[383]) );
  AND U20537 ( .A(p_input[20383]), .B(p_input[10383]), .Z(n13692) );
  AND U20538 ( .A(p_input[383]), .B(p_input[30383]), .Z(n13691) );
  AND U20539 ( .A(n13693), .B(n13694), .Z(o[3839]) );
  AND U20540 ( .A(p_input[23839]), .B(p_input[13839]), .Z(n13694) );
  AND U20541 ( .A(p_input[3839]), .B(p_input[33839]), .Z(n13693) );
  AND U20542 ( .A(n13695), .B(n13696), .Z(o[3838]) );
  AND U20543 ( .A(p_input[23838]), .B(p_input[13838]), .Z(n13696) );
  AND U20544 ( .A(p_input[3838]), .B(p_input[33838]), .Z(n13695) );
  AND U20545 ( .A(n13697), .B(n13698), .Z(o[3837]) );
  AND U20546 ( .A(p_input[23837]), .B(p_input[13837]), .Z(n13698) );
  AND U20547 ( .A(p_input[3837]), .B(p_input[33837]), .Z(n13697) );
  AND U20548 ( .A(n13699), .B(n13700), .Z(o[3836]) );
  AND U20549 ( .A(p_input[23836]), .B(p_input[13836]), .Z(n13700) );
  AND U20550 ( .A(p_input[3836]), .B(p_input[33836]), .Z(n13699) );
  AND U20551 ( .A(n13701), .B(n13702), .Z(o[3835]) );
  AND U20552 ( .A(p_input[23835]), .B(p_input[13835]), .Z(n13702) );
  AND U20553 ( .A(p_input[3835]), .B(p_input[33835]), .Z(n13701) );
  AND U20554 ( .A(n13703), .B(n13704), .Z(o[3834]) );
  AND U20555 ( .A(p_input[23834]), .B(p_input[13834]), .Z(n13704) );
  AND U20556 ( .A(p_input[3834]), .B(p_input[33834]), .Z(n13703) );
  AND U20557 ( .A(n13705), .B(n13706), .Z(o[3833]) );
  AND U20558 ( .A(p_input[23833]), .B(p_input[13833]), .Z(n13706) );
  AND U20559 ( .A(p_input[3833]), .B(p_input[33833]), .Z(n13705) );
  AND U20560 ( .A(n13707), .B(n13708), .Z(o[3832]) );
  AND U20561 ( .A(p_input[23832]), .B(p_input[13832]), .Z(n13708) );
  AND U20562 ( .A(p_input[3832]), .B(p_input[33832]), .Z(n13707) );
  AND U20563 ( .A(n13709), .B(n13710), .Z(o[3831]) );
  AND U20564 ( .A(p_input[23831]), .B(p_input[13831]), .Z(n13710) );
  AND U20565 ( .A(p_input[3831]), .B(p_input[33831]), .Z(n13709) );
  AND U20566 ( .A(n13711), .B(n13712), .Z(o[3830]) );
  AND U20567 ( .A(p_input[23830]), .B(p_input[13830]), .Z(n13712) );
  AND U20568 ( .A(p_input[3830]), .B(p_input[33830]), .Z(n13711) );
  AND U20569 ( .A(n13713), .B(n13714), .Z(o[382]) );
  AND U20570 ( .A(p_input[20382]), .B(p_input[10382]), .Z(n13714) );
  AND U20571 ( .A(p_input[382]), .B(p_input[30382]), .Z(n13713) );
  AND U20572 ( .A(n13715), .B(n13716), .Z(o[3829]) );
  AND U20573 ( .A(p_input[23829]), .B(p_input[13829]), .Z(n13716) );
  AND U20574 ( .A(p_input[3829]), .B(p_input[33829]), .Z(n13715) );
  AND U20575 ( .A(n13717), .B(n13718), .Z(o[3828]) );
  AND U20576 ( .A(p_input[23828]), .B(p_input[13828]), .Z(n13718) );
  AND U20577 ( .A(p_input[3828]), .B(p_input[33828]), .Z(n13717) );
  AND U20578 ( .A(n13719), .B(n13720), .Z(o[3827]) );
  AND U20579 ( .A(p_input[23827]), .B(p_input[13827]), .Z(n13720) );
  AND U20580 ( .A(p_input[3827]), .B(p_input[33827]), .Z(n13719) );
  AND U20581 ( .A(n13721), .B(n13722), .Z(o[3826]) );
  AND U20582 ( .A(p_input[23826]), .B(p_input[13826]), .Z(n13722) );
  AND U20583 ( .A(p_input[3826]), .B(p_input[33826]), .Z(n13721) );
  AND U20584 ( .A(n13723), .B(n13724), .Z(o[3825]) );
  AND U20585 ( .A(p_input[23825]), .B(p_input[13825]), .Z(n13724) );
  AND U20586 ( .A(p_input[3825]), .B(p_input[33825]), .Z(n13723) );
  AND U20587 ( .A(n13725), .B(n13726), .Z(o[3824]) );
  AND U20588 ( .A(p_input[23824]), .B(p_input[13824]), .Z(n13726) );
  AND U20589 ( .A(p_input[3824]), .B(p_input[33824]), .Z(n13725) );
  AND U20590 ( .A(n13727), .B(n13728), .Z(o[3823]) );
  AND U20591 ( .A(p_input[23823]), .B(p_input[13823]), .Z(n13728) );
  AND U20592 ( .A(p_input[3823]), .B(p_input[33823]), .Z(n13727) );
  AND U20593 ( .A(n13729), .B(n13730), .Z(o[3822]) );
  AND U20594 ( .A(p_input[23822]), .B(p_input[13822]), .Z(n13730) );
  AND U20595 ( .A(p_input[3822]), .B(p_input[33822]), .Z(n13729) );
  AND U20596 ( .A(n13731), .B(n13732), .Z(o[3821]) );
  AND U20597 ( .A(p_input[23821]), .B(p_input[13821]), .Z(n13732) );
  AND U20598 ( .A(p_input[3821]), .B(p_input[33821]), .Z(n13731) );
  AND U20599 ( .A(n13733), .B(n13734), .Z(o[3820]) );
  AND U20600 ( .A(p_input[23820]), .B(p_input[13820]), .Z(n13734) );
  AND U20601 ( .A(p_input[3820]), .B(p_input[33820]), .Z(n13733) );
  AND U20602 ( .A(n13735), .B(n13736), .Z(o[381]) );
  AND U20603 ( .A(p_input[20381]), .B(p_input[10381]), .Z(n13736) );
  AND U20604 ( .A(p_input[381]), .B(p_input[30381]), .Z(n13735) );
  AND U20605 ( .A(n13737), .B(n13738), .Z(o[3819]) );
  AND U20606 ( .A(p_input[23819]), .B(p_input[13819]), .Z(n13738) );
  AND U20607 ( .A(p_input[3819]), .B(p_input[33819]), .Z(n13737) );
  AND U20608 ( .A(n13739), .B(n13740), .Z(o[3818]) );
  AND U20609 ( .A(p_input[23818]), .B(p_input[13818]), .Z(n13740) );
  AND U20610 ( .A(p_input[3818]), .B(p_input[33818]), .Z(n13739) );
  AND U20611 ( .A(n13741), .B(n13742), .Z(o[3817]) );
  AND U20612 ( .A(p_input[23817]), .B(p_input[13817]), .Z(n13742) );
  AND U20613 ( .A(p_input[3817]), .B(p_input[33817]), .Z(n13741) );
  AND U20614 ( .A(n13743), .B(n13744), .Z(o[3816]) );
  AND U20615 ( .A(p_input[23816]), .B(p_input[13816]), .Z(n13744) );
  AND U20616 ( .A(p_input[3816]), .B(p_input[33816]), .Z(n13743) );
  AND U20617 ( .A(n13745), .B(n13746), .Z(o[3815]) );
  AND U20618 ( .A(p_input[23815]), .B(p_input[13815]), .Z(n13746) );
  AND U20619 ( .A(p_input[3815]), .B(p_input[33815]), .Z(n13745) );
  AND U20620 ( .A(n13747), .B(n13748), .Z(o[3814]) );
  AND U20621 ( .A(p_input[23814]), .B(p_input[13814]), .Z(n13748) );
  AND U20622 ( .A(p_input[3814]), .B(p_input[33814]), .Z(n13747) );
  AND U20623 ( .A(n13749), .B(n13750), .Z(o[3813]) );
  AND U20624 ( .A(p_input[23813]), .B(p_input[13813]), .Z(n13750) );
  AND U20625 ( .A(p_input[3813]), .B(p_input[33813]), .Z(n13749) );
  AND U20626 ( .A(n13751), .B(n13752), .Z(o[3812]) );
  AND U20627 ( .A(p_input[23812]), .B(p_input[13812]), .Z(n13752) );
  AND U20628 ( .A(p_input[3812]), .B(p_input[33812]), .Z(n13751) );
  AND U20629 ( .A(n13753), .B(n13754), .Z(o[3811]) );
  AND U20630 ( .A(p_input[23811]), .B(p_input[13811]), .Z(n13754) );
  AND U20631 ( .A(p_input[3811]), .B(p_input[33811]), .Z(n13753) );
  AND U20632 ( .A(n13755), .B(n13756), .Z(o[3810]) );
  AND U20633 ( .A(p_input[23810]), .B(p_input[13810]), .Z(n13756) );
  AND U20634 ( .A(p_input[3810]), .B(p_input[33810]), .Z(n13755) );
  AND U20635 ( .A(n13757), .B(n13758), .Z(o[380]) );
  AND U20636 ( .A(p_input[20380]), .B(p_input[10380]), .Z(n13758) );
  AND U20637 ( .A(p_input[380]), .B(p_input[30380]), .Z(n13757) );
  AND U20638 ( .A(n13759), .B(n13760), .Z(o[3809]) );
  AND U20639 ( .A(p_input[23809]), .B(p_input[13809]), .Z(n13760) );
  AND U20640 ( .A(p_input[3809]), .B(p_input[33809]), .Z(n13759) );
  AND U20641 ( .A(n13761), .B(n13762), .Z(o[3808]) );
  AND U20642 ( .A(p_input[23808]), .B(p_input[13808]), .Z(n13762) );
  AND U20643 ( .A(p_input[3808]), .B(p_input[33808]), .Z(n13761) );
  AND U20644 ( .A(n13763), .B(n13764), .Z(o[3807]) );
  AND U20645 ( .A(p_input[23807]), .B(p_input[13807]), .Z(n13764) );
  AND U20646 ( .A(p_input[3807]), .B(p_input[33807]), .Z(n13763) );
  AND U20647 ( .A(n13765), .B(n13766), .Z(o[3806]) );
  AND U20648 ( .A(p_input[23806]), .B(p_input[13806]), .Z(n13766) );
  AND U20649 ( .A(p_input[3806]), .B(p_input[33806]), .Z(n13765) );
  AND U20650 ( .A(n13767), .B(n13768), .Z(o[3805]) );
  AND U20651 ( .A(p_input[23805]), .B(p_input[13805]), .Z(n13768) );
  AND U20652 ( .A(p_input[3805]), .B(p_input[33805]), .Z(n13767) );
  AND U20653 ( .A(n13769), .B(n13770), .Z(o[3804]) );
  AND U20654 ( .A(p_input[23804]), .B(p_input[13804]), .Z(n13770) );
  AND U20655 ( .A(p_input[3804]), .B(p_input[33804]), .Z(n13769) );
  AND U20656 ( .A(n13771), .B(n13772), .Z(o[3803]) );
  AND U20657 ( .A(p_input[23803]), .B(p_input[13803]), .Z(n13772) );
  AND U20658 ( .A(p_input[3803]), .B(p_input[33803]), .Z(n13771) );
  AND U20659 ( .A(n13773), .B(n13774), .Z(o[3802]) );
  AND U20660 ( .A(p_input[23802]), .B(p_input[13802]), .Z(n13774) );
  AND U20661 ( .A(p_input[3802]), .B(p_input[33802]), .Z(n13773) );
  AND U20662 ( .A(n13775), .B(n13776), .Z(o[3801]) );
  AND U20663 ( .A(p_input[23801]), .B(p_input[13801]), .Z(n13776) );
  AND U20664 ( .A(p_input[3801]), .B(p_input[33801]), .Z(n13775) );
  AND U20665 ( .A(n13777), .B(n13778), .Z(o[3800]) );
  AND U20666 ( .A(p_input[23800]), .B(p_input[13800]), .Z(n13778) );
  AND U20667 ( .A(p_input[3800]), .B(p_input[33800]), .Z(n13777) );
  AND U20668 ( .A(n13779), .B(n13780), .Z(o[37]) );
  AND U20669 ( .A(p_input[20037]), .B(p_input[10037]), .Z(n13780) );
  AND U20670 ( .A(p_input[37]), .B(p_input[30037]), .Z(n13779) );
  AND U20671 ( .A(n13781), .B(n13782), .Z(o[379]) );
  AND U20672 ( .A(p_input[20379]), .B(p_input[10379]), .Z(n13782) );
  AND U20673 ( .A(p_input[379]), .B(p_input[30379]), .Z(n13781) );
  AND U20674 ( .A(n13783), .B(n13784), .Z(o[3799]) );
  AND U20675 ( .A(p_input[23799]), .B(p_input[13799]), .Z(n13784) );
  AND U20676 ( .A(p_input[3799]), .B(p_input[33799]), .Z(n13783) );
  AND U20677 ( .A(n13785), .B(n13786), .Z(o[3798]) );
  AND U20678 ( .A(p_input[23798]), .B(p_input[13798]), .Z(n13786) );
  AND U20679 ( .A(p_input[3798]), .B(p_input[33798]), .Z(n13785) );
  AND U20680 ( .A(n13787), .B(n13788), .Z(o[3797]) );
  AND U20681 ( .A(p_input[23797]), .B(p_input[13797]), .Z(n13788) );
  AND U20682 ( .A(p_input[3797]), .B(p_input[33797]), .Z(n13787) );
  AND U20683 ( .A(n13789), .B(n13790), .Z(o[3796]) );
  AND U20684 ( .A(p_input[23796]), .B(p_input[13796]), .Z(n13790) );
  AND U20685 ( .A(p_input[3796]), .B(p_input[33796]), .Z(n13789) );
  AND U20686 ( .A(n13791), .B(n13792), .Z(o[3795]) );
  AND U20687 ( .A(p_input[23795]), .B(p_input[13795]), .Z(n13792) );
  AND U20688 ( .A(p_input[3795]), .B(p_input[33795]), .Z(n13791) );
  AND U20689 ( .A(n13793), .B(n13794), .Z(o[3794]) );
  AND U20690 ( .A(p_input[23794]), .B(p_input[13794]), .Z(n13794) );
  AND U20691 ( .A(p_input[3794]), .B(p_input[33794]), .Z(n13793) );
  AND U20692 ( .A(n13795), .B(n13796), .Z(o[3793]) );
  AND U20693 ( .A(p_input[23793]), .B(p_input[13793]), .Z(n13796) );
  AND U20694 ( .A(p_input[3793]), .B(p_input[33793]), .Z(n13795) );
  AND U20695 ( .A(n13797), .B(n13798), .Z(o[3792]) );
  AND U20696 ( .A(p_input[23792]), .B(p_input[13792]), .Z(n13798) );
  AND U20697 ( .A(p_input[3792]), .B(p_input[33792]), .Z(n13797) );
  AND U20698 ( .A(n13799), .B(n13800), .Z(o[3791]) );
  AND U20699 ( .A(p_input[23791]), .B(p_input[13791]), .Z(n13800) );
  AND U20700 ( .A(p_input[3791]), .B(p_input[33791]), .Z(n13799) );
  AND U20701 ( .A(n13801), .B(n13802), .Z(o[3790]) );
  AND U20702 ( .A(p_input[23790]), .B(p_input[13790]), .Z(n13802) );
  AND U20703 ( .A(p_input[3790]), .B(p_input[33790]), .Z(n13801) );
  AND U20704 ( .A(n13803), .B(n13804), .Z(o[378]) );
  AND U20705 ( .A(p_input[20378]), .B(p_input[10378]), .Z(n13804) );
  AND U20706 ( .A(p_input[378]), .B(p_input[30378]), .Z(n13803) );
  AND U20707 ( .A(n13805), .B(n13806), .Z(o[3789]) );
  AND U20708 ( .A(p_input[23789]), .B(p_input[13789]), .Z(n13806) );
  AND U20709 ( .A(p_input[3789]), .B(p_input[33789]), .Z(n13805) );
  AND U20710 ( .A(n13807), .B(n13808), .Z(o[3788]) );
  AND U20711 ( .A(p_input[23788]), .B(p_input[13788]), .Z(n13808) );
  AND U20712 ( .A(p_input[3788]), .B(p_input[33788]), .Z(n13807) );
  AND U20713 ( .A(n13809), .B(n13810), .Z(o[3787]) );
  AND U20714 ( .A(p_input[23787]), .B(p_input[13787]), .Z(n13810) );
  AND U20715 ( .A(p_input[3787]), .B(p_input[33787]), .Z(n13809) );
  AND U20716 ( .A(n13811), .B(n13812), .Z(o[3786]) );
  AND U20717 ( .A(p_input[23786]), .B(p_input[13786]), .Z(n13812) );
  AND U20718 ( .A(p_input[3786]), .B(p_input[33786]), .Z(n13811) );
  AND U20719 ( .A(n13813), .B(n13814), .Z(o[3785]) );
  AND U20720 ( .A(p_input[23785]), .B(p_input[13785]), .Z(n13814) );
  AND U20721 ( .A(p_input[3785]), .B(p_input[33785]), .Z(n13813) );
  AND U20722 ( .A(n13815), .B(n13816), .Z(o[3784]) );
  AND U20723 ( .A(p_input[23784]), .B(p_input[13784]), .Z(n13816) );
  AND U20724 ( .A(p_input[3784]), .B(p_input[33784]), .Z(n13815) );
  AND U20725 ( .A(n13817), .B(n13818), .Z(o[3783]) );
  AND U20726 ( .A(p_input[23783]), .B(p_input[13783]), .Z(n13818) );
  AND U20727 ( .A(p_input[3783]), .B(p_input[33783]), .Z(n13817) );
  AND U20728 ( .A(n13819), .B(n13820), .Z(o[3782]) );
  AND U20729 ( .A(p_input[23782]), .B(p_input[13782]), .Z(n13820) );
  AND U20730 ( .A(p_input[3782]), .B(p_input[33782]), .Z(n13819) );
  AND U20731 ( .A(n13821), .B(n13822), .Z(o[3781]) );
  AND U20732 ( .A(p_input[23781]), .B(p_input[13781]), .Z(n13822) );
  AND U20733 ( .A(p_input[3781]), .B(p_input[33781]), .Z(n13821) );
  AND U20734 ( .A(n13823), .B(n13824), .Z(o[3780]) );
  AND U20735 ( .A(p_input[23780]), .B(p_input[13780]), .Z(n13824) );
  AND U20736 ( .A(p_input[3780]), .B(p_input[33780]), .Z(n13823) );
  AND U20737 ( .A(n13825), .B(n13826), .Z(o[377]) );
  AND U20738 ( .A(p_input[20377]), .B(p_input[10377]), .Z(n13826) );
  AND U20739 ( .A(p_input[377]), .B(p_input[30377]), .Z(n13825) );
  AND U20740 ( .A(n13827), .B(n13828), .Z(o[3779]) );
  AND U20741 ( .A(p_input[23779]), .B(p_input[13779]), .Z(n13828) );
  AND U20742 ( .A(p_input[3779]), .B(p_input[33779]), .Z(n13827) );
  AND U20743 ( .A(n13829), .B(n13830), .Z(o[3778]) );
  AND U20744 ( .A(p_input[23778]), .B(p_input[13778]), .Z(n13830) );
  AND U20745 ( .A(p_input[3778]), .B(p_input[33778]), .Z(n13829) );
  AND U20746 ( .A(n13831), .B(n13832), .Z(o[3777]) );
  AND U20747 ( .A(p_input[23777]), .B(p_input[13777]), .Z(n13832) );
  AND U20748 ( .A(p_input[3777]), .B(p_input[33777]), .Z(n13831) );
  AND U20749 ( .A(n13833), .B(n13834), .Z(o[3776]) );
  AND U20750 ( .A(p_input[23776]), .B(p_input[13776]), .Z(n13834) );
  AND U20751 ( .A(p_input[3776]), .B(p_input[33776]), .Z(n13833) );
  AND U20752 ( .A(n13835), .B(n13836), .Z(o[3775]) );
  AND U20753 ( .A(p_input[23775]), .B(p_input[13775]), .Z(n13836) );
  AND U20754 ( .A(p_input[3775]), .B(p_input[33775]), .Z(n13835) );
  AND U20755 ( .A(n13837), .B(n13838), .Z(o[3774]) );
  AND U20756 ( .A(p_input[23774]), .B(p_input[13774]), .Z(n13838) );
  AND U20757 ( .A(p_input[3774]), .B(p_input[33774]), .Z(n13837) );
  AND U20758 ( .A(n13839), .B(n13840), .Z(o[3773]) );
  AND U20759 ( .A(p_input[23773]), .B(p_input[13773]), .Z(n13840) );
  AND U20760 ( .A(p_input[3773]), .B(p_input[33773]), .Z(n13839) );
  AND U20761 ( .A(n13841), .B(n13842), .Z(o[3772]) );
  AND U20762 ( .A(p_input[23772]), .B(p_input[13772]), .Z(n13842) );
  AND U20763 ( .A(p_input[3772]), .B(p_input[33772]), .Z(n13841) );
  AND U20764 ( .A(n13843), .B(n13844), .Z(o[3771]) );
  AND U20765 ( .A(p_input[23771]), .B(p_input[13771]), .Z(n13844) );
  AND U20766 ( .A(p_input[3771]), .B(p_input[33771]), .Z(n13843) );
  AND U20767 ( .A(n13845), .B(n13846), .Z(o[3770]) );
  AND U20768 ( .A(p_input[23770]), .B(p_input[13770]), .Z(n13846) );
  AND U20769 ( .A(p_input[3770]), .B(p_input[33770]), .Z(n13845) );
  AND U20770 ( .A(n13847), .B(n13848), .Z(o[376]) );
  AND U20771 ( .A(p_input[20376]), .B(p_input[10376]), .Z(n13848) );
  AND U20772 ( .A(p_input[376]), .B(p_input[30376]), .Z(n13847) );
  AND U20773 ( .A(n13849), .B(n13850), .Z(o[3769]) );
  AND U20774 ( .A(p_input[23769]), .B(p_input[13769]), .Z(n13850) );
  AND U20775 ( .A(p_input[3769]), .B(p_input[33769]), .Z(n13849) );
  AND U20776 ( .A(n13851), .B(n13852), .Z(o[3768]) );
  AND U20777 ( .A(p_input[23768]), .B(p_input[13768]), .Z(n13852) );
  AND U20778 ( .A(p_input[3768]), .B(p_input[33768]), .Z(n13851) );
  AND U20779 ( .A(n13853), .B(n13854), .Z(o[3767]) );
  AND U20780 ( .A(p_input[23767]), .B(p_input[13767]), .Z(n13854) );
  AND U20781 ( .A(p_input[3767]), .B(p_input[33767]), .Z(n13853) );
  AND U20782 ( .A(n13855), .B(n13856), .Z(o[3766]) );
  AND U20783 ( .A(p_input[23766]), .B(p_input[13766]), .Z(n13856) );
  AND U20784 ( .A(p_input[3766]), .B(p_input[33766]), .Z(n13855) );
  AND U20785 ( .A(n13857), .B(n13858), .Z(o[3765]) );
  AND U20786 ( .A(p_input[23765]), .B(p_input[13765]), .Z(n13858) );
  AND U20787 ( .A(p_input[3765]), .B(p_input[33765]), .Z(n13857) );
  AND U20788 ( .A(n13859), .B(n13860), .Z(o[3764]) );
  AND U20789 ( .A(p_input[23764]), .B(p_input[13764]), .Z(n13860) );
  AND U20790 ( .A(p_input[3764]), .B(p_input[33764]), .Z(n13859) );
  AND U20791 ( .A(n13861), .B(n13862), .Z(o[3763]) );
  AND U20792 ( .A(p_input[23763]), .B(p_input[13763]), .Z(n13862) );
  AND U20793 ( .A(p_input[3763]), .B(p_input[33763]), .Z(n13861) );
  AND U20794 ( .A(n13863), .B(n13864), .Z(o[3762]) );
  AND U20795 ( .A(p_input[23762]), .B(p_input[13762]), .Z(n13864) );
  AND U20796 ( .A(p_input[3762]), .B(p_input[33762]), .Z(n13863) );
  AND U20797 ( .A(n13865), .B(n13866), .Z(o[3761]) );
  AND U20798 ( .A(p_input[23761]), .B(p_input[13761]), .Z(n13866) );
  AND U20799 ( .A(p_input[3761]), .B(p_input[33761]), .Z(n13865) );
  AND U20800 ( .A(n13867), .B(n13868), .Z(o[3760]) );
  AND U20801 ( .A(p_input[23760]), .B(p_input[13760]), .Z(n13868) );
  AND U20802 ( .A(p_input[3760]), .B(p_input[33760]), .Z(n13867) );
  AND U20803 ( .A(n13869), .B(n13870), .Z(o[375]) );
  AND U20804 ( .A(p_input[20375]), .B(p_input[10375]), .Z(n13870) );
  AND U20805 ( .A(p_input[375]), .B(p_input[30375]), .Z(n13869) );
  AND U20806 ( .A(n13871), .B(n13872), .Z(o[3759]) );
  AND U20807 ( .A(p_input[23759]), .B(p_input[13759]), .Z(n13872) );
  AND U20808 ( .A(p_input[3759]), .B(p_input[33759]), .Z(n13871) );
  AND U20809 ( .A(n13873), .B(n13874), .Z(o[3758]) );
  AND U20810 ( .A(p_input[23758]), .B(p_input[13758]), .Z(n13874) );
  AND U20811 ( .A(p_input[3758]), .B(p_input[33758]), .Z(n13873) );
  AND U20812 ( .A(n13875), .B(n13876), .Z(o[3757]) );
  AND U20813 ( .A(p_input[23757]), .B(p_input[13757]), .Z(n13876) );
  AND U20814 ( .A(p_input[3757]), .B(p_input[33757]), .Z(n13875) );
  AND U20815 ( .A(n13877), .B(n13878), .Z(o[3756]) );
  AND U20816 ( .A(p_input[23756]), .B(p_input[13756]), .Z(n13878) );
  AND U20817 ( .A(p_input[3756]), .B(p_input[33756]), .Z(n13877) );
  AND U20818 ( .A(n13879), .B(n13880), .Z(o[3755]) );
  AND U20819 ( .A(p_input[23755]), .B(p_input[13755]), .Z(n13880) );
  AND U20820 ( .A(p_input[3755]), .B(p_input[33755]), .Z(n13879) );
  AND U20821 ( .A(n13881), .B(n13882), .Z(o[3754]) );
  AND U20822 ( .A(p_input[23754]), .B(p_input[13754]), .Z(n13882) );
  AND U20823 ( .A(p_input[3754]), .B(p_input[33754]), .Z(n13881) );
  AND U20824 ( .A(n13883), .B(n13884), .Z(o[3753]) );
  AND U20825 ( .A(p_input[23753]), .B(p_input[13753]), .Z(n13884) );
  AND U20826 ( .A(p_input[3753]), .B(p_input[33753]), .Z(n13883) );
  AND U20827 ( .A(n13885), .B(n13886), .Z(o[3752]) );
  AND U20828 ( .A(p_input[23752]), .B(p_input[13752]), .Z(n13886) );
  AND U20829 ( .A(p_input[3752]), .B(p_input[33752]), .Z(n13885) );
  AND U20830 ( .A(n13887), .B(n13888), .Z(o[3751]) );
  AND U20831 ( .A(p_input[23751]), .B(p_input[13751]), .Z(n13888) );
  AND U20832 ( .A(p_input[3751]), .B(p_input[33751]), .Z(n13887) );
  AND U20833 ( .A(n13889), .B(n13890), .Z(o[3750]) );
  AND U20834 ( .A(p_input[23750]), .B(p_input[13750]), .Z(n13890) );
  AND U20835 ( .A(p_input[3750]), .B(p_input[33750]), .Z(n13889) );
  AND U20836 ( .A(n13891), .B(n13892), .Z(o[374]) );
  AND U20837 ( .A(p_input[20374]), .B(p_input[10374]), .Z(n13892) );
  AND U20838 ( .A(p_input[374]), .B(p_input[30374]), .Z(n13891) );
  AND U20839 ( .A(n13893), .B(n13894), .Z(o[3749]) );
  AND U20840 ( .A(p_input[23749]), .B(p_input[13749]), .Z(n13894) );
  AND U20841 ( .A(p_input[3749]), .B(p_input[33749]), .Z(n13893) );
  AND U20842 ( .A(n13895), .B(n13896), .Z(o[3748]) );
  AND U20843 ( .A(p_input[23748]), .B(p_input[13748]), .Z(n13896) );
  AND U20844 ( .A(p_input[3748]), .B(p_input[33748]), .Z(n13895) );
  AND U20845 ( .A(n13897), .B(n13898), .Z(o[3747]) );
  AND U20846 ( .A(p_input[23747]), .B(p_input[13747]), .Z(n13898) );
  AND U20847 ( .A(p_input[3747]), .B(p_input[33747]), .Z(n13897) );
  AND U20848 ( .A(n13899), .B(n13900), .Z(o[3746]) );
  AND U20849 ( .A(p_input[23746]), .B(p_input[13746]), .Z(n13900) );
  AND U20850 ( .A(p_input[3746]), .B(p_input[33746]), .Z(n13899) );
  AND U20851 ( .A(n13901), .B(n13902), .Z(o[3745]) );
  AND U20852 ( .A(p_input[23745]), .B(p_input[13745]), .Z(n13902) );
  AND U20853 ( .A(p_input[3745]), .B(p_input[33745]), .Z(n13901) );
  AND U20854 ( .A(n13903), .B(n13904), .Z(o[3744]) );
  AND U20855 ( .A(p_input[23744]), .B(p_input[13744]), .Z(n13904) );
  AND U20856 ( .A(p_input[3744]), .B(p_input[33744]), .Z(n13903) );
  AND U20857 ( .A(n13905), .B(n13906), .Z(o[3743]) );
  AND U20858 ( .A(p_input[23743]), .B(p_input[13743]), .Z(n13906) );
  AND U20859 ( .A(p_input[3743]), .B(p_input[33743]), .Z(n13905) );
  AND U20860 ( .A(n13907), .B(n13908), .Z(o[3742]) );
  AND U20861 ( .A(p_input[23742]), .B(p_input[13742]), .Z(n13908) );
  AND U20862 ( .A(p_input[3742]), .B(p_input[33742]), .Z(n13907) );
  AND U20863 ( .A(n13909), .B(n13910), .Z(o[3741]) );
  AND U20864 ( .A(p_input[23741]), .B(p_input[13741]), .Z(n13910) );
  AND U20865 ( .A(p_input[3741]), .B(p_input[33741]), .Z(n13909) );
  AND U20866 ( .A(n13911), .B(n13912), .Z(o[3740]) );
  AND U20867 ( .A(p_input[23740]), .B(p_input[13740]), .Z(n13912) );
  AND U20868 ( .A(p_input[3740]), .B(p_input[33740]), .Z(n13911) );
  AND U20869 ( .A(n13913), .B(n13914), .Z(o[373]) );
  AND U20870 ( .A(p_input[20373]), .B(p_input[10373]), .Z(n13914) );
  AND U20871 ( .A(p_input[373]), .B(p_input[30373]), .Z(n13913) );
  AND U20872 ( .A(n13915), .B(n13916), .Z(o[3739]) );
  AND U20873 ( .A(p_input[23739]), .B(p_input[13739]), .Z(n13916) );
  AND U20874 ( .A(p_input[3739]), .B(p_input[33739]), .Z(n13915) );
  AND U20875 ( .A(n13917), .B(n13918), .Z(o[3738]) );
  AND U20876 ( .A(p_input[23738]), .B(p_input[13738]), .Z(n13918) );
  AND U20877 ( .A(p_input[3738]), .B(p_input[33738]), .Z(n13917) );
  AND U20878 ( .A(n13919), .B(n13920), .Z(o[3737]) );
  AND U20879 ( .A(p_input[23737]), .B(p_input[13737]), .Z(n13920) );
  AND U20880 ( .A(p_input[3737]), .B(p_input[33737]), .Z(n13919) );
  AND U20881 ( .A(n13921), .B(n13922), .Z(o[3736]) );
  AND U20882 ( .A(p_input[23736]), .B(p_input[13736]), .Z(n13922) );
  AND U20883 ( .A(p_input[3736]), .B(p_input[33736]), .Z(n13921) );
  AND U20884 ( .A(n13923), .B(n13924), .Z(o[3735]) );
  AND U20885 ( .A(p_input[23735]), .B(p_input[13735]), .Z(n13924) );
  AND U20886 ( .A(p_input[3735]), .B(p_input[33735]), .Z(n13923) );
  AND U20887 ( .A(n13925), .B(n13926), .Z(o[3734]) );
  AND U20888 ( .A(p_input[23734]), .B(p_input[13734]), .Z(n13926) );
  AND U20889 ( .A(p_input[3734]), .B(p_input[33734]), .Z(n13925) );
  AND U20890 ( .A(n13927), .B(n13928), .Z(o[3733]) );
  AND U20891 ( .A(p_input[23733]), .B(p_input[13733]), .Z(n13928) );
  AND U20892 ( .A(p_input[3733]), .B(p_input[33733]), .Z(n13927) );
  AND U20893 ( .A(n13929), .B(n13930), .Z(o[3732]) );
  AND U20894 ( .A(p_input[23732]), .B(p_input[13732]), .Z(n13930) );
  AND U20895 ( .A(p_input[3732]), .B(p_input[33732]), .Z(n13929) );
  AND U20896 ( .A(n13931), .B(n13932), .Z(o[3731]) );
  AND U20897 ( .A(p_input[23731]), .B(p_input[13731]), .Z(n13932) );
  AND U20898 ( .A(p_input[3731]), .B(p_input[33731]), .Z(n13931) );
  AND U20899 ( .A(n13933), .B(n13934), .Z(o[3730]) );
  AND U20900 ( .A(p_input[23730]), .B(p_input[13730]), .Z(n13934) );
  AND U20901 ( .A(p_input[3730]), .B(p_input[33730]), .Z(n13933) );
  AND U20902 ( .A(n13935), .B(n13936), .Z(o[372]) );
  AND U20903 ( .A(p_input[20372]), .B(p_input[10372]), .Z(n13936) );
  AND U20904 ( .A(p_input[372]), .B(p_input[30372]), .Z(n13935) );
  AND U20905 ( .A(n13937), .B(n13938), .Z(o[3729]) );
  AND U20906 ( .A(p_input[23729]), .B(p_input[13729]), .Z(n13938) );
  AND U20907 ( .A(p_input[3729]), .B(p_input[33729]), .Z(n13937) );
  AND U20908 ( .A(n13939), .B(n13940), .Z(o[3728]) );
  AND U20909 ( .A(p_input[23728]), .B(p_input[13728]), .Z(n13940) );
  AND U20910 ( .A(p_input[3728]), .B(p_input[33728]), .Z(n13939) );
  AND U20911 ( .A(n13941), .B(n13942), .Z(o[3727]) );
  AND U20912 ( .A(p_input[23727]), .B(p_input[13727]), .Z(n13942) );
  AND U20913 ( .A(p_input[3727]), .B(p_input[33727]), .Z(n13941) );
  AND U20914 ( .A(n13943), .B(n13944), .Z(o[3726]) );
  AND U20915 ( .A(p_input[23726]), .B(p_input[13726]), .Z(n13944) );
  AND U20916 ( .A(p_input[3726]), .B(p_input[33726]), .Z(n13943) );
  AND U20917 ( .A(n13945), .B(n13946), .Z(o[3725]) );
  AND U20918 ( .A(p_input[23725]), .B(p_input[13725]), .Z(n13946) );
  AND U20919 ( .A(p_input[3725]), .B(p_input[33725]), .Z(n13945) );
  AND U20920 ( .A(n13947), .B(n13948), .Z(o[3724]) );
  AND U20921 ( .A(p_input[23724]), .B(p_input[13724]), .Z(n13948) );
  AND U20922 ( .A(p_input[3724]), .B(p_input[33724]), .Z(n13947) );
  AND U20923 ( .A(n13949), .B(n13950), .Z(o[3723]) );
  AND U20924 ( .A(p_input[23723]), .B(p_input[13723]), .Z(n13950) );
  AND U20925 ( .A(p_input[3723]), .B(p_input[33723]), .Z(n13949) );
  AND U20926 ( .A(n13951), .B(n13952), .Z(o[3722]) );
  AND U20927 ( .A(p_input[23722]), .B(p_input[13722]), .Z(n13952) );
  AND U20928 ( .A(p_input[3722]), .B(p_input[33722]), .Z(n13951) );
  AND U20929 ( .A(n13953), .B(n13954), .Z(o[3721]) );
  AND U20930 ( .A(p_input[23721]), .B(p_input[13721]), .Z(n13954) );
  AND U20931 ( .A(p_input[3721]), .B(p_input[33721]), .Z(n13953) );
  AND U20932 ( .A(n13955), .B(n13956), .Z(o[3720]) );
  AND U20933 ( .A(p_input[23720]), .B(p_input[13720]), .Z(n13956) );
  AND U20934 ( .A(p_input[3720]), .B(p_input[33720]), .Z(n13955) );
  AND U20935 ( .A(n13957), .B(n13958), .Z(o[371]) );
  AND U20936 ( .A(p_input[20371]), .B(p_input[10371]), .Z(n13958) );
  AND U20937 ( .A(p_input[371]), .B(p_input[30371]), .Z(n13957) );
  AND U20938 ( .A(n13959), .B(n13960), .Z(o[3719]) );
  AND U20939 ( .A(p_input[23719]), .B(p_input[13719]), .Z(n13960) );
  AND U20940 ( .A(p_input[3719]), .B(p_input[33719]), .Z(n13959) );
  AND U20941 ( .A(n13961), .B(n13962), .Z(o[3718]) );
  AND U20942 ( .A(p_input[23718]), .B(p_input[13718]), .Z(n13962) );
  AND U20943 ( .A(p_input[3718]), .B(p_input[33718]), .Z(n13961) );
  AND U20944 ( .A(n13963), .B(n13964), .Z(o[3717]) );
  AND U20945 ( .A(p_input[23717]), .B(p_input[13717]), .Z(n13964) );
  AND U20946 ( .A(p_input[3717]), .B(p_input[33717]), .Z(n13963) );
  AND U20947 ( .A(n13965), .B(n13966), .Z(o[3716]) );
  AND U20948 ( .A(p_input[23716]), .B(p_input[13716]), .Z(n13966) );
  AND U20949 ( .A(p_input[3716]), .B(p_input[33716]), .Z(n13965) );
  AND U20950 ( .A(n13967), .B(n13968), .Z(o[3715]) );
  AND U20951 ( .A(p_input[23715]), .B(p_input[13715]), .Z(n13968) );
  AND U20952 ( .A(p_input[3715]), .B(p_input[33715]), .Z(n13967) );
  AND U20953 ( .A(n13969), .B(n13970), .Z(o[3714]) );
  AND U20954 ( .A(p_input[23714]), .B(p_input[13714]), .Z(n13970) );
  AND U20955 ( .A(p_input[3714]), .B(p_input[33714]), .Z(n13969) );
  AND U20956 ( .A(n13971), .B(n13972), .Z(o[3713]) );
  AND U20957 ( .A(p_input[23713]), .B(p_input[13713]), .Z(n13972) );
  AND U20958 ( .A(p_input[3713]), .B(p_input[33713]), .Z(n13971) );
  AND U20959 ( .A(n13973), .B(n13974), .Z(o[3712]) );
  AND U20960 ( .A(p_input[23712]), .B(p_input[13712]), .Z(n13974) );
  AND U20961 ( .A(p_input[3712]), .B(p_input[33712]), .Z(n13973) );
  AND U20962 ( .A(n13975), .B(n13976), .Z(o[3711]) );
  AND U20963 ( .A(p_input[23711]), .B(p_input[13711]), .Z(n13976) );
  AND U20964 ( .A(p_input[3711]), .B(p_input[33711]), .Z(n13975) );
  AND U20965 ( .A(n13977), .B(n13978), .Z(o[3710]) );
  AND U20966 ( .A(p_input[23710]), .B(p_input[13710]), .Z(n13978) );
  AND U20967 ( .A(p_input[3710]), .B(p_input[33710]), .Z(n13977) );
  AND U20968 ( .A(n13979), .B(n13980), .Z(o[370]) );
  AND U20969 ( .A(p_input[20370]), .B(p_input[10370]), .Z(n13980) );
  AND U20970 ( .A(p_input[370]), .B(p_input[30370]), .Z(n13979) );
  AND U20971 ( .A(n13981), .B(n13982), .Z(o[3709]) );
  AND U20972 ( .A(p_input[23709]), .B(p_input[13709]), .Z(n13982) );
  AND U20973 ( .A(p_input[3709]), .B(p_input[33709]), .Z(n13981) );
  AND U20974 ( .A(n13983), .B(n13984), .Z(o[3708]) );
  AND U20975 ( .A(p_input[23708]), .B(p_input[13708]), .Z(n13984) );
  AND U20976 ( .A(p_input[3708]), .B(p_input[33708]), .Z(n13983) );
  AND U20977 ( .A(n13985), .B(n13986), .Z(o[3707]) );
  AND U20978 ( .A(p_input[23707]), .B(p_input[13707]), .Z(n13986) );
  AND U20979 ( .A(p_input[3707]), .B(p_input[33707]), .Z(n13985) );
  AND U20980 ( .A(n13987), .B(n13988), .Z(o[3706]) );
  AND U20981 ( .A(p_input[23706]), .B(p_input[13706]), .Z(n13988) );
  AND U20982 ( .A(p_input[3706]), .B(p_input[33706]), .Z(n13987) );
  AND U20983 ( .A(n13989), .B(n13990), .Z(o[3705]) );
  AND U20984 ( .A(p_input[23705]), .B(p_input[13705]), .Z(n13990) );
  AND U20985 ( .A(p_input[3705]), .B(p_input[33705]), .Z(n13989) );
  AND U20986 ( .A(n13991), .B(n13992), .Z(o[3704]) );
  AND U20987 ( .A(p_input[23704]), .B(p_input[13704]), .Z(n13992) );
  AND U20988 ( .A(p_input[3704]), .B(p_input[33704]), .Z(n13991) );
  AND U20989 ( .A(n13993), .B(n13994), .Z(o[3703]) );
  AND U20990 ( .A(p_input[23703]), .B(p_input[13703]), .Z(n13994) );
  AND U20991 ( .A(p_input[3703]), .B(p_input[33703]), .Z(n13993) );
  AND U20992 ( .A(n13995), .B(n13996), .Z(o[3702]) );
  AND U20993 ( .A(p_input[23702]), .B(p_input[13702]), .Z(n13996) );
  AND U20994 ( .A(p_input[3702]), .B(p_input[33702]), .Z(n13995) );
  AND U20995 ( .A(n13997), .B(n13998), .Z(o[3701]) );
  AND U20996 ( .A(p_input[23701]), .B(p_input[13701]), .Z(n13998) );
  AND U20997 ( .A(p_input[3701]), .B(p_input[33701]), .Z(n13997) );
  AND U20998 ( .A(n13999), .B(n14000), .Z(o[3700]) );
  AND U20999 ( .A(p_input[23700]), .B(p_input[13700]), .Z(n14000) );
  AND U21000 ( .A(p_input[3700]), .B(p_input[33700]), .Z(n13999) );
  AND U21001 ( .A(n14001), .B(n14002), .Z(o[36]) );
  AND U21002 ( .A(p_input[20036]), .B(p_input[10036]), .Z(n14002) );
  AND U21003 ( .A(p_input[36]), .B(p_input[30036]), .Z(n14001) );
  AND U21004 ( .A(n14003), .B(n14004), .Z(o[369]) );
  AND U21005 ( .A(p_input[20369]), .B(p_input[10369]), .Z(n14004) );
  AND U21006 ( .A(p_input[369]), .B(p_input[30369]), .Z(n14003) );
  AND U21007 ( .A(n14005), .B(n14006), .Z(o[3699]) );
  AND U21008 ( .A(p_input[23699]), .B(p_input[13699]), .Z(n14006) );
  AND U21009 ( .A(p_input[3699]), .B(p_input[33699]), .Z(n14005) );
  AND U21010 ( .A(n14007), .B(n14008), .Z(o[3698]) );
  AND U21011 ( .A(p_input[23698]), .B(p_input[13698]), .Z(n14008) );
  AND U21012 ( .A(p_input[3698]), .B(p_input[33698]), .Z(n14007) );
  AND U21013 ( .A(n14009), .B(n14010), .Z(o[3697]) );
  AND U21014 ( .A(p_input[23697]), .B(p_input[13697]), .Z(n14010) );
  AND U21015 ( .A(p_input[3697]), .B(p_input[33697]), .Z(n14009) );
  AND U21016 ( .A(n14011), .B(n14012), .Z(o[3696]) );
  AND U21017 ( .A(p_input[23696]), .B(p_input[13696]), .Z(n14012) );
  AND U21018 ( .A(p_input[3696]), .B(p_input[33696]), .Z(n14011) );
  AND U21019 ( .A(n14013), .B(n14014), .Z(o[3695]) );
  AND U21020 ( .A(p_input[23695]), .B(p_input[13695]), .Z(n14014) );
  AND U21021 ( .A(p_input[3695]), .B(p_input[33695]), .Z(n14013) );
  AND U21022 ( .A(n14015), .B(n14016), .Z(o[3694]) );
  AND U21023 ( .A(p_input[23694]), .B(p_input[13694]), .Z(n14016) );
  AND U21024 ( .A(p_input[3694]), .B(p_input[33694]), .Z(n14015) );
  AND U21025 ( .A(n14017), .B(n14018), .Z(o[3693]) );
  AND U21026 ( .A(p_input[23693]), .B(p_input[13693]), .Z(n14018) );
  AND U21027 ( .A(p_input[3693]), .B(p_input[33693]), .Z(n14017) );
  AND U21028 ( .A(n14019), .B(n14020), .Z(o[3692]) );
  AND U21029 ( .A(p_input[23692]), .B(p_input[13692]), .Z(n14020) );
  AND U21030 ( .A(p_input[3692]), .B(p_input[33692]), .Z(n14019) );
  AND U21031 ( .A(n14021), .B(n14022), .Z(o[3691]) );
  AND U21032 ( .A(p_input[23691]), .B(p_input[13691]), .Z(n14022) );
  AND U21033 ( .A(p_input[3691]), .B(p_input[33691]), .Z(n14021) );
  AND U21034 ( .A(n14023), .B(n14024), .Z(o[3690]) );
  AND U21035 ( .A(p_input[23690]), .B(p_input[13690]), .Z(n14024) );
  AND U21036 ( .A(p_input[3690]), .B(p_input[33690]), .Z(n14023) );
  AND U21037 ( .A(n14025), .B(n14026), .Z(o[368]) );
  AND U21038 ( .A(p_input[20368]), .B(p_input[10368]), .Z(n14026) );
  AND U21039 ( .A(p_input[368]), .B(p_input[30368]), .Z(n14025) );
  AND U21040 ( .A(n14027), .B(n14028), .Z(o[3689]) );
  AND U21041 ( .A(p_input[23689]), .B(p_input[13689]), .Z(n14028) );
  AND U21042 ( .A(p_input[3689]), .B(p_input[33689]), .Z(n14027) );
  AND U21043 ( .A(n14029), .B(n14030), .Z(o[3688]) );
  AND U21044 ( .A(p_input[23688]), .B(p_input[13688]), .Z(n14030) );
  AND U21045 ( .A(p_input[3688]), .B(p_input[33688]), .Z(n14029) );
  AND U21046 ( .A(n14031), .B(n14032), .Z(o[3687]) );
  AND U21047 ( .A(p_input[23687]), .B(p_input[13687]), .Z(n14032) );
  AND U21048 ( .A(p_input[3687]), .B(p_input[33687]), .Z(n14031) );
  AND U21049 ( .A(n14033), .B(n14034), .Z(o[3686]) );
  AND U21050 ( .A(p_input[23686]), .B(p_input[13686]), .Z(n14034) );
  AND U21051 ( .A(p_input[3686]), .B(p_input[33686]), .Z(n14033) );
  AND U21052 ( .A(n14035), .B(n14036), .Z(o[3685]) );
  AND U21053 ( .A(p_input[23685]), .B(p_input[13685]), .Z(n14036) );
  AND U21054 ( .A(p_input[3685]), .B(p_input[33685]), .Z(n14035) );
  AND U21055 ( .A(n14037), .B(n14038), .Z(o[3684]) );
  AND U21056 ( .A(p_input[23684]), .B(p_input[13684]), .Z(n14038) );
  AND U21057 ( .A(p_input[3684]), .B(p_input[33684]), .Z(n14037) );
  AND U21058 ( .A(n14039), .B(n14040), .Z(o[3683]) );
  AND U21059 ( .A(p_input[23683]), .B(p_input[13683]), .Z(n14040) );
  AND U21060 ( .A(p_input[3683]), .B(p_input[33683]), .Z(n14039) );
  AND U21061 ( .A(n14041), .B(n14042), .Z(o[3682]) );
  AND U21062 ( .A(p_input[23682]), .B(p_input[13682]), .Z(n14042) );
  AND U21063 ( .A(p_input[3682]), .B(p_input[33682]), .Z(n14041) );
  AND U21064 ( .A(n14043), .B(n14044), .Z(o[3681]) );
  AND U21065 ( .A(p_input[23681]), .B(p_input[13681]), .Z(n14044) );
  AND U21066 ( .A(p_input[3681]), .B(p_input[33681]), .Z(n14043) );
  AND U21067 ( .A(n14045), .B(n14046), .Z(o[3680]) );
  AND U21068 ( .A(p_input[23680]), .B(p_input[13680]), .Z(n14046) );
  AND U21069 ( .A(p_input[3680]), .B(p_input[33680]), .Z(n14045) );
  AND U21070 ( .A(n14047), .B(n14048), .Z(o[367]) );
  AND U21071 ( .A(p_input[20367]), .B(p_input[10367]), .Z(n14048) );
  AND U21072 ( .A(p_input[367]), .B(p_input[30367]), .Z(n14047) );
  AND U21073 ( .A(n14049), .B(n14050), .Z(o[3679]) );
  AND U21074 ( .A(p_input[23679]), .B(p_input[13679]), .Z(n14050) );
  AND U21075 ( .A(p_input[3679]), .B(p_input[33679]), .Z(n14049) );
  AND U21076 ( .A(n14051), .B(n14052), .Z(o[3678]) );
  AND U21077 ( .A(p_input[23678]), .B(p_input[13678]), .Z(n14052) );
  AND U21078 ( .A(p_input[3678]), .B(p_input[33678]), .Z(n14051) );
  AND U21079 ( .A(n14053), .B(n14054), .Z(o[3677]) );
  AND U21080 ( .A(p_input[23677]), .B(p_input[13677]), .Z(n14054) );
  AND U21081 ( .A(p_input[3677]), .B(p_input[33677]), .Z(n14053) );
  AND U21082 ( .A(n14055), .B(n14056), .Z(o[3676]) );
  AND U21083 ( .A(p_input[23676]), .B(p_input[13676]), .Z(n14056) );
  AND U21084 ( .A(p_input[3676]), .B(p_input[33676]), .Z(n14055) );
  AND U21085 ( .A(n14057), .B(n14058), .Z(o[3675]) );
  AND U21086 ( .A(p_input[23675]), .B(p_input[13675]), .Z(n14058) );
  AND U21087 ( .A(p_input[3675]), .B(p_input[33675]), .Z(n14057) );
  AND U21088 ( .A(n14059), .B(n14060), .Z(o[3674]) );
  AND U21089 ( .A(p_input[23674]), .B(p_input[13674]), .Z(n14060) );
  AND U21090 ( .A(p_input[3674]), .B(p_input[33674]), .Z(n14059) );
  AND U21091 ( .A(n14061), .B(n14062), .Z(o[3673]) );
  AND U21092 ( .A(p_input[23673]), .B(p_input[13673]), .Z(n14062) );
  AND U21093 ( .A(p_input[3673]), .B(p_input[33673]), .Z(n14061) );
  AND U21094 ( .A(n14063), .B(n14064), .Z(o[3672]) );
  AND U21095 ( .A(p_input[23672]), .B(p_input[13672]), .Z(n14064) );
  AND U21096 ( .A(p_input[3672]), .B(p_input[33672]), .Z(n14063) );
  AND U21097 ( .A(n14065), .B(n14066), .Z(o[3671]) );
  AND U21098 ( .A(p_input[23671]), .B(p_input[13671]), .Z(n14066) );
  AND U21099 ( .A(p_input[3671]), .B(p_input[33671]), .Z(n14065) );
  AND U21100 ( .A(n14067), .B(n14068), .Z(o[3670]) );
  AND U21101 ( .A(p_input[23670]), .B(p_input[13670]), .Z(n14068) );
  AND U21102 ( .A(p_input[3670]), .B(p_input[33670]), .Z(n14067) );
  AND U21103 ( .A(n14069), .B(n14070), .Z(o[366]) );
  AND U21104 ( .A(p_input[20366]), .B(p_input[10366]), .Z(n14070) );
  AND U21105 ( .A(p_input[366]), .B(p_input[30366]), .Z(n14069) );
  AND U21106 ( .A(n14071), .B(n14072), .Z(o[3669]) );
  AND U21107 ( .A(p_input[23669]), .B(p_input[13669]), .Z(n14072) );
  AND U21108 ( .A(p_input[3669]), .B(p_input[33669]), .Z(n14071) );
  AND U21109 ( .A(n14073), .B(n14074), .Z(o[3668]) );
  AND U21110 ( .A(p_input[23668]), .B(p_input[13668]), .Z(n14074) );
  AND U21111 ( .A(p_input[3668]), .B(p_input[33668]), .Z(n14073) );
  AND U21112 ( .A(n14075), .B(n14076), .Z(o[3667]) );
  AND U21113 ( .A(p_input[23667]), .B(p_input[13667]), .Z(n14076) );
  AND U21114 ( .A(p_input[3667]), .B(p_input[33667]), .Z(n14075) );
  AND U21115 ( .A(n14077), .B(n14078), .Z(o[3666]) );
  AND U21116 ( .A(p_input[23666]), .B(p_input[13666]), .Z(n14078) );
  AND U21117 ( .A(p_input[3666]), .B(p_input[33666]), .Z(n14077) );
  AND U21118 ( .A(n14079), .B(n14080), .Z(o[3665]) );
  AND U21119 ( .A(p_input[23665]), .B(p_input[13665]), .Z(n14080) );
  AND U21120 ( .A(p_input[3665]), .B(p_input[33665]), .Z(n14079) );
  AND U21121 ( .A(n14081), .B(n14082), .Z(o[3664]) );
  AND U21122 ( .A(p_input[23664]), .B(p_input[13664]), .Z(n14082) );
  AND U21123 ( .A(p_input[3664]), .B(p_input[33664]), .Z(n14081) );
  AND U21124 ( .A(n14083), .B(n14084), .Z(o[3663]) );
  AND U21125 ( .A(p_input[23663]), .B(p_input[13663]), .Z(n14084) );
  AND U21126 ( .A(p_input[3663]), .B(p_input[33663]), .Z(n14083) );
  AND U21127 ( .A(n14085), .B(n14086), .Z(o[3662]) );
  AND U21128 ( .A(p_input[23662]), .B(p_input[13662]), .Z(n14086) );
  AND U21129 ( .A(p_input[3662]), .B(p_input[33662]), .Z(n14085) );
  AND U21130 ( .A(n14087), .B(n14088), .Z(o[3661]) );
  AND U21131 ( .A(p_input[23661]), .B(p_input[13661]), .Z(n14088) );
  AND U21132 ( .A(p_input[3661]), .B(p_input[33661]), .Z(n14087) );
  AND U21133 ( .A(n14089), .B(n14090), .Z(o[3660]) );
  AND U21134 ( .A(p_input[23660]), .B(p_input[13660]), .Z(n14090) );
  AND U21135 ( .A(p_input[3660]), .B(p_input[33660]), .Z(n14089) );
  AND U21136 ( .A(n14091), .B(n14092), .Z(o[365]) );
  AND U21137 ( .A(p_input[20365]), .B(p_input[10365]), .Z(n14092) );
  AND U21138 ( .A(p_input[365]), .B(p_input[30365]), .Z(n14091) );
  AND U21139 ( .A(n14093), .B(n14094), .Z(o[3659]) );
  AND U21140 ( .A(p_input[23659]), .B(p_input[13659]), .Z(n14094) );
  AND U21141 ( .A(p_input[3659]), .B(p_input[33659]), .Z(n14093) );
  AND U21142 ( .A(n14095), .B(n14096), .Z(o[3658]) );
  AND U21143 ( .A(p_input[23658]), .B(p_input[13658]), .Z(n14096) );
  AND U21144 ( .A(p_input[3658]), .B(p_input[33658]), .Z(n14095) );
  AND U21145 ( .A(n14097), .B(n14098), .Z(o[3657]) );
  AND U21146 ( .A(p_input[23657]), .B(p_input[13657]), .Z(n14098) );
  AND U21147 ( .A(p_input[3657]), .B(p_input[33657]), .Z(n14097) );
  AND U21148 ( .A(n14099), .B(n14100), .Z(o[3656]) );
  AND U21149 ( .A(p_input[23656]), .B(p_input[13656]), .Z(n14100) );
  AND U21150 ( .A(p_input[3656]), .B(p_input[33656]), .Z(n14099) );
  AND U21151 ( .A(n14101), .B(n14102), .Z(o[3655]) );
  AND U21152 ( .A(p_input[23655]), .B(p_input[13655]), .Z(n14102) );
  AND U21153 ( .A(p_input[3655]), .B(p_input[33655]), .Z(n14101) );
  AND U21154 ( .A(n14103), .B(n14104), .Z(o[3654]) );
  AND U21155 ( .A(p_input[23654]), .B(p_input[13654]), .Z(n14104) );
  AND U21156 ( .A(p_input[3654]), .B(p_input[33654]), .Z(n14103) );
  AND U21157 ( .A(n14105), .B(n14106), .Z(o[3653]) );
  AND U21158 ( .A(p_input[23653]), .B(p_input[13653]), .Z(n14106) );
  AND U21159 ( .A(p_input[3653]), .B(p_input[33653]), .Z(n14105) );
  AND U21160 ( .A(n14107), .B(n14108), .Z(o[3652]) );
  AND U21161 ( .A(p_input[23652]), .B(p_input[13652]), .Z(n14108) );
  AND U21162 ( .A(p_input[3652]), .B(p_input[33652]), .Z(n14107) );
  AND U21163 ( .A(n14109), .B(n14110), .Z(o[3651]) );
  AND U21164 ( .A(p_input[23651]), .B(p_input[13651]), .Z(n14110) );
  AND U21165 ( .A(p_input[3651]), .B(p_input[33651]), .Z(n14109) );
  AND U21166 ( .A(n14111), .B(n14112), .Z(o[3650]) );
  AND U21167 ( .A(p_input[23650]), .B(p_input[13650]), .Z(n14112) );
  AND U21168 ( .A(p_input[3650]), .B(p_input[33650]), .Z(n14111) );
  AND U21169 ( .A(n14113), .B(n14114), .Z(o[364]) );
  AND U21170 ( .A(p_input[20364]), .B(p_input[10364]), .Z(n14114) );
  AND U21171 ( .A(p_input[364]), .B(p_input[30364]), .Z(n14113) );
  AND U21172 ( .A(n14115), .B(n14116), .Z(o[3649]) );
  AND U21173 ( .A(p_input[23649]), .B(p_input[13649]), .Z(n14116) );
  AND U21174 ( .A(p_input[3649]), .B(p_input[33649]), .Z(n14115) );
  AND U21175 ( .A(n14117), .B(n14118), .Z(o[3648]) );
  AND U21176 ( .A(p_input[23648]), .B(p_input[13648]), .Z(n14118) );
  AND U21177 ( .A(p_input[3648]), .B(p_input[33648]), .Z(n14117) );
  AND U21178 ( .A(n14119), .B(n14120), .Z(o[3647]) );
  AND U21179 ( .A(p_input[23647]), .B(p_input[13647]), .Z(n14120) );
  AND U21180 ( .A(p_input[3647]), .B(p_input[33647]), .Z(n14119) );
  AND U21181 ( .A(n14121), .B(n14122), .Z(o[3646]) );
  AND U21182 ( .A(p_input[23646]), .B(p_input[13646]), .Z(n14122) );
  AND U21183 ( .A(p_input[3646]), .B(p_input[33646]), .Z(n14121) );
  AND U21184 ( .A(n14123), .B(n14124), .Z(o[3645]) );
  AND U21185 ( .A(p_input[23645]), .B(p_input[13645]), .Z(n14124) );
  AND U21186 ( .A(p_input[3645]), .B(p_input[33645]), .Z(n14123) );
  AND U21187 ( .A(n14125), .B(n14126), .Z(o[3644]) );
  AND U21188 ( .A(p_input[23644]), .B(p_input[13644]), .Z(n14126) );
  AND U21189 ( .A(p_input[3644]), .B(p_input[33644]), .Z(n14125) );
  AND U21190 ( .A(n14127), .B(n14128), .Z(o[3643]) );
  AND U21191 ( .A(p_input[23643]), .B(p_input[13643]), .Z(n14128) );
  AND U21192 ( .A(p_input[3643]), .B(p_input[33643]), .Z(n14127) );
  AND U21193 ( .A(n14129), .B(n14130), .Z(o[3642]) );
  AND U21194 ( .A(p_input[23642]), .B(p_input[13642]), .Z(n14130) );
  AND U21195 ( .A(p_input[3642]), .B(p_input[33642]), .Z(n14129) );
  AND U21196 ( .A(n14131), .B(n14132), .Z(o[3641]) );
  AND U21197 ( .A(p_input[23641]), .B(p_input[13641]), .Z(n14132) );
  AND U21198 ( .A(p_input[3641]), .B(p_input[33641]), .Z(n14131) );
  AND U21199 ( .A(n14133), .B(n14134), .Z(o[3640]) );
  AND U21200 ( .A(p_input[23640]), .B(p_input[13640]), .Z(n14134) );
  AND U21201 ( .A(p_input[3640]), .B(p_input[33640]), .Z(n14133) );
  AND U21202 ( .A(n14135), .B(n14136), .Z(o[363]) );
  AND U21203 ( .A(p_input[20363]), .B(p_input[10363]), .Z(n14136) );
  AND U21204 ( .A(p_input[363]), .B(p_input[30363]), .Z(n14135) );
  AND U21205 ( .A(n14137), .B(n14138), .Z(o[3639]) );
  AND U21206 ( .A(p_input[23639]), .B(p_input[13639]), .Z(n14138) );
  AND U21207 ( .A(p_input[3639]), .B(p_input[33639]), .Z(n14137) );
  AND U21208 ( .A(n14139), .B(n14140), .Z(o[3638]) );
  AND U21209 ( .A(p_input[23638]), .B(p_input[13638]), .Z(n14140) );
  AND U21210 ( .A(p_input[3638]), .B(p_input[33638]), .Z(n14139) );
  AND U21211 ( .A(n14141), .B(n14142), .Z(o[3637]) );
  AND U21212 ( .A(p_input[23637]), .B(p_input[13637]), .Z(n14142) );
  AND U21213 ( .A(p_input[3637]), .B(p_input[33637]), .Z(n14141) );
  AND U21214 ( .A(n14143), .B(n14144), .Z(o[3636]) );
  AND U21215 ( .A(p_input[23636]), .B(p_input[13636]), .Z(n14144) );
  AND U21216 ( .A(p_input[3636]), .B(p_input[33636]), .Z(n14143) );
  AND U21217 ( .A(n14145), .B(n14146), .Z(o[3635]) );
  AND U21218 ( .A(p_input[23635]), .B(p_input[13635]), .Z(n14146) );
  AND U21219 ( .A(p_input[3635]), .B(p_input[33635]), .Z(n14145) );
  AND U21220 ( .A(n14147), .B(n14148), .Z(o[3634]) );
  AND U21221 ( .A(p_input[23634]), .B(p_input[13634]), .Z(n14148) );
  AND U21222 ( .A(p_input[3634]), .B(p_input[33634]), .Z(n14147) );
  AND U21223 ( .A(n14149), .B(n14150), .Z(o[3633]) );
  AND U21224 ( .A(p_input[23633]), .B(p_input[13633]), .Z(n14150) );
  AND U21225 ( .A(p_input[3633]), .B(p_input[33633]), .Z(n14149) );
  AND U21226 ( .A(n14151), .B(n14152), .Z(o[3632]) );
  AND U21227 ( .A(p_input[23632]), .B(p_input[13632]), .Z(n14152) );
  AND U21228 ( .A(p_input[3632]), .B(p_input[33632]), .Z(n14151) );
  AND U21229 ( .A(n14153), .B(n14154), .Z(o[3631]) );
  AND U21230 ( .A(p_input[23631]), .B(p_input[13631]), .Z(n14154) );
  AND U21231 ( .A(p_input[3631]), .B(p_input[33631]), .Z(n14153) );
  AND U21232 ( .A(n14155), .B(n14156), .Z(o[3630]) );
  AND U21233 ( .A(p_input[23630]), .B(p_input[13630]), .Z(n14156) );
  AND U21234 ( .A(p_input[3630]), .B(p_input[33630]), .Z(n14155) );
  AND U21235 ( .A(n14157), .B(n14158), .Z(o[362]) );
  AND U21236 ( .A(p_input[20362]), .B(p_input[10362]), .Z(n14158) );
  AND U21237 ( .A(p_input[362]), .B(p_input[30362]), .Z(n14157) );
  AND U21238 ( .A(n14159), .B(n14160), .Z(o[3629]) );
  AND U21239 ( .A(p_input[23629]), .B(p_input[13629]), .Z(n14160) );
  AND U21240 ( .A(p_input[3629]), .B(p_input[33629]), .Z(n14159) );
  AND U21241 ( .A(n14161), .B(n14162), .Z(o[3628]) );
  AND U21242 ( .A(p_input[23628]), .B(p_input[13628]), .Z(n14162) );
  AND U21243 ( .A(p_input[3628]), .B(p_input[33628]), .Z(n14161) );
  AND U21244 ( .A(n14163), .B(n14164), .Z(o[3627]) );
  AND U21245 ( .A(p_input[23627]), .B(p_input[13627]), .Z(n14164) );
  AND U21246 ( .A(p_input[3627]), .B(p_input[33627]), .Z(n14163) );
  AND U21247 ( .A(n14165), .B(n14166), .Z(o[3626]) );
  AND U21248 ( .A(p_input[23626]), .B(p_input[13626]), .Z(n14166) );
  AND U21249 ( .A(p_input[3626]), .B(p_input[33626]), .Z(n14165) );
  AND U21250 ( .A(n14167), .B(n14168), .Z(o[3625]) );
  AND U21251 ( .A(p_input[23625]), .B(p_input[13625]), .Z(n14168) );
  AND U21252 ( .A(p_input[3625]), .B(p_input[33625]), .Z(n14167) );
  AND U21253 ( .A(n14169), .B(n14170), .Z(o[3624]) );
  AND U21254 ( .A(p_input[23624]), .B(p_input[13624]), .Z(n14170) );
  AND U21255 ( .A(p_input[3624]), .B(p_input[33624]), .Z(n14169) );
  AND U21256 ( .A(n14171), .B(n14172), .Z(o[3623]) );
  AND U21257 ( .A(p_input[23623]), .B(p_input[13623]), .Z(n14172) );
  AND U21258 ( .A(p_input[3623]), .B(p_input[33623]), .Z(n14171) );
  AND U21259 ( .A(n14173), .B(n14174), .Z(o[3622]) );
  AND U21260 ( .A(p_input[23622]), .B(p_input[13622]), .Z(n14174) );
  AND U21261 ( .A(p_input[3622]), .B(p_input[33622]), .Z(n14173) );
  AND U21262 ( .A(n14175), .B(n14176), .Z(o[3621]) );
  AND U21263 ( .A(p_input[23621]), .B(p_input[13621]), .Z(n14176) );
  AND U21264 ( .A(p_input[3621]), .B(p_input[33621]), .Z(n14175) );
  AND U21265 ( .A(n14177), .B(n14178), .Z(o[3620]) );
  AND U21266 ( .A(p_input[23620]), .B(p_input[13620]), .Z(n14178) );
  AND U21267 ( .A(p_input[3620]), .B(p_input[33620]), .Z(n14177) );
  AND U21268 ( .A(n14179), .B(n14180), .Z(o[361]) );
  AND U21269 ( .A(p_input[20361]), .B(p_input[10361]), .Z(n14180) );
  AND U21270 ( .A(p_input[361]), .B(p_input[30361]), .Z(n14179) );
  AND U21271 ( .A(n14181), .B(n14182), .Z(o[3619]) );
  AND U21272 ( .A(p_input[23619]), .B(p_input[13619]), .Z(n14182) );
  AND U21273 ( .A(p_input[3619]), .B(p_input[33619]), .Z(n14181) );
  AND U21274 ( .A(n14183), .B(n14184), .Z(o[3618]) );
  AND U21275 ( .A(p_input[23618]), .B(p_input[13618]), .Z(n14184) );
  AND U21276 ( .A(p_input[3618]), .B(p_input[33618]), .Z(n14183) );
  AND U21277 ( .A(n14185), .B(n14186), .Z(o[3617]) );
  AND U21278 ( .A(p_input[23617]), .B(p_input[13617]), .Z(n14186) );
  AND U21279 ( .A(p_input[3617]), .B(p_input[33617]), .Z(n14185) );
  AND U21280 ( .A(n14187), .B(n14188), .Z(o[3616]) );
  AND U21281 ( .A(p_input[23616]), .B(p_input[13616]), .Z(n14188) );
  AND U21282 ( .A(p_input[3616]), .B(p_input[33616]), .Z(n14187) );
  AND U21283 ( .A(n14189), .B(n14190), .Z(o[3615]) );
  AND U21284 ( .A(p_input[23615]), .B(p_input[13615]), .Z(n14190) );
  AND U21285 ( .A(p_input[3615]), .B(p_input[33615]), .Z(n14189) );
  AND U21286 ( .A(n14191), .B(n14192), .Z(o[3614]) );
  AND U21287 ( .A(p_input[23614]), .B(p_input[13614]), .Z(n14192) );
  AND U21288 ( .A(p_input[3614]), .B(p_input[33614]), .Z(n14191) );
  AND U21289 ( .A(n14193), .B(n14194), .Z(o[3613]) );
  AND U21290 ( .A(p_input[23613]), .B(p_input[13613]), .Z(n14194) );
  AND U21291 ( .A(p_input[3613]), .B(p_input[33613]), .Z(n14193) );
  AND U21292 ( .A(n14195), .B(n14196), .Z(o[3612]) );
  AND U21293 ( .A(p_input[23612]), .B(p_input[13612]), .Z(n14196) );
  AND U21294 ( .A(p_input[3612]), .B(p_input[33612]), .Z(n14195) );
  AND U21295 ( .A(n14197), .B(n14198), .Z(o[3611]) );
  AND U21296 ( .A(p_input[23611]), .B(p_input[13611]), .Z(n14198) );
  AND U21297 ( .A(p_input[3611]), .B(p_input[33611]), .Z(n14197) );
  AND U21298 ( .A(n14199), .B(n14200), .Z(o[3610]) );
  AND U21299 ( .A(p_input[23610]), .B(p_input[13610]), .Z(n14200) );
  AND U21300 ( .A(p_input[3610]), .B(p_input[33610]), .Z(n14199) );
  AND U21301 ( .A(n14201), .B(n14202), .Z(o[360]) );
  AND U21302 ( .A(p_input[20360]), .B(p_input[10360]), .Z(n14202) );
  AND U21303 ( .A(p_input[360]), .B(p_input[30360]), .Z(n14201) );
  AND U21304 ( .A(n14203), .B(n14204), .Z(o[3609]) );
  AND U21305 ( .A(p_input[23609]), .B(p_input[13609]), .Z(n14204) );
  AND U21306 ( .A(p_input[3609]), .B(p_input[33609]), .Z(n14203) );
  AND U21307 ( .A(n14205), .B(n14206), .Z(o[3608]) );
  AND U21308 ( .A(p_input[23608]), .B(p_input[13608]), .Z(n14206) );
  AND U21309 ( .A(p_input[3608]), .B(p_input[33608]), .Z(n14205) );
  AND U21310 ( .A(n14207), .B(n14208), .Z(o[3607]) );
  AND U21311 ( .A(p_input[23607]), .B(p_input[13607]), .Z(n14208) );
  AND U21312 ( .A(p_input[3607]), .B(p_input[33607]), .Z(n14207) );
  AND U21313 ( .A(n14209), .B(n14210), .Z(o[3606]) );
  AND U21314 ( .A(p_input[23606]), .B(p_input[13606]), .Z(n14210) );
  AND U21315 ( .A(p_input[3606]), .B(p_input[33606]), .Z(n14209) );
  AND U21316 ( .A(n14211), .B(n14212), .Z(o[3605]) );
  AND U21317 ( .A(p_input[23605]), .B(p_input[13605]), .Z(n14212) );
  AND U21318 ( .A(p_input[3605]), .B(p_input[33605]), .Z(n14211) );
  AND U21319 ( .A(n14213), .B(n14214), .Z(o[3604]) );
  AND U21320 ( .A(p_input[23604]), .B(p_input[13604]), .Z(n14214) );
  AND U21321 ( .A(p_input[3604]), .B(p_input[33604]), .Z(n14213) );
  AND U21322 ( .A(n14215), .B(n14216), .Z(o[3603]) );
  AND U21323 ( .A(p_input[23603]), .B(p_input[13603]), .Z(n14216) );
  AND U21324 ( .A(p_input[3603]), .B(p_input[33603]), .Z(n14215) );
  AND U21325 ( .A(n14217), .B(n14218), .Z(o[3602]) );
  AND U21326 ( .A(p_input[23602]), .B(p_input[13602]), .Z(n14218) );
  AND U21327 ( .A(p_input[3602]), .B(p_input[33602]), .Z(n14217) );
  AND U21328 ( .A(n14219), .B(n14220), .Z(o[3601]) );
  AND U21329 ( .A(p_input[23601]), .B(p_input[13601]), .Z(n14220) );
  AND U21330 ( .A(p_input[3601]), .B(p_input[33601]), .Z(n14219) );
  AND U21331 ( .A(n14221), .B(n14222), .Z(o[3600]) );
  AND U21332 ( .A(p_input[23600]), .B(p_input[13600]), .Z(n14222) );
  AND U21333 ( .A(p_input[3600]), .B(p_input[33600]), .Z(n14221) );
  AND U21334 ( .A(n14223), .B(n14224), .Z(o[35]) );
  AND U21335 ( .A(p_input[20035]), .B(p_input[10035]), .Z(n14224) );
  AND U21336 ( .A(p_input[35]), .B(p_input[30035]), .Z(n14223) );
  AND U21337 ( .A(n14225), .B(n14226), .Z(o[359]) );
  AND U21338 ( .A(p_input[20359]), .B(p_input[10359]), .Z(n14226) );
  AND U21339 ( .A(p_input[359]), .B(p_input[30359]), .Z(n14225) );
  AND U21340 ( .A(n14227), .B(n14228), .Z(o[3599]) );
  AND U21341 ( .A(p_input[23599]), .B(p_input[13599]), .Z(n14228) );
  AND U21342 ( .A(p_input[3599]), .B(p_input[33599]), .Z(n14227) );
  AND U21343 ( .A(n14229), .B(n14230), .Z(o[3598]) );
  AND U21344 ( .A(p_input[23598]), .B(p_input[13598]), .Z(n14230) );
  AND U21345 ( .A(p_input[3598]), .B(p_input[33598]), .Z(n14229) );
  AND U21346 ( .A(n14231), .B(n14232), .Z(o[3597]) );
  AND U21347 ( .A(p_input[23597]), .B(p_input[13597]), .Z(n14232) );
  AND U21348 ( .A(p_input[3597]), .B(p_input[33597]), .Z(n14231) );
  AND U21349 ( .A(n14233), .B(n14234), .Z(o[3596]) );
  AND U21350 ( .A(p_input[23596]), .B(p_input[13596]), .Z(n14234) );
  AND U21351 ( .A(p_input[3596]), .B(p_input[33596]), .Z(n14233) );
  AND U21352 ( .A(n14235), .B(n14236), .Z(o[3595]) );
  AND U21353 ( .A(p_input[23595]), .B(p_input[13595]), .Z(n14236) );
  AND U21354 ( .A(p_input[3595]), .B(p_input[33595]), .Z(n14235) );
  AND U21355 ( .A(n14237), .B(n14238), .Z(o[3594]) );
  AND U21356 ( .A(p_input[23594]), .B(p_input[13594]), .Z(n14238) );
  AND U21357 ( .A(p_input[3594]), .B(p_input[33594]), .Z(n14237) );
  AND U21358 ( .A(n14239), .B(n14240), .Z(o[3593]) );
  AND U21359 ( .A(p_input[23593]), .B(p_input[13593]), .Z(n14240) );
  AND U21360 ( .A(p_input[3593]), .B(p_input[33593]), .Z(n14239) );
  AND U21361 ( .A(n14241), .B(n14242), .Z(o[3592]) );
  AND U21362 ( .A(p_input[23592]), .B(p_input[13592]), .Z(n14242) );
  AND U21363 ( .A(p_input[3592]), .B(p_input[33592]), .Z(n14241) );
  AND U21364 ( .A(n14243), .B(n14244), .Z(o[3591]) );
  AND U21365 ( .A(p_input[23591]), .B(p_input[13591]), .Z(n14244) );
  AND U21366 ( .A(p_input[3591]), .B(p_input[33591]), .Z(n14243) );
  AND U21367 ( .A(n14245), .B(n14246), .Z(o[3590]) );
  AND U21368 ( .A(p_input[23590]), .B(p_input[13590]), .Z(n14246) );
  AND U21369 ( .A(p_input[3590]), .B(p_input[33590]), .Z(n14245) );
  AND U21370 ( .A(n14247), .B(n14248), .Z(o[358]) );
  AND U21371 ( .A(p_input[20358]), .B(p_input[10358]), .Z(n14248) );
  AND U21372 ( .A(p_input[358]), .B(p_input[30358]), .Z(n14247) );
  AND U21373 ( .A(n14249), .B(n14250), .Z(o[3589]) );
  AND U21374 ( .A(p_input[23589]), .B(p_input[13589]), .Z(n14250) );
  AND U21375 ( .A(p_input[3589]), .B(p_input[33589]), .Z(n14249) );
  AND U21376 ( .A(n14251), .B(n14252), .Z(o[3588]) );
  AND U21377 ( .A(p_input[23588]), .B(p_input[13588]), .Z(n14252) );
  AND U21378 ( .A(p_input[3588]), .B(p_input[33588]), .Z(n14251) );
  AND U21379 ( .A(n14253), .B(n14254), .Z(o[3587]) );
  AND U21380 ( .A(p_input[23587]), .B(p_input[13587]), .Z(n14254) );
  AND U21381 ( .A(p_input[3587]), .B(p_input[33587]), .Z(n14253) );
  AND U21382 ( .A(n14255), .B(n14256), .Z(o[3586]) );
  AND U21383 ( .A(p_input[23586]), .B(p_input[13586]), .Z(n14256) );
  AND U21384 ( .A(p_input[3586]), .B(p_input[33586]), .Z(n14255) );
  AND U21385 ( .A(n14257), .B(n14258), .Z(o[3585]) );
  AND U21386 ( .A(p_input[23585]), .B(p_input[13585]), .Z(n14258) );
  AND U21387 ( .A(p_input[3585]), .B(p_input[33585]), .Z(n14257) );
  AND U21388 ( .A(n14259), .B(n14260), .Z(o[3584]) );
  AND U21389 ( .A(p_input[23584]), .B(p_input[13584]), .Z(n14260) );
  AND U21390 ( .A(p_input[3584]), .B(p_input[33584]), .Z(n14259) );
  AND U21391 ( .A(n14261), .B(n14262), .Z(o[3583]) );
  AND U21392 ( .A(p_input[23583]), .B(p_input[13583]), .Z(n14262) );
  AND U21393 ( .A(p_input[3583]), .B(p_input[33583]), .Z(n14261) );
  AND U21394 ( .A(n14263), .B(n14264), .Z(o[3582]) );
  AND U21395 ( .A(p_input[23582]), .B(p_input[13582]), .Z(n14264) );
  AND U21396 ( .A(p_input[3582]), .B(p_input[33582]), .Z(n14263) );
  AND U21397 ( .A(n14265), .B(n14266), .Z(o[3581]) );
  AND U21398 ( .A(p_input[23581]), .B(p_input[13581]), .Z(n14266) );
  AND U21399 ( .A(p_input[3581]), .B(p_input[33581]), .Z(n14265) );
  AND U21400 ( .A(n14267), .B(n14268), .Z(o[3580]) );
  AND U21401 ( .A(p_input[23580]), .B(p_input[13580]), .Z(n14268) );
  AND U21402 ( .A(p_input[3580]), .B(p_input[33580]), .Z(n14267) );
  AND U21403 ( .A(n14269), .B(n14270), .Z(o[357]) );
  AND U21404 ( .A(p_input[20357]), .B(p_input[10357]), .Z(n14270) );
  AND U21405 ( .A(p_input[357]), .B(p_input[30357]), .Z(n14269) );
  AND U21406 ( .A(n14271), .B(n14272), .Z(o[3579]) );
  AND U21407 ( .A(p_input[23579]), .B(p_input[13579]), .Z(n14272) );
  AND U21408 ( .A(p_input[3579]), .B(p_input[33579]), .Z(n14271) );
  AND U21409 ( .A(n14273), .B(n14274), .Z(o[3578]) );
  AND U21410 ( .A(p_input[23578]), .B(p_input[13578]), .Z(n14274) );
  AND U21411 ( .A(p_input[3578]), .B(p_input[33578]), .Z(n14273) );
  AND U21412 ( .A(n14275), .B(n14276), .Z(o[3577]) );
  AND U21413 ( .A(p_input[23577]), .B(p_input[13577]), .Z(n14276) );
  AND U21414 ( .A(p_input[3577]), .B(p_input[33577]), .Z(n14275) );
  AND U21415 ( .A(n14277), .B(n14278), .Z(o[3576]) );
  AND U21416 ( .A(p_input[23576]), .B(p_input[13576]), .Z(n14278) );
  AND U21417 ( .A(p_input[3576]), .B(p_input[33576]), .Z(n14277) );
  AND U21418 ( .A(n14279), .B(n14280), .Z(o[3575]) );
  AND U21419 ( .A(p_input[23575]), .B(p_input[13575]), .Z(n14280) );
  AND U21420 ( .A(p_input[3575]), .B(p_input[33575]), .Z(n14279) );
  AND U21421 ( .A(n14281), .B(n14282), .Z(o[3574]) );
  AND U21422 ( .A(p_input[23574]), .B(p_input[13574]), .Z(n14282) );
  AND U21423 ( .A(p_input[3574]), .B(p_input[33574]), .Z(n14281) );
  AND U21424 ( .A(n14283), .B(n14284), .Z(o[3573]) );
  AND U21425 ( .A(p_input[23573]), .B(p_input[13573]), .Z(n14284) );
  AND U21426 ( .A(p_input[3573]), .B(p_input[33573]), .Z(n14283) );
  AND U21427 ( .A(n14285), .B(n14286), .Z(o[3572]) );
  AND U21428 ( .A(p_input[23572]), .B(p_input[13572]), .Z(n14286) );
  AND U21429 ( .A(p_input[3572]), .B(p_input[33572]), .Z(n14285) );
  AND U21430 ( .A(n14287), .B(n14288), .Z(o[3571]) );
  AND U21431 ( .A(p_input[23571]), .B(p_input[13571]), .Z(n14288) );
  AND U21432 ( .A(p_input[3571]), .B(p_input[33571]), .Z(n14287) );
  AND U21433 ( .A(n14289), .B(n14290), .Z(o[3570]) );
  AND U21434 ( .A(p_input[23570]), .B(p_input[13570]), .Z(n14290) );
  AND U21435 ( .A(p_input[3570]), .B(p_input[33570]), .Z(n14289) );
  AND U21436 ( .A(n14291), .B(n14292), .Z(o[356]) );
  AND U21437 ( .A(p_input[20356]), .B(p_input[10356]), .Z(n14292) );
  AND U21438 ( .A(p_input[356]), .B(p_input[30356]), .Z(n14291) );
  AND U21439 ( .A(n14293), .B(n14294), .Z(o[3569]) );
  AND U21440 ( .A(p_input[23569]), .B(p_input[13569]), .Z(n14294) );
  AND U21441 ( .A(p_input[3569]), .B(p_input[33569]), .Z(n14293) );
  AND U21442 ( .A(n14295), .B(n14296), .Z(o[3568]) );
  AND U21443 ( .A(p_input[23568]), .B(p_input[13568]), .Z(n14296) );
  AND U21444 ( .A(p_input[3568]), .B(p_input[33568]), .Z(n14295) );
  AND U21445 ( .A(n14297), .B(n14298), .Z(o[3567]) );
  AND U21446 ( .A(p_input[23567]), .B(p_input[13567]), .Z(n14298) );
  AND U21447 ( .A(p_input[3567]), .B(p_input[33567]), .Z(n14297) );
  AND U21448 ( .A(n14299), .B(n14300), .Z(o[3566]) );
  AND U21449 ( .A(p_input[23566]), .B(p_input[13566]), .Z(n14300) );
  AND U21450 ( .A(p_input[3566]), .B(p_input[33566]), .Z(n14299) );
  AND U21451 ( .A(n14301), .B(n14302), .Z(o[3565]) );
  AND U21452 ( .A(p_input[23565]), .B(p_input[13565]), .Z(n14302) );
  AND U21453 ( .A(p_input[3565]), .B(p_input[33565]), .Z(n14301) );
  AND U21454 ( .A(n14303), .B(n14304), .Z(o[3564]) );
  AND U21455 ( .A(p_input[23564]), .B(p_input[13564]), .Z(n14304) );
  AND U21456 ( .A(p_input[3564]), .B(p_input[33564]), .Z(n14303) );
  AND U21457 ( .A(n14305), .B(n14306), .Z(o[3563]) );
  AND U21458 ( .A(p_input[23563]), .B(p_input[13563]), .Z(n14306) );
  AND U21459 ( .A(p_input[3563]), .B(p_input[33563]), .Z(n14305) );
  AND U21460 ( .A(n14307), .B(n14308), .Z(o[3562]) );
  AND U21461 ( .A(p_input[23562]), .B(p_input[13562]), .Z(n14308) );
  AND U21462 ( .A(p_input[3562]), .B(p_input[33562]), .Z(n14307) );
  AND U21463 ( .A(n14309), .B(n14310), .Z(o[3561]) );
  AND U21464 ( .A(p_input[23561]), .B(p_input[13561]), .Z(n14310) );
  AND U21465 ( .A(p_input[3561]), .B(p_input[33561]), .Z(n14309) );
  AND U21466 ( .A(n14311), .B(n14312), .Z(o[3560]) );
  AND U21467 ( .A(p_input[23560]), .B(p_input[13560]), .Z(n14312) );
  AND U21468 ( .A(p_input[3560]), .B(p_input[33560]), .Z(n14311) );
  AND U21469 ( .A(n14313), .B(n14314), .Z(o[355]) );
  AND U21470 ( .A(p_input[20355]), .B(p_input[10355]), .Z(n14314) );
  AND U21471 ( .A(p_input[355]), .B(p_input[30355]), .Z(n14313) );
  AND U21472 ( .A(n14315), .B(n14316), .Z(o[3559]) );
  AND U21473 ( .A(p_input[23559]), .B(p_input[13559]), .Z(n14316) );
  AND U21474 ( .A(p_input[3559]), .B(p_input[33559]), .Z(n14315) );
  AND U21475 ( .A(n14317), .B(n14318), .Z(o[3558]) );
  AND U21476 ( .A(p_input[23558]), .B(p_input[13558]), .Z(n14318) );
  AND U21477 ( .A(p_input[3558]), .B(p_input[33558]), .Z(n14317) );
  AND U21478 ( .A(n14319), .B(n14320), .Z(o[3557]) );
  AND U21479 ( .A(p_input[23557]), .B(p_input[13557]), .Z(n14320) );
  AND U21480 ( .A(p_input[3557]), .B(p_input[33557]), .Z(n14319) );
  AND U21481 ( .A(n14321), .B(n14322), .Z(o[3556]) );
  AND U21482 ( .A(p_input[23556]), .B(p_input[13556]), .Z(n14322) );
  AND U21483 ( .A(p_input[3556]), .B(p_input[33556]), .Z(n14321) );
  AND U21484 ( .A(n14323), .B(n14324), .Z(o[3555]) );
  AND U21485 ( .A(p_input[23555]), .B(p_input[13555]), .Z(n14324) );
  AND U21486 ( .A(p_input[3555]), .B(p_input[33555]), .Z(n14323) );
  AND U21487 ( .A(n14325), .B(n14326), .Z(o[3554]) );
  AND U21488 ( .A(p_input[23554]), .B(p_input[13554]), .Z(n14326) );
  AND U21489 ( .A(p_input[3554]), .B(p_input[33554]), .Z(n14325) );
  AND U21490 ( .A(n14327), .B(n14328), .Z(o[3553]) );
  AND U21491 ( .A(p_input[23553]), .B(p_input[13553]), .Z(n14328) );
  AND U21492 ( .A(p_input[3553]), .B(p_input[33553]), .Z(n14327) );
  AND U21493 ( .A(n14329), .B(n14330), .Z(o[3552]) );
  AND U21494 ( .A(p_input[23552]), .B(p_input[13552]), .Z(n14330) );
  AND U21495 ( .A(p_input[3552]), .B(p_input[33552]), .Z(n14329) );
  AND U21496 ( .A(n14331), .B(n14332), .Z(o[3551]) );
  AND U21497 ( .A(p_input[23551]), .B(p_input[13551]), .Z(n14332) );
  AND U21498 ( .A(p_input[3551]), .B(p_input[33551]), .Z(n14331) );
  AND U21499 ( .A(n14333), .B(n14334), .Z(o[3550]) );
  AND U21500 ( .A(p_input[23550]), .B(p_input[13550]), .Z(n14334) );
  AND U21501 ( .A(p_input[3550]), .B(p_input[33550]), .Z(n14333) );
  AND U21502 ( .A(n14335), .B(n14336), .Z(o[354]) );
  AND U21503 ( .A(p_input[20354]), .B(p_input[10354]), .Z(n14336) );
  AND U21504 ( .A(p_input[354]), .B(p_input[30354]), .Z(n14335) );
  AND U21505 ( .A(n14337), .B(n14338), .Z(o[3549]) );
  AND U21506 ( .A(p_input[23549]), .B(p_input[13549]), .Z(n14338) );
  AND U21507 ( .A(p_input[3549]), .B(p_input[33549]), .Z(n14337) );
  AND U21508 ( .A(n14339), .B(n14340), .Z(o[3548]) );
  AND U21509 ( .A(p_input[23548]), .B(p_input[13548]), .Z(n14340) );
  AND U21510 ( .A(p_input[3548]), .B(p_input[33548]), .Z(n14339) );
  AND U21511 ( .A(n14341), .B(n14342), .Z(o[3547]) );
  AND U21512 ( .A(p_input[23547]), .B(p_input[13547]), .Z(n14342) );
  AND U21513 ( .A(p_input[3547]), .B(p_input[33547]), .Z(n14341) );
  AND U21514 ( .A(n14343), .B(n14344), .Z(o[3546]) );
  AND U21515 ( .A(p_input[23546]), .B(p_input[13546]), .Z(n14344) );
  AND U21516 ( .A(p_input[3546]), .B(p_input[33546]), .Z(n14343) );
  AND U21517 ( .A(n14345), .B(n14346), .Z(o[3545]) );
  AND U21518 ( .A(p_input[23545]), .B(p_input[13545]), .Z(n14346) );
  AND U21519 ( .A(p_input[3545]), .B(p_input[33545]), .Z(n14345) );
  AND U21520 ( .A(n14347), .B(n14348), .Z(o[3544]) );
  AND U21521 ( .A(p_input[23544]), .B(p_input[13544]), .Z(n14348) );
  AND U21522 ( .A(p_input[3544]), .B(p_input[33544]), .Z(n14347) );
  AND U21523 ( .A(n14349), .B(n14350), .Z(o[3543]) );
  AND U21524 ( .A(p_input[23543]), .B(p_input[13543]), .Z(n14350) );
  AND U21525 ( .A(p_input[3543]), .B(p_input[33543]), .Z(n14349) );
  AND U21526 ( .A(n14351), .B(n14352), .Z(o[3542]) );
  AND U21527 ( .A(p_input[23542]), .B(p_input[13542]), .Z(n14352) );
  AND U21528 ( .A(p_input[3542]), .B(p_input[33542]), .Z(n14351) );
  AND U21529 ( .A(n14353), .B(n14354), .Z(o[3541]) );
  AND U21530 ( .A(p_input[23541]), .B(p_input[13541]), .Z(n14354) );
  AND U21531 ( .A(p_input[3541]), .B(p_input[33541]), .Z(n14353) );
  AND U21532 ( .A(n14355), .B(n14356), .Z(o[3540]) );
  AND U21533 ( .A(p_input[23540]), .B(p_input[13540]), .Z(n14356) );
  AND U21534 ( .A(p_input[3540]), .B(p_input[33540]), .Z(n14355) );
  AND U21535 ( .A(n14357), .B(n14358), .Z(o[353]) );
  AND U21536 ( .A(p_input[20353]), .B(p_input[10353]), .Z(n14358) );
  AND U21537 ( .A(p_input[353]), .B(p_input[30353]), .Z(n14357) );
  AND U21538 ( .A(n14359), .B(n14360), .Z(o[3539]) );
  AND U21539 ( .A(p_input[23539]), .B(p_input[13539]), .Z(n14360) );
  AND U21540 ( .A(p_input[3539]), .B(p_input[33539]), .Z(n14359) );
  AND U21541 ( .A(n14361), .B(n14362), .Z(o[3538]) );
  AND U21542 ( .A(p_input[23538]), .B(p_input[13538]), .Z(n14362) );
  AND U21543 ( .A(p_input[3538]), .B(p_input[33538]), .Z(n14361) );
  AND U21544 ( .A(n14363), .B(n14364), .Z(o[3537]) );
  AND U21545 ( .A(p_input[23537]), .B(p_input[13537]), .Z(n14364) );
  AND U21546 ( .A(p_input[3537]), .B(p_input[33537]), .Z(n14363) );
  AND U21547 ( .A(n14365), .B(n14366), .Z(o[3536]) );
  AND U21548 ( .A(p_input[23536]), .B(p_input[13536]), .Z(n14366) );
  AND U21549 ( .A(p_input[3536]), .B(p_input[33536]), .Z(n14365) );
  AND U21550 ( .A(n14367), .B(n14368), .Z(o[3535]) );
  AND U21551 ( .A(p_input[23535]), .B(p_input[13535]), .Z(n14368) );
  AND U21552 ( .A(p_input[3535]), .B(p_input[33535]), .Z(n14367) );
  AND U21553 ( .A(n14369), .B(n14370), .Z(o[3534]) );
  AND U21554 ( .A(p_input[23534]), .B(p_input[13534]), .Z(n14370) );
  AND U21555 ( .A(p_input[3534]), .B(p_input[33534]), .Z(n14369) );
  AND U21556 ( .A(n14371), .B(n14372), .Z(o[3533]) );
  AND U21557 ( .A(p_input[23533]), .B(p_input[13533]), .Z(n14372) );
  AND U21558 ( .A(p_input[3533]), .B(p_input[33533]), .Z(n14371) );
  AND U21559 ( .A(n14373), .B(n14374), .Z(o[3532]) );
  AND U21560 ( .A(p_input[23532]), .B(p_input[13532]), .Z(n14374) );
  AND U21561 ( .A(p_input[3532]), .B(p_input[33532]), .Z(n14373) );
  AND U21562 ( .A(n14375), .B(n14376), .Z(o[3531]) );
  AND U21563 ( .A(p_input[23531]), .B(p_input[13531]), .Z(n14376) );
  AND U21564 ( .A(p_input[3531]), .B(p_input[33531]), .Z(n14375) );
  AND U21565 ( .A(n14377), .B(n14378), .Z(o[3530]) );
  AND U21566 ( .A(p_input[23530]), .B(p_input[13530]), .Z(n14378) );
  AND U21567 ( .A(p_input[3530]), .B(p_input[33530]), .Z(n14377) );
  AND U21568 ( .A(n14379), .B(n14380), .Z(o[352]) );
  AND U21569 ( .A(p_input[20352]), .B(p_input[10352]), .Z(n14380) );
  AND U21570 ( .A(p_input[352]), .B(p_input[30352]), .Z(n14379) );
  AND U21571 ( .A(n14381), .B(n14382), .Z(o[3529]) );
  AND U21572 ( .A(p_input[23529]), .B(p_input[13529]), .Z(n14382) );
  AND U21573 ( .A(p_input[3529]), .B(p_input[33529]), .Z(n14381) );
  AND U21574 ( .A(n14383), .B(n14384), .Z(o[3528]) );
  AND U21575 ( .A(p_input[23528]), .B(p_input[13528]), .Z(n14384) );
  AND U21576 ( .A(p_input[3528]), .B(p_input[33528]), .Z(n14383) );
  AND U21577 ( .A(n14385), .B(n14386), .Z(o[3527]) );
  AND U21578 ( .A(p_input[23527]), .B(p_input[13527]), .Z(n14386) );
  AND U21579 ( .A(p_input[3527]), .B(p_input[33527]), .Z(n14385) );
  AND U21580 ( .A(n14387), .B(n14388), .Z(o[3526]) );
  AND U21581 ( .A(p_input[23526]), .B(p_input[13526]), .Z(n14388) );
  AND U21582 ( .A(p_input[3526]), .B(p_input[33526]), .Z(n14387) );
  AND U21583 ( .A(n14389), .B(n14390), .Z(o[3525]) );
  AND U21584 ( .A(p_input[23525]), .B(p_input[13525]), .Z(n14390) );
  AND U21585 ( .A(p_input[3525]), .B(p_input[33525]), .Z(n14389) );
  AND U21586 ( .A(n14391), .B(n14392), .Z(o[3524]) );
  AND U21587 ( .A(p_input[23524]), .B(p_input[13524]), .Z(n14392) );
  AND U21588 ( .A(p_input[3524]), .B(p_input[33524]), .Z(n14391) );
  AND U21589 ( .A(n14393), .B(n14394), .Z(o[3523]) );
  AND U21590 ( .A(p_input[23523]), .B(p_input[13523]), .Z(n14394) );
  AND U21591 ( .A(p_input[3523]), .B(p_input[33523]), .Z(n14393) );
  AND U21592 ( .A(n14395), .B(n14396), .Z(o[3522]) );
  AND U21593 ( .A(p_input[23522]), .B(p_input[13522]), .Z(n14396) );
  AND U21594 ( .A(p_input[3522]), .B(p_input[33522]), .Z(n14395) );
  AND U21595 ( .A(n14397), .B(n14398), .Z(o[3521]) );
  AND U21596 ( .A(p_input[23521]), .B(p_input[13521]), .Z(n14398) );
  AND U21597 ( .A(p_input[3521]), .B(p_input[33521]), .Z(n14397) );
  AND U21598 ( .A(n14399), .B(n14400), .Z(o[3520]) );
  AND U21599 ( .A(p_input[23520]), .B(p_input[13520]), .Z(n14400) );
  AND U21600 ( .A(p_input[3520]), .B(p_input[33520]), .Z(n14399) );
  AND U21601 ( .A(n14401), .B(n14402), .Z(o[351]) );
  AND U21602 ( .A(p_input[20351]), .B(p_input[10351]), .Z(n14402) );
  AND U21603 ( .A(p_input[351]), .B(p_input[30351]), .Z(n14401) );
  AND U21604 ( .A(n14403), .B(n14404), .Z(o[3519]) );
  AND U21605 ( .A(p_input[23519]), .B(p_input[13519]), .Z(n14404) );
  AND U21606 ( .A(p_input[3519]), .B(p_input[33519]), .Z(n14403) );
  AND U21607 ( .A(n14405), .B(n14406), .Z(o[3518]) );
  AND U21608 ( .A(p_input[23518]), .B(p_input[13518]), .Z(n14406) );
  AND U21609 ( .A(p_input[3518]), .B(p_input[33518]), .Z(n14405) );
  AND U21610 ( .A(n14407), .B(n14408), .Z(o[3517]) );
  AND U21611 ( .A(p_input[23517]), .B(p_input[13517]), .Z(n14408) );
  AND U21612 ( .A(p_input[3517]), .B(p_input[33517]), .Z(n14407) );
  AND U21613 ( .A(n14409), .B(n14410), .Z(o[3516]) );
  AND U21614 ( .A(p_input[23516]), .B(p_input[13516]), .Z(n14410) );
  AND U21615 ( .A(p_input[3516]), .B(p_input[33516]), .Z(n14409) );
  AND U21616 ( .A(n14411), .B(n14412), .Z(o[3515]) );
  AND U21617 ( .A(p_input[23515]), .B(p_input[13515]), .Z(n14412) );
  AND U21618 ( .A(p_input[3515]), .B(p_input[33515]), .Z(n14411) );
  AND U21619 ( .A(n14413), .B(n14414), .Z(o[3514]) );
  AND U21620 ( .A(p_input[23514]), .B(p_input[13514]), .Z(n14414) );
  AND U21621 ( .A(p_input[3514]), .B(p_input[33514]), .Z(n14413) );
  AND U21622 ( .A(n14415), .B(n14416), .Z(o[3513]) );
  AND U21623 ( .A(p_input[23513]), .B(p_input[13513]), .Z(n14416) );
  AND U21624 ( .A(p_input[3513]), .B(p_input[33513]), .Z(n14415) );
  AND U21625 ( .A(n14417), .B(n14418), .Z(o[3512]) );
  AND U21626 ( .A(p_input[23512]), .B(p_input[13512]), .Z(n14418) );
  AND U21627 ( .A(p_input[3512]), .B(p_input[33512]), .Z(n14417) );
  AND U21628 ( .A(n14419), .B(n14420), .Z(o[3511]) );
  AND U21629 ( .A(p_input[23511]), .B(p_input[13511]), .Z(n14420) );
  AND U21630 ( .A(p_input[3511]), .B(p_input[33511]), .Z(n14419) );
  AND U21631 ( .A(n14421), .B(n14422), .Z(o[3510]) );
  AND U21632 ( .A(p_input[23510]), .B(p_input[13510]), .Z(n14422) );
  AND U21633 ( .A(p_input[3510]), .B(p_input[33510]), .Z(n14421) );
  AND U21634 ( .A(n14423), .B(n14424), .Z(o[350]) );
  AND U21635 ( .A(p_input[20350]), .B(p_input[10350]), .Z(n14424) );
  AND U21636 ( .A(p_input[350]), .B(p_input[30350]), .Z(n14423) );
  AND U21637 ( .A(n14425), .B(n14426), .Z(o[3509]) );
  AND U21638 ( .A(p_input[23509]), .B(p_input[13509]), .Z(n14426) );
  AND U21639 ( .A(p_input[3509]), .B(p_input[33509]), .Z(n14425) );
  AND U21640 ( .A(n14427), .B(n14428), .Z(o[3508]) );
  AND U21641 ( .A(p_input[23508]), .B(p_input[13508]), .Z(n14428) );
  AND U21642 ( .A(p_input[3508]), .B(p_input[33508]), .Z(n14427) );
  AND U21643 ( .A(n14429), .B(n14430), .Z(o[3507]) );
  AND U21644 ( .A(p_input[23507]), .B(p_input[13507]), .Z(n14430) );
  AND U21645 ( .A(p_input[3507]), .B(p_input[33507]), .Z(n14429) );
  AND U21646 ( .A(n14431), .B(n14432), .Z(o[3506]) );
  AND U21647 ( .A(p_input[23506]), .B(p_input[13506]), .Z(n14432) );
  AND U21648 ( .A(p_input[3506]), .B(p_input[33506]), .Z(n14431) );
  AND U21649 ( .A(n14433), .B(n14434), .Z(o[3505]) );
  AND U21650 ( .A(p_input[23505]), .B(p_input[13505]), .Z(n14434) );
  AND U21651 ( .A(p_input[3505]), .B(p_input[33505]), .Z(n14433) );
  AND U21652 ( .A(n14435), .B(n14436), .Z(o[3504]) );
  AND U21653 ( .A(p_input[23504]), .B(p_input[13504]), .Z(n14436) );
  AND U21654 ( .A(p_input[3504]), .B(p_input[33504]), .Z(n14435) );
  AND U21655 ( .A(n14437), .B(n14438), .Z(o[3503]) );
  AND U21656 ( .A(p_input[23503]), .B(p_input[13503]), .Z(n14438) );
  AND U21657 ( .A(p_input[3503]), .B(p_input[33503]), .Z(n14437) );
  AND U21658 ( .A(n14439), .B(n14440), .Z(o[3502]) );
  AND U21659 ( .A(p_input[23502]), .B(p_input[13502]), .Z(n14440) );
  AND U21660 ( .A(p_input[3502]), .B(p_input[33502]), .Z(n14439) );
  AND U21661 ( .A(n14441), .B(n14442), .Z(o[3501]) );
  AND U21662 ( .A(p_input[23501]), .B(p_input[13501]), .Z(n14442) );
  AND U21663 ( .A(p_input[3501]), .B(p_input[33501]), .Z(n14441) );
  AND U21664 ( .A(n14443), .B(n14444), .Z(o[3500]) );
  AND U21665 ( .A(p_input[23500]), .B(p_input[13500]), .Z(n14444) );
  AND U21666 ( .A(p_input[3500]), .B(p_input[33500]), .Z(n14443) );
  AND U21667 ( .A(n14445), .B(n14446), .Z(o[34]) );
  AND U21668 ( .A(p_input[20034]), .B(p_input[10034]), .Z(n14446) );
  AND U21669 ( .A(p_input[34]), .B(p_input[30034]), .Z(n14445) );
  AND U21670 ( .A(n14447), .B(n14448), .Z(o[349]) );
  AND U21671 ( .A(p_input[20349]), .B(p_input[10349]), .Z(n14448) );
  AND U21672 ( .A(p_input[349]), .B(p_input[30349]), .Z(n14447) );
  AND U21673 ( .A(n14449), .B(n14450), .Z(o[3499]) );
  AND U21674 ( .A(p_input[23499]), .B(p_input[13499]), .Z(n14450) );
  AND U21675 ( .A(p_input[3499]), .B(p_input[33499]), .Z(n14449) );
  AND U21676 ( .A(n14451), .B(n14452), .Z(o[3498]) );
  AND U21677 ( .A(p_input[23498]), .B(p_input[13498]), .Z(n14452) );
  AND U21678 ( .A(p_input[3498]), .B(p_input[33498]), .Z(n14451) );
  AND U21679 ( .A(n14453), .B(n14454), .Z(o[3497]) );
  AND U21680 ( .A(p_input[23497]), .B(p_input[13497]), .Z(n14454) );
  AND U21681 ( .A(p_input[3497]), .B(p_input[33497]), .Z(n14453) );
  AND U21682 ( .A(n14455), .B(n14456), .Z(o[3496]) );
  AND U21683 ( .A(p_input[23496]), .B(p_input[13496]), .Z(n14456) );
  AND U21684 ( .A(p_input[3496]), .B(p_input[33496]), .Z(n14455) );
  AND U21685 ( .A(n14457), .B(n14458), .Z(o[3495]) );
  AND U21686 ( .A(p_input[23495]), .B(p_input[13495]), .Z(n14458) );
  AND U21687 ( .A(p_input[3495]), .B(p_input[33495]), .Z(n14457) );
  AND U21688 ( .A(n14459), .B(n14460), .Z(o[3494]) );
  AND U21689 ( .A(p_input[23494]), .B(p_input[13494]), .Z(n14460) );
  AND U21690 ( .A(p_input[3494]), .B(p_input[33494]), .Z(n14459) );
  AND U21691 ( .A(n14461), .B(n14462), .Z(o[3493]) );
  AND U21692 ( .A(p_input[23493]), .B(p_input[13493]), .Z(n14462) );
  AND U21693 ( .A(p_input[3493]), .B(p_input[33493]), .Z(n14461) );
  AND U21694 ( .A(n14463), .B(n14464), .Z(o[3492]) );
  AND U21695 ( .A(p_input[23492]), .B(p_input[13492]), .Z(n14464) );
  AND U21696 ( .A(p_input[3492]), .B(p_input[33492]), .Z(n14463) );
  AND U21697 ( .A(n14465), .B(n14466), .Z(o[3491]) );
  AND U21698 ( .A(p_input[23491]), .B(p_input[13491]), .Z(n14466) );
  AND U21699 ( .A(p_input[3491]), .B(p_input[33491]), .Z(n14465) );
  AND U21700 ( .A(n14467), .B(n14468), .Z(o[3490]) );
  AND U21701 ( .A(p_input[23490]), .B(p_input[13490]), .Z(n14468) );
  AND U21702 ( .A(p_input[3490]), .B(p_input[33490]), .Z(n14467) );
  AND U21703 ( .A(n14469), .B(n14470), .Z(o[348]) );
  AND U21704 ( .A(p_input[20348]), .B(p_input[10348]), .Z(n14470) );
  AND U21705 ( .A(p_input[348]), .B(p_input[30348]), .Z(n14469) );
  AND U21706 ( .A(n14471), .B(n14472), .Z(o[3489]) );
  AND U21707 ( .A(p_input[23489]), .B(p_input[13489]), .Z(n14472) );
  AND U21708 ( .A(p_input[3489]), .B(p_input[33489]), .Z(n14471) );
  AND U21709 ( .A(n14473), .B(n14474), .Z(o[3488]) );
  AND U21710 ( .A(p_input[23488]), .B(p_input[13488]), .Z(n14474) );
  AND U21711 ( .A(p_input[3488]), .B(p_input[33488]), .Z(n14473) );
  AND U21712 ( .A(n14475), .B(n14476), .Z(o[3487]) );
  AND U21713 ( .A(p_input[23487]), .B(p_input[13487]), .Z(n14476) );
  AND U21714 ( .A(p_input[3487]), .B(p_input[33487]), .Z(n14475) );
  AND U21715 ( .A(n14477), .B(n14478), .Z(o[3486]) );
  AND U21716 ( .A(p_input[23486]), .B(p_input[13486]), .Z(n14478) );
  AND U21717 ( .A(p_input[3486]), .B(p_input[33486]), .Z(n14477) );
  AND U21718 ( .A(n14479), .B(n14480), .Z(o[3485]) );
  AND U21719 ( .A(p_input[23485]), .B(p_input[13485]), .Z(n14480) );
  AND U21720 ( .A(p_input[3485]), .B(p_input[33485]), .Z(n14479) );
  AND U21721 ( .A(n14481), .B(n14482), .Z(o[3484]) );
  AND U21722 ( .A(p_input[23484]), .B(p_input[13484]), .Z(n14482) );
  AND U21723 ( .A(p_input[3484]), .B(p_input[33484]), .Z(n14481) );
  AND U21724 ( .A(n14483), .B(n14484), .Z(o[3483]) );
  AND U21725 ( .A(p_input[23483]), .B(p_input[13483]), .Z(n14484) );
  AND U21726 ( .A(p_input[3483]), .B(p_input[33483]), .Z(n14483) );
  AND U21727 ( .A(n14485), .B(n14486), .Z(o[3482]) );
  AND U21728 ( .A(p_input[23482]), .B(p_input[13482]), .Z(n14486) );
  AND U21729 ( .A(p_input[3482]), .B(p_input[33482]), .Z(n14485) );
  AND U21730 ( .A(n14487), .B(n14488), .Z(o[3481]) );
  AND U21731 ( .A(p_input[23481]), .B(p_input[13481]), .Z(n14488) );
  AND U21732 ( .A(p_input[3481]), .B(p_input[33481]), .Z(n14487) );
  AND U21733 ( .A(n14489), .B(n14490), .Z(o[3480]) );
  AND U21734 ( .A(p_input[23480]), .B(p_input[13480]), .Z(n14490) );
  AND U21735 ( .A(p_input[3480]), .B(p_input[33480]), .Z(n14489) );
  AND U21736 ( .A(n14491), .B(n14492), .Z(o[347]) );
  AND U21737 ( .A(p_input[20347]), .B(p_input[10347]), .Z(n14492) );
  AND U21738 ( .A(p_input[347]), .B(p_input[30347]), .Z(n14491) );
  AND U21739 ( .A(n14493), .B(n14494), .Z(o[3479]) );
  AND U21740 ( .A(p_input[23479]), .B(p_input[13479]), .Z(n14494) );
  AND U21741 ( .A(p_input[3479]), .B(p_input[33479]), .Z(n14493) );
  AND U21742 ( .A(n14495), .B(n14496), .Z(o[3478]) );
  AND U21743 ( .A(p_input[23478]), .B(p_input[13478]), .Z(n14496) );
  AND U21744 ( .A(p_input[3478]), .B(p_input[33478]), .Z(n14495) );
  AND U21745 ( .A(n14497), .B(n14498), .Z(o[3477]) );
  AND U21746 ( .A(p_input[23477]), .B(p_input[13477]), .Z(n14498) );
  AND U21747 ( .A(p_input[3477]), .B(p_input[33477]), .Z(n14497) );
  AND U21748 ( .A(n14499), .B(n14500), .Z(o[3476]) );
  AND U21749 ( .A(p_input[23476]), .B(p_input[13476]), .Z(n14500) );
  AND U21750 ( .A(p_input[3476]), .B(p_input[33476]), .Z(n14499) );
  AND U21751 ( .A(n14501), .B(n14502), .Z(o[3475]) );
  AND U21752 ( .A(p_input[23475]), .B(p_input[13475]), .Z(n14502) );
  AND U21753 ( .A(p_input[3475]), .B(p_input[33475]), .Z(n14501) );
  AND U21754 ( .A(n14503), .B(n14504), .Z(o[3474]) );
  AND U21755 ( .A(p_input[23474]), .B(p_input[13474]), .Z(n14504) );
  AND U21756 ( .A(p_input[3474]), .B(p_input[33474]), .Z(n14503) );
  AND U21757 ( .A(n14505), .B(n14506), .Z(o[3473]) );
  AND U21758 ( .A(p_input[23473]), .B(p_input[13473]), .Z(n14506) );
  AND U21759 ( .A(p_input[3473]), .B(p_input[33473]), .Z(n14505) );
  AND U21760 ( .A(n14507), .B(n14508), .Z(o[3472]) );
  AND U21761 ( .A(p_input[23472]), .B(p_input[13472]), .Z(n14508) );
  AND U21762 ( .A(p_input[3472]), .B(p_input[33472]), .Z(n14507) );
  AND U21763 ( .A(n14509), .B(n14510), .Z(o[3471]) );
  AND U21764 ( .A(p_input[23471]), .B(p_input[13471]), .Z(n14510) );
  AND U21765 ( .A(p_input[3471]), .B(p_input[33471]), .Z(n14509) );
  AND U21766 ( .A(n14511), .B(n14512), .Z(o[3470]) );
  AND U21767 ( .A(p_input[23470]), .B(p_input[13470]), .Z(n14512) );
  AND U21768 ( .A(p_input[3470]), .B(p_input[33470]), .Z(n14511) );
  AND U21769 ( .A(n14513), .B(n14514), .Z(o[346]) );
  AND U21770 ( .A(p_input[20346]), .B(p_input[10346]), .Z(n14514) );
  AND U21771 ( .A(p_input[346]), .B(p_input[30346]), .Z(n14513) );
  AND U21772 ( .A(n14515), .B(n14516), .Z(o[3469]) );
  AND U21773 ( .A(p_input[23469]), .B(p_input[13469]), .Z(n14516) );
  AND U21774 ( .A(p_input[3469]), .B(p_input[33469]), .Z(n14515) );
  AND U21775 ( .A(n14517), .B(n14518), .Z(o[3468]) );
  AND U21776 ( .A(p_input[23468]), .B(p_input[13468]), .Z(n14518) );
  AND U21777 ( .A(p_input[3468]), .B(p_input[33468]), .Z(n14517) );
  AND U21778 ( .A(n14519), .B(n14520), .Z(o[3467]) );
  AND U21779 ( .A(p_input[23467]), .B(p_input[13467]), .Z(n14520) );
  AND U21780 ( .A(p_input[3467]), .B(p_input[33467]), .Z(n14519) );
  AND U21781 ( .A(n14521), .B(n14522), .Z(o[3466]) );
  AND U21782 ( .A(p_input[23466]), .B(p_input[13466]), .Z(n14522) );
  AND U21783 ( .A(p_input[3466]), .B(p_input[33466]), .Z(n14521) );
  AND U21784 ( .A(n14523), .B(n14524), .Z(o[3465]) );
  AND U21785 ( .A(p_input[23465]), .B(p_input[13465]), .Z(n14524) );
  AND U21786 ( .A(p_input[3465]), .B(p_input[33465]), .Z(n14523) );
  AND U21787 ( .A(n14525), .B(n14526), .Z(o[3464]) );
  AND U21788 ( .A(p_input[23464]), .B(p_input[13464]), .Z(n14526) );
  AND U21789 ( .A(p_input[3464]), .B(p_input[33464]), .Z(n14525) );
  AND U21790 ( .A(n14527), .B(n14528), .Z(o[3463]) );
  AND U21791 ( .A(p_input[23463]), .B(p_input[13463]), .Z(n14528) );
  AND U21792 ( .A(p_input[3463]), .B(p_input[33463]), .Z(n14527) );
  AND U21793 ( .A(n14529), .B(n14530), .Z(o[3462]) );
  AND U21794 ( .A(p_input[23462]), .B(p_input[13462]), .Z(n14530) );
  AND U21795 ( .A(p_input[3462]), .B(p_input[33462]), .Z(n14529) );
  AND U21796 ( .A(n14531), .B(n14532), .Z(o[3461]) );
  AND U21797 ( .A(p_input[23461]), .B(p_input[13461]), .Z(n14532) );
  AND U21798 ( .A(p_input[3461]), .B(p_input[33461]), .Z(n14531) );
  AND U21799 ( .A(n14533), .B(n14534), .Z(o[3460]) );
  AND U21800 ( .A(p_input[23460]), .B(p_input[13460]), .Z(n14534) );
  AND U21801 ( .A(p_input[3460]), .B(p_input[33460]), .Z(n14533) );
  AND U21802 ( .A(n14535), .B(n14536), .Z(o[345]) );
  AND U21803 ( .A(p_input[20345]), .B(p_input[10345]), .Z(n14536) );
  AND U21804 ( .A(p_input[345]), .B(p_input[30345]), .Z(n14535) );
  AND U21805 ( .A(n14537), .B(n14538), .Z(o[3459]) );
  AND U21806 ( .A(p_input[23459]), .B(p_input[13459]), .Z(n14538) );
  AND U21807 ( .A(p_input[3459]), .B(p_input[33459]), .Z(n14537) );
  AND U21808 ( .A(n14539), .B(n14540), .Z(o[3458]) );
  AND U21809 ( .A(p_input[23458]), .B(p_input[13458]), .Z(n14540) );
  AND U21810 ( .A(p_input[3458]), .B(p_input[33458]), .Z(n14539) );
  AND U21811 ( .A(n14541), .B(n14542), .Z(o[3457]) );
  AND U21812 ( .A(p_input[23457]), .B(p_input[13457]), .Z(n14542) );
  AND U21813 ( .A(p_input[3457]), .B(p_input[33457]), .Z(n14541) );
  AND U21814 ( .A(n14543), .B(n14544), .Z(o[3456]) );
  AND U21815 ( .A(p_input[23456]), .B(p_input[13456]), .Z(n14544) );
  AND U21816 ( .A(p_input[3456]), .B(p_input[33456]), .Z(n14543) );
  AND U21817 ( .A(n14545), .B(n14546), .Z(o[3455]) );
  AND U21818 ( .A(p_input[23455]), .B(p_input[13455]), .Z(n14546) );
  AND U21819 ( .A(p_input[3455]), .B(p_input[33455]), .Z(n14545) );
  AND U21820 ( .A(n14547), .B(n14548), .Z(o[3454]) );
  AND U21821 ( .A(p_input[23454]), .B(p_input[13454]), .Z(n14548) );
  AND U21822 ( .A(p_input[3454]), .B(p_input[33454]), .Z(n14547) );
  AND U21823 ( .A(n14549), .B(n14550), .Z(o[3453]) );
  AND U21824 ( .A(p_input[23453]), .B(p_input[13453]), .Z(n14550) );
  AND U21825 ( .A(p_input[3453]), .B(p_input[33453]), .Z(n14549) );
  AND U21826 ( .A(n14551), .B(n14552), .Z(o[3452]) );
  AND U21827 ( .A(p_input[23452]), .B(p_input[13452]), .Z(n14552) );
  AND U21828 ( .A(p_input[3452]), .B(p_input[33452]), .Z(n14551) );
  AND U21829 ( .A(n14553), .B(n14554), .Z(o[3451]) );
  AND U21830 ( .A(p_input[23451]), .B(p_input[13451]), .Z(n14554) );
  AND U21831 ( .A(p_input[3451]), .B(p_input[33451]), .Z(n14553) );
  AND U21832 ( .A(n14555), .B(n14556), .Z(o[3450]) );
  AND U21833 ( .A(p_input[23450]), .B(p_input[13450]), .Z(n14556) );
  AND U21834 ( .A(p_input[3450]), .B(p_input[33450]), .Z(n14555) );
  AND U21835 ( .A(n14557), .B(n14558), .Z(o[344]) );
  AND U21836 ( .A(p_input[20344]), .B(p_input[10344]), .Z(n14558) );
  AND U21837 ( .A(p_input[344]), .B(p_input[30344]), .Z(n14557) );
  AND U21838 ( .A(n14559), .B(n14560), .Z(o[3449]) );
  AND U21839 ( .A(p_input[23449]), .B(p_input[13449]), .Z(n14560) );
  AND U21840 ( .A(p_input[3449]), .B(p_input[33449]), .Z(n14559) );
  AND U21841 ( .A(n14561), .B(n14562), .Z(o[3448]) );
  AND U21842 ( .A(p_input[23448]), .B(p_input[13448]), .Z(n14562) );
  AND U21843 ( .A(p_input[3448]), .B(p_input[33448]), .Z(n14561) );
  AND U21844 ( .A(n14563), .B(n14564), .Z(o[3447]) );
  AND U21845 ( .A(p_input[23447]), .B(p_input[13447]), .Z(n14564) );
  AND U21846 ( .A(p_input[3447]), .B(p_input[33447]), .Z(n14563) );
  AND U21847 ( .A(n14565), .B(n14566), .Z(o[3446]) );
  AND U21848 ( .A(p_input[23446]), .B(p_input[13446]), .Z(n14566) );
  AND U21849 ( .A(p_input[3446]), .B(p_input[33446]), .Z(n14565) );
  AND U21850 ( .A(n14567), .B(n14568), .Z(o[3445]) );
  AND U21851 ( .A(p_input[23445]), .B(p_input[13445]), .Z(n14568) );
  AND U21852 ( .A(p_input[3445]), .B(p_input[33445]), .Z(n14567) );
  AND U21853 ( .A(n14569), .B(n14570), .Z(o[3444]) );
  AND U21854 ( .A(p_input[23444]), .B(p_input[13444]), .Z(n14570) );
  AND U21855 ( .A(p_input[3444]), .B(p_input[33444]), .Z(n14569) );
  AND U21856 ( .A(n14571), .B(n14572), .Z(o[3443]) );
  AND U21857 ( .A(p_input[23443]), .B(p_input[13443]), .Z(n14572) );
  AND U21858 ( .A(p_input[3443]), .B(p_input[33443]), .Z(n14571) );
  AND U21859 ( .A(n14573), .B(n14574), .Z(o[3442]) );
  AND U21860 ( .A(p_input[23442]), .B(p_input[13442]), .Z(n14574) );
  AND U21861 ( .A(p_input[3442]), .B(p_input[33442]), .Z(n14573) );
  AND U21862 ( .A(n14575), .B(n14576), .Z(o[3441]) );
  AND U21863 ( .A(p_input[23441]), .B(p_input[13441]), .Z(n14576) );
  AND U21864 ( .A(p_input[3441]), .B(p_input[33441]), .Z(n14575) );
  AND U21865 ( .A(n14577), .B(n14578), .Z(o[3440]) );
  AND U21866 ( .A(p_input[23440]), .B(p_input[13440]), .Z(n14578) );
  AND U21867 ( .A(p_input[3440]), .B(p_input[33440]), .Z(n14577) );
  AND U21868 ( .A(n14579), .B(n14580), .Z(o[343]) );
  AND U21869 ( .A(p_input[20343]), .B(p_input[10343]), .Z(n14580) );
  AND U21870 ( .A(p_input[343]), .B(p_input[30343]), .Z(n14579) );
  AND U21871 ( .A(n14581), .B(n14582), .Z(o[3439]) );
  AND U21872 ( .A(p_input[23439]), .B(p_input[13439]), .Z(n14582) );
  AND U21873 ( .A(p_input[3439]), .B(p_input[33439]), .Z(n14581) );
  AND U21874 ( .A(n14583), .B(n14584), .Z(o[3438]) );
  AND U21875 ( .A(p_input[23438]), .B(p_input[13438]), .Z(n14584) );
  AND U21876 ( .A(p_input[3438]), .B(p_input[33438]), .Z(n14583) );
  AND U21877 ( .A(n14585), .B(n14586), .Z(o[3437]) );
  AND U21878 ( .A(p_input[23437]), .B(p_input[13437]), .Z(n14586) );
  AND U21879 ( .A(p_input[3437]), .B(p_input[33437]), .Z(n14585) );
  AND U21880 ( .A(n14587), .B(n14588), .Z(o[3436]) );
  AND U21881 ( .A(p_input[23436]), .B(p_input[13436]), .Z(n14588) );
  AND U21882 ( .A(p_input[3436]), .B(p_input[33436]), .Z(n14587) );
  AND U21883 ( .A(n14589), .B(n14590), .Z(o[3435]) );
  AND U21884 ( .A(p_input[23435]), .B(p_input[13435]), .Z(n14590) );
  AND U21885 ( .A(p_input[3435]), .B(p_input[33435]), .Z(n14589) );
  AND U21886 ( .A(n14591), .B(n14592), .Z(o[3434]) );
  AND U21887 ( .A(p_input[23434]), .B(p_input[13434]), .Z(n14592) );
  AND U21888 ( .A(p_input[3434]), .B(p_input[33434]), .Z(n14591) );
  AND U21889 ( .A(n14593), .B(n14594), .Z(o[3433]) );
  AND U21890 ( .A(p_input[23433]), .B(p_input[13433]), .Z(n14594) );
  AND U21891 ( .A(p_input[3433]), .B(p_input[33433]), .Z(n14593) );
  AND U21892 ( .A(n14595), .B(n14596), .Z(o[3432]) );
  AND U21893 ( .A(p_input[23432]), .B(p_input[13432]), .Z(n14596) );
  AND U21894 ( .A(p_input[3432]), .B(p_input[33432]), .Z(n14595) );
  AND U21895 ( .A(n14597), .B(n14598), .Z(o[3431]) );
  AND U21896 ( .A(p_input[23431]), .B(p_input[13431]), .Z(n14598) );
  AND U21897 ( .A(p_input[3431]), .B(p_input[33431]), .Z(n14597) );
  AND U21898 ( .A(n14599), .B(n14600), .Z(o[3430]) );
  AND U21899 ( .A(p_input[23430]), .B(p_input[13430]), .Z(n14600) );
  AND U21900 ( .A(p_input[3430]), .B(p_input[33430]), .Z(n14599) );
  AND U21901 ( .A(n14601), .B(n14602), .Z(o[342]) );
  AND U21902 ( .A(p_input[20342]), .B(p_input[10342]), .Z(n14602) );
  AND U21903 ( .A(p_input[342]), .B(p_input[30342]), .Z(n14601) );
  AND U21904 ( .A(n14603), .B(n14604), .Z(o[3429]) );
  AND U21905 ( .A(p_input[23429]), .B(p_input[13429]), .Z(n14604) );
  AND U21906 ( .A(p_input[3429]), .B(p_input[33429]), .Z(n14603) );
  AND U21907 ( .A(n14605), .B(n14606), .Z(o[3428]) );
  AND U21908 ( .A(p_input[23428]), .B(p_input[13428]), .Z(n14606) );
  AND U21909 ( .A(p_input[3428]), .B(p_input[33428]), .Z(n14605) );
  AND U21910 ( .A(n14607), .B(n14608), .Z(o[3427]) );
  AND U21911 ( .A(p_input[23427]), .B(p_input[13427]), .Z(n14608) );
  AND U21912 ( .A(p_input[3427]), .B(p_input[33427]), .Z(n14607) );
  AND U21913 ( .A(n14609), .B(n14610), .Z(o[3426]) );
  AND U21914 ( .A(p_input[23426]), .B(p_input[13426]), .Z(n14610) );
  AND U21915 ( .A(p_input[3426]), .B(p_input[33426]), .Z(n14609) );
  AND U21916 ( .A(n14611), .B(n14612), .Z(o[3425]) );
  AND U21917 ( .A(p_input[23425]), .B(p_input[13425]), .Z(n14612) );
  AND U21918 ( .A(p_input[3425]), .B(p_input[33425]), .Z(n14611) );
  AND U21919 ( .A(n14613), .B(n14614), .Z(o[3424]) );
  AND U21920 ( .A(p_input[23424]), .B(p_input[13424]), .Z(n14614) );
  AND U21921 ( .A(p_input[3424]), .B(p_input[33424]), .Z(n14613) );
  AND U21922 ( .A(n14615), .B(n14616), .Z(o[3423]) );
  AND U21923 ( .A(p_input[23423]), .B(p_input[13423]), .Z(n14616) );
  AND U21924 ( .A(p_input[3423]), .B(p_input[33423]), .Z(n14615) );
  AND U21925 ( .A(n14617), .B(n14618), .Z(o[3422]) );
  AND U21926 ( .A(p_input[23422]), .B(p_input[13422]), .Z(n14618) );
  AND U21927 ( .A(p_input[3422]), .B(p_input[33422]), .Z(n14617) );
  AND U21928 ( .A(n14619), .B(n14620), .Z(o[3421]) );
  AND U21929 ( .A(p_input[23421]), .B(p_input[13421]), .Z(n14620) );
  AND U21930 ( .A(p_input[3421]), .B(p_input[33421]), .Z(n14619) );
  AND U21931 ( .A(n14621), .B(n14622), .Z(o[3420]) );
  AND U21932 ( .A(p_input[23420]), .B(p_input[13420]), .Z(n14622) );
  AND U21933 ( .A(p_input[3420]), .B(p_input[33420]), .Z(n14621) );
  AND U21934 ( .A(n14623), .B(n14624), .Z(o[341]) );
  AND U21935 ( .A(p_input[20341]), .B(p_input[10341]), .Z(n14624) );
  AND U21936 ( .A(p_input[341]), .B(p_input[30341]), .Z(n14623) );
  AND U21937 ( .A(n14625), .B(n14626), .Z(o[3419]) );
  AND U21938 ( .A(p_input[23419]), .B(p_input[13419]), .Z(n14626) );
  AND U21939 ( .A(p_input[3419]), .B(p_input[33419]), .Z(n14625) );
  AND U21940 ( .A(n14627), .B(n14628), .Z(o[3418]) );
  AND U21941 ( .A(p_input[23418]), .B(p_input[13418]), .Z(n14628) );
  AND U21942 ( .A(p_input[3418]), .B(p_input[33418]), .Z(n14627) );
  AND U21943 ( .A(n14629), .B(n14630), .Z(o[3417]) );
  AND U21944 ( .A(p_input[23417]), .B(p_input[13417]), .Z(n14630) );
  AND U21945 ( .A(p_input[3417]), .B(p_input[33417]), .Z(n14629) );
  AND U21946 ( .A(n14631), .B(n14632), .Z(o[3416]) );
  AND U21947 ( .A(p_input[23416]), .B(p_input[13416]), .Z(n14632) );
  AND U21948 ( .A(p_input[3416]), .B(p_input[33416]), .Z(n14631) );
  AND U21949 ( .A(n14633), .B(n14634), .Z(o[3415]) );
  AND U21950 ( .A(p_input[23415]), .B(p_input[13415]), .Z(n14634) );
  AND U21951 ( .A(p_input[3415]), .B(p_input[33415]), .Z(n14633) );
  AND U21952 ( .A(n14635), .B(n14636), .Z(o[3414]) );
  AND U21953 ( .A(p_input[23414]), .B(p_input[13414]), .Z(n14636) );
  AND U21954 ( .A(p_input[3414]), .B(p_input[33414]), .Z(n14635) );
  AND U21955 ( .A(n14637), .B(n14638), .Z(o[3413]) );
  AND U21956 ( .A(p_input[23413]), .B(p_input[13413]), .Z(n14638) );
  AND U21957 ( .A(p_input[3413]), .B(p_input[33413]), .Z(n14637) );
  AND U21958 ( .A(n14639), .B(n14640), .Z(o[3412]) );
  AND U21959 ( .A(p_input[23412]), .B(p_input[13412]), .Z(n14640) );
  AND U21960 ( .A(p_input[3412]), .B(p_input[33412]), .Z(n14639) );
  AND U21961 ( .A(n14641), .B(n14642), .Z(o[3411]) );
  AND U21962 ( .A(p_input[23411]), .B(p_input[13411]), .Z(n14642) );
  AND U21963 ( .A(p_input[3411]), .B(p_input[33411]), .Z(n14641) );
  AND U21964 ( .A(n14643), .B(n14644), .Z(o[3410]) );
  AND U21965 ( .A(p_input[23410]), .B(p_input[13410]), .Z(n14644) );
  AND U21966 ( .A(p_input[3410]), .B(p_input[33410]), .Z(n14643) );
  AND U21967 ( .A(n14645), .B(n14646), .Z(o[340]) );
  AND U21968 ( .A(p_input[20340]), .B(p_input[10340]), .Z(n14646) );
  AND U21969 ( .A(p_input[340]), .B(p_input[30340]), .Z(n14645) );
  AND U21970 ( .A(n14647), .B(n14648), .Z(o[3409]) );
  AND U21971 ( .A(p_input[23409]), .B(p_input[13409]), .Z(n14648) );
  AND U21972 ( .A(p_input[3409]), .B(p_input[33409]), .Z(n14647) );
  AND U21973 ( .A(n14649), .B(n14650), .Z(o[3408]) );
  AND U21974 ( .A(p_input[23408]), .B(p_input[13408]), .Z(n14650) );
  AND U21975 ( .A(p_input[3408]), .B(p_input[33408]), .Z(n14649) );
  AND U21976 ( .A(n14651), .B(n14652), .Z(o[3407]) );
  AND U21977 ( .A(p_input[23407]), .B(p_input[13407]), .Z(n14652) );
  AND U21978 ( .A(p_input[3407]), .B(p_input[33407]), .Z(n14651) );
  AND U21979 ( .A(n14653), .B(n14654), .Z(o[3406]) );
  AND U21980 ( .A(p_input[23406]), .B(p_input[13406]), .Z(n14654) );
  AND U21981 ( .A(p_input[3406]), .B(p_input[33406]), .Z(n14653) );
  AND U21982 ( .A(n14655), .B(n14656), .Z(o[3405]) );
  AND U21983 ( .A(p_input[23405]), .B(p_input[13405]), .Z(n14656) );
  AND U21984 ( .A(p_input[3405]), .B(p_input[33405]), .Z(n14655) );
  AND U21985 ( .A(n14657), .B(n14658), .Z(o[3404]) );
  AND U21986 ( .A(p_input[23404]), .B(p_input[13404]), .Z(n14658) );
  AND U21987 ( .A(p_input[3404]), .B(p_input[33404]), .Z(n14657) );
  AND U21988 ( .A(n14659), .B(n14660), .Z(o[3403]) );
  AND U21989 ( .A(p_input[23403]), .B(p_input[13403]), .Z(n14660) );
  AND U21990 ( .A(p_input[3403]), .B(p_input[33403]), .Z(n14659) );
  AND U21991 ( .A(n14661), .B(n14662), .Z(o[3402]) );
  AND U21992 ( .A(p_input[23402]), .B(p_input[13402]), .Z(n14662) );
  AND U21993 ( .A(p_input[3402]), .B(p_input[33402]), .Z(n14661) );
  AND U21994 ( .A(n14663), .B(n14664), .Z(o[3401]) );
  AND U21995 ( .A(p_input[23401]), .B(p_input[13401]), .Z(n14664) );
  AND U21996 ( .A(p_input[3401]), .B(p_input[33401]), .Z(n14663) );
  AND U21997 ( .A(n14665), .B(n14666), .Z(o[3400]) );
  AND U21998 ( .A(p_input[23400]), .B(p_input[13400]), .Z(n14666) );
  AND U21999 ( .A(p_input[3400]), .B(p_input[33400]), .Z(n14665) );
  AND U22000 ( .A(n14667), .B(n14668), .Z(o[33]) );
  AND U22001 ( .A(p_input[20033]), .B(p_input[10033]), .Z(n14668) );
  AND U22002 ( .A(p_input[33]), .B(p_input[30033]), .Z(n14667) );
  AND U22003 ( .A(n14669), .B(n14670), .Z(o[339]) );
  AND U22004 ( .A(p_input[20339]), .B(p_input[10339]), .Z(n14670) );
  AND U22005 ( .A(p_input[339]), .B(p_input[30339]), .Z(n14669) );
  AND U22006 ( .A(n14671), .B(n14672), .Z(o[3399]) );
  AND U22007 ( .A(p_input[23399]), .B(p_input[13399]), .Z(n14672) );
  AND U22008 ( .A(p_input[3399]), .B(p_input[33399]), .Z(n14671) );
  AND U22009 ( .A(n14673), .B(n14674), .Z(o[3398]) );
  AND U22010 ( .A(p_input[23398]), .B(p_input[13398]), .Z(n14674) );
  AND U22011 ( .A(p_input[3398]), .B(p_input[33398]), .Z(n14673) );
  AND U22012 ( .A(n14675), .B(n14676), .Z(o[3397]) );
  AND U22013 ( .A(p_input[23397]), .B(p_input[13397]), .Z(n14676) );
  AND U22014 ( .A(p_input[3397]), .B(p_input[33397]), .Z(n14675) );
  AND U22015 ( .A(n14677), .B(n14678), .Z(o[3396]) );
  AND U22016 ( .A(p_input[23396]), .B(p_input[13396]), .Z(n14678) );
  AND U22017 ( .A(p_input[3396]), .B(p_input[33396]), .Z(n14677) );
  AND U22018 ( .A(n14679), .B(n14680), .Z(o[3395]) );
  AND U22019 ( .A(p_input[23395]), .B(p_input[13395]), .Z(n14680) );
  AND U22020 ( .A(p_input[3395]), .B(p_input[33395]), .Z(n14679) );
  AND U22021 ( .A(n14681), .B(n14682), .Z(o[3394]) );
  AND U22022 ( .A(p_input[23394]), .B(p_input[13394]), .Z(n14682) );
  AND U22023 ( .A(p_input[3394]), .B(p_input[33394]), .Z(n14681) );
  AND U22024 ( .A(n14683), .B(n14684), .Z(o[3393]) );
  AND U22025 ( .A(p_input[23393]), .B(p_input[13393]), .Z(n14684) );
  AND U22026 ( .A(p_input[3393]), .B(p_input[33393]), .Z(n14683) );
  AND U22027 ( .A(n14685), .B(n14686), .Z(o[3392]) );
  AND U22028 ( .A(p_input[23392]), .B(p_input[13392]), .Z(n14686) );
  AND U22029 ( .A(p_input[3392]), .B(p_input[33392]), .Z(n14685) );
  AND U22030 ( .A(n14687), .B(n14688), .Z(o[3391]) );
  AND U22031 ( .A(p_input[23391]), .B(p_input[13391]), .Z(n14688) );
  AND U22032 ( .A(p_input[3391]), .B(p_input[33391]), .Z(n14687) );
  AND U22033 ( .A(n14689), .B(n14690), .Z(o[3390]) );
  AND U22034 ( .A(p_input[23390]), .B(p_input[13390]), .Z(n14690) );
  AND U22035 ( .A(p_input[3390]), .B(p_input[33390]), .Z(n14689) );
  AND U22036 ( .A(n14691), .B(n14692), .Z(o[338]) );
  AND U22037 ( .A(p_input[20338]), .B(p_input[10338]), .Z(n14692) );
  AND U22038 ( .A(p_input[338]), .B(p_input[30338]), .Z(n14691) );
  AND U22039 ( .A(n14693), .B(n14694), .Z(o[3389]) );
  AND U22040 ( .A(p_input[23389]), .B(p_input[13389]), .Z(n14694) );
  AND U22041 ( .A(p_input[3389]), .B(p_input[33389]), .Z(n14693) );
  AND U22042 ( .A(n14695), .B(n14696), .Z(o[3388]) );
  AND U22043 ( .A(p_input[23388]), .B(p_input[13388]), .Z(n14696) );
  AND U22044 ( .A(p_input[3388]), .B(p_input[33388]), .Z(n14695) );
  AND U22045 ( .A(n14697), .B(n14698), .Z(o[3387]) );
  AND U22046 ( .A(p_input[23387]), .B(p_input[13387]), .Z(n14698) );
  AND U22047 ( .A(p_input[3387]), .B(p_input[33387]), .Z(n14697) );
  AND U22048 ( .A(n14699), .B(n14700), .Z(o[3386]) );
  AND U22049 ( .A(p_input[23386]), .B(p_input[13386]), .Z(n14700) );
  AND U22050 ( .A(p_input[3386]), .B(p_input[33386]), .Z(n14699) );
  AND U22051 ( .A(n14701), .B(n14702), .Z(o[3385]) );
  AND U22052 ( .A(p_input[23385]), .B(p_input[13385]), .Z(n14702) );
  AND U22053 ( .A(p_input[3385]), .B(p_input[33385]), .Z(n14701) );
  AND U22054 ( .A(n14703), .B(n14704), .Z(o[3384]) );
  AND U22055 ( .A(p_input[23384]), .B(p_input[13384]), .Z(n14704) );
  AND U22056 ( .A(p_input[3384]), .B(p_input[33384]), .Z(n14703) );
  AND U22057 ( .A(n14705), .B(n14706), .Z(o[3383]) );
  AND U22058 ( .A(p_input[23383]), .B(p_input[13383]), .Z(n14706) );
  AND U22059 ( .A(p_input[3383]), .B(p_input[33383]), .Z(n14705) );
  AND U22060 ( .A(n14707), .B(n14708), .Z(o[3382]) );
  AND U22061 ( .A(p_input[23382]), .B(p_input[13382]), .Z(n14708) );
  AND U22062 ( .A(p_input[3382]), .B(p_input[33382]), .Z(n14707) );
  AND U22063 ( .A(n14709), .B(n14710), .Z(o[3381]) );
  AND U22064 ( .A(p_input[23381]), .B(p_input[13381]), .Z(n14710) );
  AND U22065 ( .A(p_input[3381]), .B(p_input[33381]), .Z(n14709) );
  AND U22066 ( .A(n14711), .B(n14712), .Z(o[3380]) );
  AND U22067 ( .A(p_input[23380]), .B(p_input[13380]), .Z(n14712) );
  AND U22068 ( .A(p_input[3380]), .B(p_input[33380]), .Z(n14711) );
  AND U22069 ( .A(n14713), .B(n14714), .Z(o[337]) );
  AND U22070 ( .A(p_input[20337]), .B(p_input[10337]), .Z(n14714) );
  AND U22071 ( .A(p_input[337]), .B(p_input[30337]), .Z(n14713) );
  AND U22072 ( .A(n14715), .B(n14716), .Z(o[3379]) );
  AND U22073 ( .A(p_input[23379]), .B(p_input[13379]), .Z(n14716) );
  AND U22074 ( .A(p_input[3379]), .B(p_input[33379]), .Z(n14715) );
  AND U22075 ( .A(n14717), .B(n14718), .Z(o[3378]) );
  AND U22076 ( .A(p_input[23378]), .B(p_input[13378]), .Z(n14718) );
  AND U22077 ( .A(p_input[3378]), .B(p_input[33378]), .Z(n14717) );
  AND U22078 ( .A(n14719), .B(n14720), .Z(o[3377]) );
  AND U22079 ( .A(p_input[23377]), .B(p_input[13377]), .Z(n14720) );
  AND U22080 ( .A(p_input[3377]), .B(p_input[33377]), .Z(n14719) );
  AND U22081 ( .A(n14721), .B(n14722), .Z(o[3376]) );
  AND U22082 ( .A(p_input[23376]), .B(p_input[13376]), .Z(n14722) );
  AND U22083 ( .A(p_input[3376]), .B(p_input[33376]), .Z(n14721) );
  AND U22084 ( .A(n14723), .B(n14724), .Z(o[3375]) );
  AND U22085 ( .A(p_input[23375]), .B(p_input[13375]), .Z(n14724) );
  AND U22086 ( .A(p_input[3375]), .B(p_input[33375]), .Z(n14723) );
  AND U22087 ( .A(n14725), .B(n14726), .Z(o[3374]) );
  AND U22088 ( .A(p_input[23374]), .B(p_input[13374]), .Z(n14726) );
  AND U22089 ( .A(p_input[3374]), .B(p_input[33374]), .Z(n14725) );
  AND U22090 ( .A(n14727), .B(n14728), .Z(o[3373]) );
  AND U22091 ( .A(p_input[23373]), .B(p_input[13373]), .Z(n14728) );
  AND U22092 ( .A(p_input[3373]), .B(p_input[33373]), .Z(n14727) );
  AND U22093 ( .A(n14729), .B(n14730), .Z(o[3372]) );
  AND U22094 ( .A(p_input[23372]), .B(p_input[13372]), .Z(n14730) );
  AND U22095 ( .A(p_input[3372]), .B(p_input[33372]), .Z(n14729) );
  AND U22096 ( .A(n14731), .B(n14732), .Z(o[3371]) );
  AND U22097 ( .A(p_input[23371]), .B(p_input[13371]), .Z(n14732) );
  AND U22098 ( .A(p_input[3371]), .B(p_input[33371]), .Z(n14731) );
  AND U22099 ( .A(n14733), .B(n14734), .Z(o[3370]) );
  AND U22100 ( .A(p_input[23370]), .B(p_input[13370]), .Z(n14734) );
  AND U22101 ( .A(p_input[3370]), .B(p_input[33370]), .Z(n14733) );
  AND U22102 ( .A(n14735), .B(n14736), .Z(o[336]) );
  AND U22103 ( .A(p_input[20336]), .B(p_input[10336]), .Z(n14736) );
  AND U22104 ( .A(p_input[336]), .B(p_input[30336]), .Z(n14735) );
  AND U22105 ( .A(n14737), .B(n14738), .Z(o[3369]) );
  AND U22106 ( .A(p_input[23369]), .B(p_input[13369]), .Z(n14738) );
  AND U22107 ( .A(p_input[3369]), .B(p_input[33369]), .Z(n14737) );
  AND U22108 ( .A(n14739), .B(n14740), .Z(o[3368]) );
  AND U22109 ( .A(p_input[23368]), .B(p_input[13368]), .Z(n14740) );
  AND U22110 ( .A(p_input[3368]), .B(p_input[33368]), .Z(n14739) );
  AND U22111 ( .A(n14741), .B(n14742), .Z(o[3367]) );
  AND U22112 ( .A(p_input[23367]), .B(p_input[13367]), .Z(n14742) );
  AND U22113 ( .A(p_input[3367]), .B(p_input[33367]), .Z(n14741) );
  AND U22114 ( .A(n14743), .B(n14744), .Z(o[3366]) );
  AND U22115 ( .A(p_input[23366]), .B(p_input[13366]), .Z(n14744) );
  AND U22116 ( .A(p_input[3366]), .B(p_input[33366]), .Z(n14743) );
  AND U22117 ( .A(n14745), .B(n14746), .Z(o[3365]) );
  AND U22118 ( .A(p_input[23365]), .B(p_input[13365]), .Z(n14746) );
  AND U22119 ( .A(p_input[3365]), .B(p_input[33365]), .Z(n14745) );
  AND U22120 ( .A(n14747), .B(n14748), .Z(o[3364]) );
  AND U22121 ( .A(p_input[23364]), .B(p_input[13364]), .Z(n14748) );
  AND U22122 ( .A(p_input[3364]), .B(p_input[33364]), .Z(n14747) );
  AND U22123 ( .A(n14749), .B(n14750), .Z(o[3363]) );
  AND U22124 ( .A(p_input[23363]), .B(p_input[13363]), .Z(n14750) );
  AND U22125 ( .A(p_input[3363]), .B(p_input[33363]), .Z(n14749) );
  AND U22126 ( .A(n14751), .B(n14752), .Z(o[3362]) );
  AND U22127 ( .A(p_input[23362]), .B(p_input[13362]), .Z(n14752) );
  AND U22128 ( .A(p_input[3362]), .B(p_input[33362]), .Z(n14751) );
  AND U22129 ( .A(n14753), .B(n14754), .Z(o[3361]) );
  AND U22130 ( .A(p_input[23361]), .B(p_input[13361]), .Z(n14754) );
  AND U22131 ( .A(p_input[3361]), .B(p_input[33361]), .Z(n14753) );
  AND U22132 ( .A(n14755), .B(n14756), .Z(o[3360]) );
  AND U22133 ( .A(p_input[23360]), .B(p_input[13360]), .Z(n14756) );
  AND U22134 ( .A(p_input[3360]), .B(p_input[33360]), .Z(n14755) );
  AND U22135 ( .A(n14757), .B(n14758), .Z(o[335]) );
  AND U22136 ( .A(p_input[20335]), .B(p_input[10335]), .Z(n14758) );
  AND U22137 ( .A(p_input[335]), .B(p_input[30335]), .Z(n14757) );
  AND U22138 ( .A(n14759), .B(n14760), .Z(o[3359]) );
  AND U22139 ( .A(p_input[23359]), .B(p_input[13359]), .Z(n14760) );
  AND U22140 ( .A(p_input[3359]), .B(p_input[33359]), .Z(n14759) );
  AND U22141 ( .A(n14761), .B(n14762), .Z(o[3358]) );
  AND U22142 ( .A(p_input[23358]), .B(p_input[13358]), .Z(n14762) );
  AND U22143 ( .A(p_input[3358]), .B(p_input[33358]), .Z(n14761) );
  AND U22144 ( .A(n14763), .B(n14764), .Z(o[3357]) );
  AND U22145 ( .A(p_input[23357]), .B(p_input[13357]), .Z(n14764) );
  AND U22146 ( .A(p_input[3357]), .B(p_input[33357]), .Z(n14763) );
  AND U22147 ( .A(n14765), .B(n14766), .Z(o[3356]) );
  AND U22148 ( .A(p_input[23356]), .B(p_input[13356]), .Z(n14766) );
  AND U22149 ( .A(p_input[3356]), .B(p_input[33356]), .Z(n14765) );
  AND U22150 ( .A(n14767), .B(n14768), .Z(o[3355]) );
  AND U22151 ( .A(p_input[23355]), .B(p_input[13355]), .Z(n14768) );
  AND U22152 ( .A(p_input[3355]), .B(p_input[33355]), .Z(n14767) );
  AND U22153 ( .A(n14769), .B(n14770), .Z(o[3354]) );
  AND U22154 ( .A(p_input[23354]), .B(p_input[13354]), .Z(n14770) );
  AND U22155 ( .A(p_input[3354]), .B(p_input[33354]), .Z(n14769) );
  AND U22156 ( .A(n14771), .B(n14772), .Z(o[3353]) );
  AND U22157 ( .A(p_input[23353]), .B(p_input[13353]), .Z(n14772) );
  AND U22158 ( .A(p_input[3353]), .B(p_input[33353]), .Z(n14771) );
  AND U22159 ( .A(n14773), .B(n14774), .Z(o[3352]) );
  AND U22160 ( .A(p_input[23352]), .B(p_input[13352]), .Z(n14774) );
  AND U22161 ( .A(p_input[3352]), .B(p_input[33352]), .Z(n14773) );
  AND U22162 ( .A(n14775), .B(n14776), .Z(o[3351]) );
  AND U22163 ( .A(p_input[23351]), .B(p_input[13351]), .Z(n14776) );
  AND U22164 ( .A(p_input[3351]), .B(p_input[33351]), .Z(n14775) );
  AND U22165 ( .A(n14777), .B(n14778), .Z(o[3350]) );
  AND U22166 ( .A(p_input[23350]), .B(p_input[13350]), .Z(n14778) );
  AND U22167 ( .A(p_input[3350]), .B(p_input[33350]), .Z(n14777) );
  AND U22168 ( .A(n14779), .B(n14780), .Z(o[334]) );
  AND U22169 ( .A(p_input[20334]), .B(p_input[10334]), .Z(n14780) );
  AND U22170 ( .A(p_input[334]), .B(p_input[30334]), .Z(n14779) );
  AND U22171 ( .A(n14781), .B(n14782), .Z(o[3349]) );
  AND U22172 ( .A(p_input[23349]), .B(p_input[13349]), .Z(n14782) );
  AND U22173 ( .A(p_input[3349]), .B(p_input[33349]), .Z(n14781) );
  AND U22174 ( .A(n14783), .B(n14784), .Z(o[3348]) );
  AND U22175 ( .A(p_input[23348]), .B(p_input[13348]), .Z(n14784) );
  AND U22176 ( .A(p_input[3348]), .B(p_input[33348]), .Z(n14783) );
  AND U22177 ( .A(n14785), .B(n14786), .Z(o[3347]) );
  AND U22178 ( .A(p_input[23347]), .B(p_input[13347]), .Z(n14786) );
  AND U22179 ( .A(p_input[3347]), .B(p_input[33347]), .Z(n14785) );
  AND U22180 ( .A(n14787), .B(n14788), .Z(o[3346]) );
  AND U22181 ( .A(p_input[23346]), .B(p_input[13346]), .Z(n14788) );
  AND U22182 ( .A(p_input[3346]), .B(p_input[33346]), .Z(n14787) );
  AND U22183 ( .A(n14789), .B(n14790), .Z(o[3345]) );
  AND U22184 ( .A(p_input[23345]), .B(p_input[13345]), .Z(n14790) );
  AND U22185 ( .A(p_input[3345]), .B(p_input[33345]), .Z(n14789) );
  AND U22186 ( .A(n14791), .B(n14792), .Z(o[3344]) );
  AND U22187 ( .A(p_input[23344]), .B(p_input[13344]), .Z(n14792) );
  AND U22188 ( .A(p_input[3344]), .B(p_input[33344]), .Z(n14791) );
  AND U22189 ( .A(n14793), .B(n14794), .Z(o[3343]) );
  AND U22190 ( .A(p_input[23343]), .B(p_input[13343]), .Z(n14794) );
  AND U22191 ( .A(p_input[3343]), .B(p_input[33343]), .Z(n14793) );
  AND U22192 ( .A(n14795), .B(n14796), .Z(o[3342]) );
  AND U22193 ( .A(p_input[23342]), .B(p_input[13342]), .Z(n14796) );
  AND U22194 ( .A(p_input[3342]), .B(p_input[33342]), .Z(n14795) );
  AND U22195 ( .A(n14797), .B(n14798), .Z(o[3341]) );
  AND U22196 ( .A(p_input[23341]), .B(p_input[13341]), .Z(n14798) );
  AND U22197 ( .A(p_input[3341]), .B(p_input[33341]), .Z(n14797) );
  AND U22198 ( .A(n14799), .B(n14800), .Z(o[3340]) );
  AND U22199 ( .A(p_input[23340]), .B(p_input[13340]), .Z(n14800) );
  AND U22200 ( .A(p_input[3340]), .B(p_input[33340]), .Z(n14799) );
  AND U22201 ( .A(n14801), .B(n14802), .Z(o[333]) );
  AND U22202 ( .A(p_input[20333]), .B(p_input[10333]), .Z(n14802) );
  AND U22203 ( .A(p_input[333]), .B(p_input[30333]), .Z(n14801) );
  AND U22204 ( .A(n14803), .B(n14804), .Z(o[3339]) );
  AND U22205 ( .A(p_input[23339]), .B(p_input[13339]), .Z(n14804) );
  AND U22206 ( .A(p_input[3339]), .B(p_input[33339]), .Z(n14803) );
  AND U22207 ( .A(n14805), .B(n14806), .Z(o[3338]) );
  AND U22208 ( .A(p_input[23338]), .B(p_input[13338]), .Z(n14806) );
  AND U22209 ( .A(p_input[3338]), .B(p_input[33338]), .Z(n14805) );
  AND U22210 ( .A(n14807), .B(n14808), .Z(o[3337]) );
  AND U22211 ( .A(p_input[23337]), .B(p_input[13337]), .Z(n14808) );
  AND U22212 ( .A(p_input[3337]), .B(p_input[33337]), .Z(n14807) );
  AND U22213 ( .A(n14809), .B(n14810), .Z(o[3336]) );
  AND U22214 ( .A(p_input[23336]), .B(p_input[13336]), .Z(n14810) );
  AND U22215 ( .A(p_input[3336]), .B(p_input[33336]), .Z(n14809) );
  AND U22216 ( .A(n14811), .B(n14812), .Z(o[3335]) );
  AND U22217 ( .A(p_input[23335]), .B(p_input[13335]), .Z(n14812) );
  AND U22218 ( .A(p_input[3335]), .B(p_input[33335]), .Z(n14811) );
  AND U22219 ( .A(n14813), .B(n14814), .Z(o[3334]) );
  AND U22220 ( .A(p_input[23334]), .B(p_input[13334]), .Z(n14814) );
  AND U22221 ( .A(p_input[3334]), .B(p_input[33334]), .Z(n14813) );
  AND U22222 ( .A(n14815), .B(n14816), .Z(o[3333]) );
  AND U22223 ( .A(p_input[23333]), .B(p_input[13333]), .Z(n14816) );
  AND U22224 ( .A(p_input[3333]), .B(p_input[33333]), .Z(n14815) );
  AND U22225 ( .A(n14817), .B(n14818), .Z(o[3332]) );
  AND U22226 ( .A(p_input[23332]), .B(p_input[13332]), .Z(n14818) );
  AND U22227 ( .A(p_input[33332]), .B(p_input[3332]), .Z(n14817) );
  AND U22228 ( .A(n14819), .B(n14820), .Z(o[3331]) );
  AND U22229 ( .A(p_input[23331]), .B(p_input[13331]), .Z(n14820) );
  AND U22230 ( .A(p_input[33331]), .B(p_input[3331]), .Z(n14819) );
  AND U22231 ( .A(n14821), .B(n14822), .Z(o[3330]) );
  AND U22232 ( .A(p_input[23330]), .B(p_input[13330]), .Z(n14822) );
  AND U22233 ( .A(p_input[33330]), .B(p_input[3330]), .Z(n14821) );
  AND U22234 ( .A(n14823), .B(n14824), .Z(o[332]) );
  AND U22235 ( .A(p_input[20332]), .B(p_input[10332]), .Z(n14824) );
  AND U22236 ( .A(p_input[332]), .B(p_input[30332]), .Z(n14823) );
  AND U22237 ( .A(n14825), .B(n14826), .Z(o[3329]) );
  AND U22238 ( .A(p_input[23329]), .B(p_input[13329]), .Z(n14826) );
  AND U22239 ( .A(p_input[33329]), .B(p_input[3329]), .Z(n14825) );
  AND U22240 ( .A(n14827), .B(n14828), .Z(o[3328]) );
  AND U22241 ( .A(p_input[23328]), .B(p_input[13328]), .Z(n14828) );
  AND U22242 ( .A(p_input[33328]), .B(p_input[3328]), .Z(n14827) );
  AND U22243 ( .A(n14829), .B(n14830), .Z(o[3327]) );
  AND U22244 ( .A(p_input[23327]), .B(p_input[13327]), .Z(n14830) );
  AND U22245 ( .A(p_input[33327]), .B(p_input[3327]), .Z(n14829) );
  AND U22246 ( .A(n14831), .B(n14832), .Z(o[3326]) );
  AND U22247 ( .A(p_input[23326]), .B(p_input[13326]), .Z(n14832) );
  AND U22248 ( .A(p_input[33326]), .B(p_input[3326]), .Z(n14831) );
  AND U22249 ( .A(n14833), .B(n14834), .Z(o[3325]) );
  AND U22250 ( .A(p_input[23325]), .B(p_input[13325]), .Z(n14834) );
  AND U22251 ( .A(p_input[33325]), .B(p_input[3325]), .Z(n14833) );
  AND U22252 ( .A(n14835), .B(n14836), .Z(o[3324]) );
  AND U22253 ( .A(p_input[23324]), .B(p_input[13324]), .Z(n14836) );
  AND U22254 ( .A(p_input[33324]), .B(p_input[3324]), .Z(n14835) );
  AND U22255 ( .A(n14837), .B(n14838), .Z(o[3323]) );
  AND U22256 ( .A(p_input[23323]), .B(p_input[13323]), .Z(n14838) );
  AND U22257 ( .A(p_input[33323]), .B(p_input[3323]), .Z(n14837) );
  AND U22258 ( .A(n14839), .B(n14840), .Z(o[3322]) );
  AND U22259 ( .A(p_input[23322]), .B(p_input[13322]), .Z(n14840) );
  AND U22260 ( .A(p_input[33322]), .B(p_input[3322]), .Z(n14839) );
  AND U22261 ( .A(n14841), .B(n14842), .Z(o[3321]) );
  AND U22262 ( .A(p_input[23321]), .B(p_input[13321]), .Z(n14842) );
  AND U22263 ( .A(p_input[33321]), .B(p_input[3321]), .Z(n14841) );
  AND U22264 ( .A(n14843), .B(n14844), .Z(o[3320]) );
  AND U22265 ( .A(p_input[23320]), .B(p_input[13320]), .Z(n14844) );
  AND U22266 ( .A(p_input[33320]), .B(p_input[3320]), .Z(n14843) );
  AND U22267 ( .A(n14845), .B(n14846), .Z(o[331]) );
  AND U22268 ( .A(p_input[20331]), .B(p_input[10331]), .Z(n14846) );
  AND U22269 ( .A(p_input[331]), .B(p_input[30331]), .Z(n14845) );
  AND U22270 ( .A(n14847), .B(n14848), .Z(o[3319]) );
  AND U22271 ( .A(p_input[23319]), .B(p_input[13319]), .Z(n14848) );
  AND U22272 ( .A(p_input[33319]), .B(p_input[3319]), .Z(n14847) );
  AND U22273 ( .A(n14849), .B(n14850), .Z(o[3318]) );
  AND U22274 ( .A(p_input[23318]), .B(p_input[13318]), .Z(n14850) );
  AND U22275 ( .A(p_input[33318]), .B(p_input[3318]), .Z(n14849) );
  AND U22276 ( .A(n14851), .B(n14852), .Z(o[3317]) );
  AND U22277 ( .A(p_input[23317]), .B(p_input[13317]), .Z(n14852) );
  AND U22278 ( .A(p_input[33317]), .B(p_input[3317]), .Z(n14851) );
  AND U22279 ( .A(n14853), .B(n14854), .Z(o[3316]) );
  AND U22280 ( .A(p_input[23316]), .B(p_input[13316]), .Z(n14854) );
  AND U22281 ( .A(p_input[33316]), .B(p_input[3316]), .Z(n14853) );
  AND U22282 ( .A(n14855), .B(n14856), .Z(o[3315]) );
  AND U22283 ( .A(p_input[23315]), .B(p_input[13315]), .Z(n14856) );
  AND U22284 ( .A(p_input[33315]), .B(p_input[3315]), .Z(n14855) );
  AND U22285 ( .A(n14857), .B(n14858), .Z(o[3314]) );
  AND U22286 ( .A(p_input[23314]), .B(p_input[13314]), .Z(n14858) );
  AND U22287 ( .A(p_input[33314]), .B(p_input[3314]), .Z(n14857) );
  AND U22288 ( .A(n14859), .B(n14860), .Z(o[3313]) );
  AND U22289 ( .A(p_input[23313]), .B(p_input[13313]), .Z(n14860) );
  AND U22290 ( .A(p_input[33313]), .B(p_input[3313]), .Z(n14859) );
  AND U22291 ( .A(n14861), .B(n14862), .Z(o[3312]) );
  AND U22292 ( .A(p_input[23312]), .B(p_input[13312]), .Z(n14862) );
  AND U22293 ( .A(p_input[33312]), .B(p_input[3312]), .Z(n14861) );
  AND U22294 ( .A(n14863), .B(n14864), .Z(o[3311]) );
  AND U22295 ( .A(p_input[23311]), .B(p_input[13311]), .Z(n14864) );
  AND U22296 ( .A(p_input[33311]), .B(p_input[3311]), .Z(n14863) );
  AND U22297 ( .A(n14865), .B(n14866), .Z(o[3310]) );
  AND U22298 ( .A(p_input[23310]), .B(p_input[13310]), .Z(n14866) );
  AND U22299 ( .A(p_input[33310]), .B(p_input[3310]), .Z(n14865) );
  AND U22300 ( .A(n14867), .B(n14868), .Z(o[330]) );
  AND U22301 ( .A(p_input[20330]), .B(p_input[10330]), .Z(n14868) );
  AND U22302 ( .A(p_input[330]), .B(p_input[30330]), .Z(n14867) );
  AND U22303 ( .A(n14869), .B(n14870), .Z(o[3309]) );
  AND U22304 ( .A(p_input[23309]), .B(p_input[13309]), .Z(n14870) );
  AND U22305 ( .A(p_input[33309]), .B(p_input[3309]), .Z(n14869) );
  AND U22306 ( .A(n14871), .B(n14872), .Z(o[3308]) );
  AND U22307 ( .A(p_input[23308]), .B(p_input[13308]), .Z(n14872) );
  AND U22308 ( .A(p_input[33308]), .B(p_input[3308]), .Z(n14871) );
  AND U22309 ( .A(n14873), .B(n14874), .Z(o[3307]) );
  AND U22310 ( .A(p_input[23307]), .B(p_input[13307]), .Z(n14874) );
  AND U22311 ( .A(p_input[33307]), .B(p_input[3307]), .Z(n14873) );
  AND U22312 ( .A(n14875), .B(n14876), .Z(o[3306]) );
  AND U22313 ( .A(p_input[23306]), .B(p_input[13306]), .Z(n14876) );
  AND U22314 ( .A(p_input[33306]), .B(p_input[3306]), .Z(n14875) );
  AND U22315 ( .A(n14877), .B(n14878), .Z(o[3305]) );
  AND U22316 ( .A(p_input[23305]), .B(p_input[13305]), .Z(n14878) );
  AND U22317 ( .A(p_input[33305]), .B(p_input[3305]), .Z(n14877) );
  AND U22318 ( .A(n14879), .B(n14880), .Z(o[3304]) );
  AND U22319 ( .A(p_input[23304]), .B(p_input[13304]), .Z(n14880) );
  AND U22320 ( .A(p_input[33304]), .B(p_input[3304]), .Z(n14879) );
  AND U22321 ( .A(n14881), .B(n14882), .Z(o[3303]) );
  AND U22322 ( .A(p_input[23303]), .B(p_input[13303]), .Z(n14882) );
  AND U22323 ( .A(p_input[33303]), .B(p_input[3303]), .Z(n14881) );
  AND U22324 ( .A(n14883), .B(n14884), .Z(o[3302]) );
  AND U22325 ( .A(p_input[23302]), .B(p_input[13302]), .Z(n14884) );
  AND U22326 ( .A(p_input[33302]), .B(p_input[3302]), .Z(n14883) );
  AND U22327 ( .A(n14885), .B(n14886), .Z(o[3301]) );
  AND U22328 ( .A(p_input[23301]), .B(p_input[13301]), .Z(n14886) );
  AND U22329 ( .A(p_input[33301]), .B(p_input[3301]), .Z(n14885) );
  AND U22330 ( .A(n14887), .B(n14888), .Z(o[3300]) );
  AND U22331 ( .A(p_input[23300]), .B(p_input[13300]), .Z(n14888) );
  AND U22332 ( .A(p_input[33300]), .B(p_input[3300]), .Z(n14887) );
  AND U22333 ( .A(n14889), .B(n14890), .Z(o[32]) );
  AND U22334 ( .A(p_input[20032]), .B(p_input[10032]), .Z(n14890) );
  AND U22335 ( .A(p_input[32]), .B(p_input[30032]), .Z(n14889) );
  AND U22336 ( .A(n14891), .B(n14892), .Z(o[329]) );
  AND U22337 ( .A(p_input[20329]), .B(p_input[10329]), .Z(n14892) );
  AND U22338 ( .A(p_input[329]), .B(p_input[30329]), .Z(n14891) );
  AND U22339 ( .A(n14893), .B(n14894), .Z(o[3299]) );
  AND U22340 ( .A(p_input[23299]), .B(p_input[13299]), .Z(n14894) );
  AND U22341 ( .A(p_input[33299]), .B(p_input[3299]), .Z(n14893) );
  AND U22342 ( .A(n14895), .B(n14896), .Z(o[3298]) );
  AND U22343 ( .A(p_input[23298]), .B(p_input[13298]), .Z(n14896) );
  AND U22344 ( .A(p_input[33298]), .B(p_input[3298]), .Z(n14895) );
  AND U22345 ( .A(n14897), .B(n14898), .Z(o[3297]) );
  AND U22346 ( .A(p_input[23297]), .B(p_input[13297]), .Z(n14898) );
  AND U22347 ( .A(p_input[33297]), .B(p_input[3297]), .Z(n14897) );
  AND U22348 ( .A(n14899), .B(n14900), .Z(o[3296]) );
  AND U22349 ( .A(p_input[23296]), .B(p_input[13296]), .Z(n14900) );
  AND U22350 ( .A(p_input[33296]), .B(p_input[3296]), .Z(n14899) );
  AND U22351 ( .A(n14901), .B(n14902), .Z(o[3295]) );
  AND U22352 ( .A(p_input[23295]), .B(p_input[13295]), .Z(n14902) );
  AND U22353 ( .A(p_input[33295]), .B(p_input[3295]), .Z(n14901) );
  AND U22354 ( .A(n14903), .B(n14904), .Z(o[3294]) );
  AND U22355 ( .A(p_input[23294]), .B(p_input[13294]), .Z(n14904) );
  AND U22356 ( .A(p_input[33294]), .B(p_input[3294]), .Z(n14903) );
  AND U22357 ( .A(n14905), .B(n14906), .Z(o[3293]) );
  AND U22358 ( .A(p_input[23293]), .B(p_input[13293]), .Z(n14906) );
  AND U22359 ( .A(p_input[33293]), .B(p_input[3293]), .Z(n14905) );
  AND U22360 ( .A(n14907), .B(n14908), .Z(o[3292]) );
  AND U22361 ( .A(p_input[23292]), .B(p_input[13292]), .Z(n14908) );
  AND U22362 ( .A(p_input[33292]), .B(p_input[3292]), .Z(n14907) );
  AND U22363 ( .A(n14909), .B(n14910), .Z(o[3291]) );
  AND U22364 ( .A(p_input[23291]), .B(p_input[13291]), .Z(n14910) );
  AND U22365 ( .A(p_input[33291]), .B(p_input[3291]), .Z(n14909) );
  AND U22366 ( .A(n14911), .B(n14912), .Z(o[3290]) );
  AND U22367 ( .A(p_input[23290]), .B(p_input[13290]), .Z(n14912) );
  AND U22368 ( .A(p_input[33290]), .B(p_input[3290]), .Z(n14911) );
  AND U22369 ( .A(n14913), .B(n14914), .Z(o[328]) );
  AND U22370 ( .A(p_input[20328]), .B(p_input[10328]), .Z(n14914) );
  AND U22371 ( .A(p_input[328]), .B(p_input[30328]), .Z(n14913) );
  AND U22372 ( .A(n14915), .B(n14916), .Z(o[3289]) );
  AND U22373 ( .A(p_input[23289]), .B(p_input[13289]), .Z(n14916) );
  AND U22374 ( .A(p_input[33289]), .B(p_input[3289]), .Z(n14915) );
  AND U22375 ( .A(n14917), .B(n14918), .Z(o[3288]) );
  AND U22376 ( .A(p_input[23288]), .B(p_input[13288]), .Z(n14918) );
  AND U22377 ( .A(p_input[33288]), .B(p_input[3288]), .Z(n14917) );
  AND U22378 ( .A(n14919), .B(n14920), .Z(o[3287]) );
  AND U22379 ( .A(p_input[23287]), .B(p_input[13287]), .Z(n14920) );
  AND U22380 ( .A(p_input[33287]), .B(p_input[3287]), .Z(n14919) );
  AND U22381 ( .A(n14921), .B(n14922), .Z(o[3286]) );
  AND U22382 ( .A(p_input[23286]), .B(p_input[13286]), .Z(n14922) );
  AND U22383 ( .A(p_input[33286]), .B(p_input[3286]), .Z(n14921) );
  AND U22384 ( .A(n14923), .B(n14924), .Z(o[3285]) );
  AND U22385 ( .A(p_input[23285]), .B(p_input[13285]), .Z(n14924) );
  AND U22386 ( .A(p_input[33285]), .B(p_input[3285]), .Z(n14923) );
  AND U22387 ( .A(n14925), .B(n14926), .Z(o[3284]) );
  AND U22388 ( .A(p_input[23284]), .B(p_input[13284]), .Z(n14926) );
  AND U22389 ( .A(p_input[33284]), .B(p_input[3284]), .Z(n14925) );
  AND U22390 ( .A(n14927), .B(n14928), .Z(o[3283]) );
  AND U22391 ( .A(p_input[23283]), .B(p_input[13283]), .Z(n14928) );
  AND U22392 ( .A(p_input[33283]), .B(p_input[3283]), .Z(n14927) );
  AND U22393 ( .A(n14929), .B(n14930), .Z(o[3282]) );
  AND U22394 ( .A(p_input[23282]), .B(p_input[13282]), .Z(n14930) );
  AND U22395 ( .A(p_input[33282]), .B(p_input[3282]), .Z(n14929) );
  AND U22396 ( .A(n14931), .B(n14932), .Z(o[3281]) );
  AND U22397 ( .A(p_input[23281]), .B(p_input[13281]), .Z(n14932) );
  AND U22398 ( .A(p_input[33281]), .B(p_input[3281]), .Z(n14931) );
  AND U22399 ( .A(n14933), .B(n14934), .Z(o[3280]) );
  AND U22400 ( .A(p_input[23280]), .B(p_input[13280]), .Z(n14934) );
  AND U22401 ( .A(p_input[33280]), .B(p_input[3280]), .Z(n14933) );
  AND U22402 ( .A(n14935), .B(n14936), .Z(o[327]) );
  AND U22403 ( .A(p_input[20327]), .B(p_input[10327]), .Z(n14936) );
  AND U22404 ( .A(p_input[327]), .B(p_input[30327]), .Z(n14935) );
  AND U22405 ( .A(n14937), .B(n14938), .Z(o[3279]) );
  AND U22406 ( .A(p_input[23279]), .B(p_input[13279]), .Z(n14938) );
  AND U22407 ( .A(p_input[33279]), .B(p_input[3279]), .Z(n14937) );
  AND U22408 ( .A(n14939), .B(n14940), .Z(o[3278]) );
  AND U22409 ( .A(p_input[23278]), .B(p_input[13278]), .Z(n14940) );
  AND U22410 ( .A(p_input[33278]), .B(p_input[3278]), .Z(n14939) );
  AND U22411 ( .A(n14941), .B(n14942), .Z(o[3277]) );
  AND U22412 ( .A(p_input[23277]), .B(p_input[13277]), .Z(n14942) );
  AND U22413 ( .A(p_input[33277]), .B(p_input[3277]), .Z(n14941) );
  AND U22414 ( .A(n14943), .B(n14944), .Z(o[3276]) );
  AND U22415 ( .A(p_input[23276]), .B(p_input[13276]), .Z(n14944) );
  AND U22416 ( .A(p_input[33276]), .B(p_input[3276]), .Z(n14943) );
  AND U22417 ( .A(n14945), .B(n14946), .Z(o[3275]) );
  AND U22418 ( .A(p_input[23275]), .B(p_input[13275]), .Z(n14946) );
  AND U22419 ( .A(p_input[33275]), .B(p_input[3275]), .Z(n14945) );
  AND U22420 ( .A(n14947), .B(n14948), .Z(o[3274]) );
  AND U22421 ( .A(p_input[23274]), .B(p_input[13274]), .Z(n14948) );
  AND U22422 ( .A(p_input[33274]), .B(p_input[3274]), .Z(n14947) );
  AND U22423 ( .A(n14949), .B(n14950), .Z(o[3273]) );
  AND U22424 ( .A(p_input[23273]), .B(p_input[13273]), .Z(n14950) );
  AND U22425 ( .A(p_input[33273]), .B(p_input[3273]), .Z(n14949) );
  AND U22426 ( .A(n14951), .B(n14952), .Z(o[3272]) );
  AND U22427 ( .A(p_input[23272]), .B(p_input[13272]), .Z(n14952) );
  AND U22428 ( .A(p_input[33272]), .B(p_input[3272]), .Z(n14951) );
  AND U22429 ( .A(n14953), .B(n14954), .Z(o[3271]) );
  AND U22430 ( .A(p_input[23271]), .B(p_input[13271]), .Z(n14954) );
  AND U22431 ( .A(p_input[33271]), .B(p_input[3271]), .Z(n14953) );
  AND U22432 ( .A(n14955), .B(n14956), .Z(o[3270]) );
  AND U22433 ( .A(p_input[23270]), .B(p_input[13270]), .Z(n14956) );
  AND U22434 ( .A(p_input[33270]), .B(p_input[3270]), .Z(n14955) );
  AND U22435 ( .A(n14957), .B(n14958), .Z(o[326]) );
  AND U22436 ( .A(p_input[20326]), .B(p_input[10326]), .Z(n14958) );
  AND U22437 ( .A(p_input[326]), .B(p_input[30326]), .Z(n14957) );
  AND U22438 ( .A(n14959), .B(n14960), .Z(o[3269]) );
  AND U22439 ( .A(p_input[23269]), .B(p_input[13269]), .Z(n14960) );
  AND U22440 ( .A(p_input[33269]), .B(p_input[3269]), .Z(n14959) );
  AND U22441 ( .A(n14961), .B(n14962), .Z(o[3268]) );
  AND U22442 ( .A(p_input[23268]), .B(p_input[13268]), .Z(n14962) );
  AND U22443 ( .A(p_input[33268]), .B(p_input[3268]), .Z(n14961) );
  AND U22444 ( .A(n14963), .B(n14964), .Z(o[3267]) );
  AND U22445 ( .A(p_input[23267]), .B(p_input[13267]), .Z(n14964) );
  AND U22446 ( .A(p_input[33267]), .B(p_input[3267]), .Z(n14963) );
  AND U22447 ( .A(n14965), .B(n14966), .Z(o[3266]) );
  AND U22448 ( .A(p_input[23266]), .B(p_input[13266]), .Z(n14966) );
  AND U22449 ( .A(p_input[33266]), .B(p_input[3266]), .Z(n14965) );
  AND U22450 ( .A(n14967), .B(n14968), .Z(o[3265]) );
  AND U22451 ( .A(p_input[23265]), .B(p_input[13265]), .Z(n14968) );
  AND U22452 ( .A(p_input[33265]), .B(p_input[3265]), .Z(n14967) );
  AND U22453 ( .A(n14969), .B(n14970), .Z(o[3264]) );
  AND U22454 ( .A(p_input[23264]), .B(p_input[13264]), .Z(n14970) );
  AND U22455 ( .A(p_input[33264]), .B(p_input[3264]), .Z(n14969) );
  AND U22456 ( .A(n14971), .B(n14972), .Z(o[3263]) );
  AND U22457 ( .A(p_input[23263]), .B(p_input[13263]), .Z(n14972) );
  AND U22458 ( .A(p_input[33263]), .B(p_input[3263]), .Z(n14971) );
  AND U22459 ( .A(n14973), .B(n14974), .Z(o[3262]) );
  AND U22460 ( .A(p_input[23262]), .B(p_input[13262]), .Z(n14974) );
  AND U22461 ( .A(p_input[33262]), .B(p_input[3262]), .Z(n14973) );
  AND U22462 ( .A(n14975), .B(n14976), .Z(o[3261]) );
  AND U22463 ( .A(p_input[23261]), .B(p_input[13261]), .Z(n14976) );
  AND U22464 ( .A(p_input[33261]), .B(p_input[3261]), .Z(n14975) );
  AND U22465 ( .A(n14977), .B(n14978), .Z(o[3260]) );
  AND U22466 ( .A(p_input[23260]), .B(p_input[13260]), .Z(n14978) );
  AND U22467 ( .A(p_input[33260]), .B(p_input[3260]), .Z(n14977) );
  AND U22468 ( .A(n14979), .B(n14980), .Z(o[325]) );
  AND U22469 ( .A(p_input[20325]), .B(p_input[10325]), .Z(n14980) );
  AND U22470 ( .A(p_input[325]), .B(p_input[30325]), .Z(n14979) );
  AND U22471 ( .A(n14981), .B(n14982), .Z(o[3259]) );
  AND U22472 ( .A(p_input[23259]), .B(p_input[13259]), .Z(n14982) );
  AND U22473 ( .A(p_input[33259]), .B(p_input[3259]), .Z(n14981) );
  AND U22474 ( .A(n14983), .B(n14984), .Z(o[3258]) );
  AND U22475 ( .A(p_input[23258]), .B(p_input[13258]), .Z(n14984) );
  AND U22476 ( .A(p_input[33258]), .B(p_input[3258]), .Z(n14983) );
  AND U22477 ( .A(n14985), .B(n14986), .Z(o[3257]) );
  AND U22478 ( .A(p_input[23257]), .B(p_input[13257]), .Z(n14986) );
  AND U22479 ( .A(p_input[33257]), .B(p_input[3257]), .Z(n14985) );
  AND U22480 ( .A(n14987), .B(n14988), .Z(o[3256]) );
  AND U22481 ( .A(p_input[23256]), .B(p_input[13256]), .Z(n14988) );
  AND U22482 ( .A(p_input[33256]), .B(p_input[3256]), .Z(n14987) );
  AND U22483 ( .A(n14989), .B(n14990), .Z(o[3255]) );
  AND U22484 ( .A(p_input[23255]), .B(p_input[13255]), .Z(n14990) );
  AND U22485 ( .A(p_input[33255]), .B(p_input[3255]), .Z(n14989) );
  AND U22486 ( .A(n14991), .B(n14992), .Z(o[3254]) );
  AND U22487 ( .A(p_input[23254]), .B(p_input[13254]), .Z(n14992) );
  AND U22488 ( .A(p_input[33254]), .B(p_input[3254]), .Z(n14991) );
  AND U22489 ( .A(n14993), .B(n14994), .Z(o[3253]) );
  AND U22490 ( .A(p_input[23253]), .B(p_input[13253]), .Z(n14994) );
  AND U22491 ( .A(p_input[33253]), .B(p_input[3253]), .Z(n14993) );
  AND U22492 ( .A(n14995), .B(n14996), .Z(o[3252]) );
  AND U22493 ( .A(p_input[23252]), .B(p_input[13252]), .Z(n14996) );
  AND U22494 ( .A(p_input[33252]), .B(p_input[3252]), .Z(n14995) );
  AND U22495 ( .A(n14997), .B(n14998), .Z(o[3251]) );
  AND U22496 ( .A(p_input[23251]), .B(p_input[13251]), .Z(n14998) );
  AND U22497 ( .A(p_input[33251]), .B(p_input[3251]), .Z(n14997) );
  AND U22498 ( .A(n14999), .B(n15000), .Z(o[3250]) );
  AND U22499 ( .A(p_input[23250]), .B(p_input[13250]), .Z(n15000) );
  AND U22500 ( .A(p_input[33250]), .B(p_input[3250]), .Z(n14999) );
  AND U22501 ( .A(n15001), .B(n15002), .Z(o[324]) );
  AND U22502 ( .A(p_input[20324]), .B(p_input[10324]), .Z(n15002) );
  AND U22503 ( .A(p_input[324]), .B(p_input[30324]), .Z(n15001) );
  AND U22504 ( .A(n15003), .B(n15004), .Z(o[3249]) );
  AND U22505 ( .A(p_input[23249]), .B(p_input[13249]), .Z(n15004) );
  AND U22506 ( .A(p_input[33249]), .B(p_input[3249]), .Z(n15003) );
  AND U22507 ( .A(n15005), .B(n15006), .Z(o[3248]) );
  AND U22508 ( .A(p_input[23248]), .B(p_input[13248]), .Z(n15006) );
  AND U22509 ( .A(p_input[33248]), .B(p_input[3248]), .Z(n15005) );
  AND U22510 ( .A(n15007), .B(n15008), .Z(o[3247]) );
  AND U22511 ( .A(p_input[23247]), .B(p_input[13247]), .Z(n15008) );
  AND U22512 ( .A(p_input[33247]), .B(p_input[3247]), .Z(n15007) );
  AND U22513 ( .A(n15009), .B(n15010), .Z(o[3246]) );
  AND U22514 ( .A(p_input[23246]), .B(p_input[13246]), .Z(n15010) );
  AND U22515 ( .A(p_input[33246]), .B(p_input[3246]), .Z(n15009) );
  AND U22516 ( .A(n15011), .B(n15012), .Z(o[3245]) );
  AND U22517 ( .A(p_input[23245]), .B(p_input[13245]), .Z(n15012) );
  AND U22518 ( .A(p_input[33245]), .B(p_input[3245]), .Z(n15011) );
  AND U22519 ( .A(n15013), .B(n15014), .Z(o[3244]) );
  AND U22520 ( .A(p_input[23244]), .B(p_input[13244]), .Z(n15014) );
  AND U22521 ( .A(p_input[33244]), .B(p_input[3244]), .Z(n15013) );
  AND U22522 ( .A(n15015), .B(n15016), .Z(o[3243]) );
  AND U22523 ( .A(p_input[23243]), .B(p_input[13243]), .Z(n15016) );
  AND U22524 ( .A(p_input[33243]), .B(p_input[3243]), .Z(n15015) );
  AND U22525 ( .A(n15017), .B(n15018), .Z(o[3242]) );
  AND U22526 ( .A(p_input[23242]), .B(p_input[13242]), .Z(n15018) );
  AND U22527 ( .A(p_input[33242]), .B(p_input[3242]), .Z(n15017) );
  AND U22528 ( .A(n15019), .B(n15020), .Z(o[3241]) );
  AND U22529 ( .A(p_input[23241]), .B(p_input[13241]), .Z(n15020) );
  AND U22530 ( .A(p_input[33241]), .B(p_input[3241]), .Z(n15019) );
  AND U22531 ( .A(n15021), .B(n15022), .Z(o[3240]) );
  AND U22532 ( .A(p_input[23240]), .B(p_input[13240]), .Z(n15022) );
  AND U22533 ( .A(p_input[33240]), .B(p_input[3240]), .Z(n15021) );
  AND U22534 ( .A(n15023), .B(n15024), .Z(o[323]) );
  AND U22535 ( .A(p_input[20323]), .B(p_input[10323]), .Z(n15024) );
  AND U22536 ( .A(p_input[323]), .B(p_input[30323]), .Z(n15023) );
  AND U22537 ( .A(n15025), .B(n15026), .Z(o[3239]) );
  AND U22538 ( .A(p_input[23239]), .B(p_input[13239]), .Z(n15026) );
  AND U22539 ( .A(p_input[33239]), .B(p_input[3239]), .Z(n15025) );
  AND U22540 ( .A(n15027), .B(n15028), .Z(o[3238]) );
  AND U22541 ( .A(p_input[23238]), .B(p_input[13238]), .Z(n15028) );
  AND U22542 ( .A(p_input[33238]), .B(p_input[3238]), .Z(n15027) );
  AND U22543 ( .A(n15029), .B(n15030), .Z(o[3237]) );
  AND U22544 ( .A(p_input[23237]), .B(p_input[13237]), .Z(n15030) );
  AND U22545 ( .A(p_input[33237]), .B(p_input[3237]), .Z(n15029) );
  AND U22546 ( .A(n15031), .B(n15032), .Z(o[3236]) );
  AND U22547 ( .A(p_input[23236]), .B(p_input[13236]), .Z(n15032) );
  AND U22548 ( .A(p_input[33236]), .B(p_input[3236]), .Z(n15031) );
  AND U22549 ( .A(n15033), .B(n15034), .Z(o[3235]) );
  AND U22550 ( .A(p_input[23235]), .B(p_input[13235]), .Z(n15034) );
  AND U22551 ( .A(p_input[33235]), .B(p_input[3235]), .Z(n15033) );
  AND U22552 ( .A(n15035), .B(n15036), .Z(o[3234]) );
  AND U22553 ( .A(p_input[23234]), .B(p_input[13234]), .Z(n15036) );
  AND U22554 ( .A(p_input[33234]), .B(p_input[3234]), .Z(n15035) );
  AND U22555 ( .A(n15037), .B(n15038), .Z(o[3233]) );
  AND U22556 ( .A(p_input[23233]), .B(p_input[13233]), .Z(n15038) );
  AND U22557 ( .A(p_input[33233]), .B(p_input[3233]), .Z(n15037) );
  AND U22558 ( .A(n15039), .B(n15040), .Z(o[3232]) );
  AND U22559 ( .A(p_input[23232]), .B(p_input[13232]), .Z(n15040) );
  AND U22560 ( .A(p_input[33232]), .B(p_input[3232]), .Z(n15039) );
  AND U22561 ( .A(n15041), .B(n15042), .Z(o[3231]) );
  AND U22562 ( .A(p_input[23231]), .B(p_input[13231]), .Z(n15042) );
  AND U22563 ( .A(p_input[33231]), .B(p_input[3231]), .Z(n15041) );
  AND U22564 ( .A(n15043), .B(n15044), .Z(o[3230]) );
  AND U22565 ( .A(p_input[23230]), .B(p_input[13230]), .Z(n15044) );
  AND U22566 ( .A(p_input[33230]), .B(p_input[3230]), .Z(n15043) );
  AND U22567 ( .A(n15045), .B(n15046), .Z(o[322]) );
  AND U22568 ( .A(p_input[20322]), .B(p_input[10322]), .Z(n15046) );
  AND U22569 ( .A(p_input[322]), .B(p_input[30322]), .Z(n15045) );
  AND U22570 ( .A(n15047), .B(n15048), .Z(o[3229]) );
  AND U22571 ( .A(p_input[23229]), .B(p_input[13229]), .Z(n15048) );
  AND U22572 ( .A(p_input[33229]), .B(p_input[3229]), .Z(n15047) );
  AND U22573 ( .A(n15049), .B(n15050), .Z(o[3228]) );
  AND U22574 ( .A(p_input[23228]), .B(p_input[13228]), .Z(n15050) );
  AND U22575 ( .A(p_input[33228]), .B(p_input[3228]), .Z(n15049) );
  AND U22576 ( .A(n15051), .B(n15052), .Z(o[3227]) );
  AND U22577 ( .A(p_input[23227]), .B(p_input[13227]), .Z(n15052) );
  AND U22578 ( .A(p_input[33227]), .B(p_input[3227]), .Z(n15051) );
  AND U22579 ( .A(n15053), .B(n15054), .Z(o[3226]) );
  AND U22580 ( .A(p_input[23226]), .B(p_input[13226]), .Z(n15054) );
  AND U22581 ( .A(p_input[33226]), .B(p_input[3226]), .Z(n15053) );
  AND U22582 ( .A(n15055), .B(n15056), .Z(o[3225]) );
  AND U22583 ( .A(p_input[23225]), .B(p_input[13225]), .Z(n15056) );
  AND U22584 ( .A(p_input[33225]), .B(p_input[3225]), .Z(n15055) );
  AND U22585 ( .A(n15057), .B(n15058), .Z(o[3224]) );
  AND U22586 ( .A(p_input[23224]), .B(p_input[13224]), .Z(n15058) );
  AND U22587 ( .A(p_input[33224]), .B(p_input[3224]), .Z(n15057) );
  AND U22588 ( .A(n15059), .B(n15060), .Z(o[3223]) );
  AND U22589 ( .A(p_input[23223]), .B(p_input[13223]), .Z(n15060) );
  AND U22590 ( .A(p_input[33223]), .B(p_input[3223]), .Z(n15059) );
  AND U22591 ( .A(n15061), .B(n15062), .Z(o[3222]) );
  AND U22592 ( .A(p_input[23222]), .B(p_input[13222]), .Z(n15062) );
  AND U22593 ( .A(p_input[33222]), .B(p_input[3222]), .Z(n15061) );
  AND U22594 ( .A(n15063), .B(n15064), .Z(o[3221]) );
  AND U22595 ( .A(p_input[23221]), .B(p_input[13221]), .Z(n15064) );
  AND U22596 ( .A(p_input[33221]), .B(p_input[3221]), .Z(n15063) );
  AND U22597 ( .A(n15065), .B(n15066), .Z(o[3220]) );
  AND U22598 ( .A(p_input[23220]), .B(p_input[13220]), .Z(n15066) );
  AND U22599 ( .A(p_input[33220]), .B(p_input[3220]), .Z(n15065) );
  AND U22600 ( .A(n15067), .B(n15068), .Z(o[321]) );
  AND U22601 ( .A(p_input[20321]), .B(p_input[10321]), .Z(n15068) );
  AND U22602 ( .A(p_input[321]), .B(p_input[30321]), .Z(n15067) );
  AND U22603 ( .A(n15069), .B(n15070), .Z(o[3219]) );
  AND U22604 ( .A(p_input[23219]), .B(p_input[13219]), .Z(n15070) );
  AND U22605 ( .A(p_input[33219]), .B(p_input[3219]), .Z(n15069) );
  AND U22606 ( .A(n15071), .B(n15072), .Z(o[3218]) );
  AND U22607 ( .A(p_input[23218]), .B(p_input[13218]), .Z(n15072) );
  AND U22608 ( .A(p_input[33218]), .B(p_input[3218]), .Z(n15071) );
  AND U22609 ( .A(n15073), .B(n15074), .Z(o[3217]) );
  AND U22610 ( .A(p_input[23217]), .B(p_input[13217]), .Z(n15074) );
  AND U22611 ( .A(p_input[33217]), .B(p_input[3217]), .Z(n15073) );
  AND U22612 ( .A(n15075), .B(n15076), .Z(o[3216]) );
  AND U22613 ( .A(p_input[23216]), .B(p_input[13216]), .Z(n15076) );
  AND U22614 ( .A(p_input[33216]), .B(p_input[3216]), .Z(n15075) );
  AND U22615 ( .A(n15077), .B(n15078), .Z(o[3215]) );
  AND U22616 ( .A(p_input[23215]), .B(p_input[13215]), .Z(n15078) );
  AND U22617 ( .A(p_input[33215]), .B(p_input[3215]), .Z(n15077) );
  AND U22618 ( .A(n15079), .B(n15080), .Z(o[3214]) );
  AND U22619 ( .A(p_input[23214]), .B(p_input[13214]), .Z(n15080) );
  AND U22620 ( .A(p_input[33214]), .B(p_input[3214]), .Z(n15079) );
  AND U22621 ( .A(n15081), .B(n15082), .Z(o[3213]) );
  AND U22622 ( .A(p_input[23213]), .B(p_input[13213]), .Z(n15082) );
  AND U22623 ( .A(p_input[33213]), .B(p_input[3213]), .Z(n15081) );
  AND U22624 ( .A(n15083), .B(n15084), .Z(o[3212]) );
  AND U22625 ( .A(p_input[23212]), .B(p_input[13212]), .Z(n15084) );
  AND U22626 ( .A(p_input[33212]), .B(p_input[3212]), .Z(n15083) );
  AND U22627 ( .A(n15085), .B(n15086), .Z(o[3211]) );
  AND U22628 ( .A(p_input[23211]), .B(p_input[13211]), .Z(n15086) );
  AND U22629 ( .A(p_input[33211]), .B(p_input[3211]), .Z(n15085) );
  AND U22630 ( .A(n15087), .B(n15088), .Z(o[3210]) );
  AND U22631 ( .A(p_input[23210]), .B(p_input[13210]), .Z(n15088) );
  AND U22632 ( .A(p_input[33210]), .B(p_input[3210]), .Z(n15087) );
  AND U22633 ( .A(n15089), .B(n15090), .Z(o[320]) );
  AND U22634 ( .A(p_input[20320]), .B(p_input[10320]), .Z(n15090) );
  AND U22635 ( .A(p_input[320]), .B(p_input[30320]), .Z(n15089) );
  AND U22636 ( .A(n15091), .B(n15092), .Z(o[3209]) );
  AND U22637 ( .A(p_input[23209]), .B(p_input[13209]), .Z(n15092) );
  AND U22638 ( .A(p_input[33209]), .B(p_input[3209]), .Z(n15091) );
  AND U22639 ( .A(n15093), .B(n15094), .Z(o[3208]) );
  AND U22640 ( .A(p_input[23208]), .B(p_input[13208]), .Z(n15094) );
  AND U22641 ( .A(p_input[33208]), .B(p_input[3208]), .Z(n15093) );
  AND U22642 ( .A(n15095), .B(n15096), .Z(o[3207]) );
  AND U22643 ( .A(p_input[23207]), .B(p_input[13207]), .Z(n15096) );
  AND U22644 ( .A(p_input[33207]), .B(p_input[3207]), .Z(n15095) );
  AND U22645 ( .A(n15097), .B(n15098), .Z(o[3206]) );
  AND U22646 ( .A(p_input[23206]), .B(p_input[13206]), .Z(n15098) );
  AND U22647 ( .A(p_input[33206]), .B(p_input[3206]), .Z(n15097) );
  AND U22648 ( .A(n15099), .B(n15100), .Z(o[3205]) );
  AND U22649 ( .A(p_input[23205]), .B(p_input[13205]), .Z(n15100) );
  AND U22650 ( .A(p_input[33205]), .B(p_input[3205]), .Z(n15099) );
  AND U22651 ( .A(n15101), .B(n15102), .Z(o[3204]) );
  AND U22652 ( .A(p_input[23204]), .B(p_input[13204]), .Z(n15102) );
  AND U22653 ( .A(p_input[33204]), .B(p_input[3204]), .Z(n15101) );
  AND U22654 ( .A(n15103), .B(n15104), .Z(o[3203]) );
  AND U22655 ( .A(p_input[23203]), .B(p_input[13203]), .Z(n15104) );
  AND U22656 ( .A(p_input[33203]), .B(p_input[3203]), .Z(n15103) );
  AND U22657 ( .A(n15105), .B(n15106), .Z(o[3202]) );
  AND U22658 ( .A(p_input[23202]), .B(p_input[13202]), .Z(n15106) );
  AND U22659 ( .A(p_input[33202]), .B(p_input[3202]), .Z(n15105) );
  AND U22660 ( .A(n15107), .B(n15108), .Z(o[3201]) );
  AND U22661 ( .A(p_input[23201]), .B(p_input[13201]), .Z(n15108) );
  AND U22662 ( .A(p_input[33201]), .B(p_input[3201]), .Z(n15107) );
  AND U22663 ( .A(n15109), .B(n15110), .Z(o[3200]) );
  AND U22664 ( .A(p_input[23200]), .B(p_input[13200]), .Z(n15110) );
  AND U22665 ( .A(p_input[33200]), .B(p_input[3200]), .Z(n15109) );
  AND U22666 ( .A(n15111), .B(n15112), .Z(o[31]) );
  AND U22667 ( .A(p_input[20031]), .B(p_input[10031]), .Z(n15112) );
  AND U22668 ( .A(p_input[31]), .B(p_input[30031]), .Z(n15111) );
  AND U22669 ( .A(n15113), .B(n15114), .Z(o[319]) );
  AND U22670 ( .A(p_input[20319]), .B(p_input[10319]), .Z(n15114) );
  AND U22671 ( .A(p_input[319]), .B(p_input[30319]), .Z(n15113) );
  AND U22672 ( .A(n15115), .B(n15116), .Z(o[3199]) );
  AND U22673 ( .A(p_input[23199]), .B(p_input[13199]), .Z(n15116) );
  AND U22674 ( .A(p_input[33199]), .B(p_input[3199]), .Z(n15115) );
  AND U22675 ( .A(n15117), .B(n15118), .Z(o[3198]) );
  AND U22676 ( .A(p_input[23198]), .B(p_input[13198]), .Z(n15118) );
  AND U22677 ( .A(p_input[33198]), .B(p_input[3198]), .Z(n15117) );
  AND U22678 ( .A(n15119), .B(n15120), .Z(o[3197]) );
  AND U22679 ( .A(p_input[23197]), .B(p_input[13197]), .Z(n15120) );
  AND U22680 ( .A(p_input[33197]), .B(p_input[3197]), .Z(n15119) );
  AND U22681 ( .A(n15121), .B(n15122), .Z(o[3196]) );
  AND U22682 ( .A(p_input[23196]), .B(p_input[13196]), .Z(n15122) );
  AND U22683 ( .A(p_input[33196]), .B(p_input[3196]), .Z(n15121) );
  AND U22684 ( .A(n15123), .B(n15124), .Z(o[3195]) );
  AND U22685 ( .A(p_input[23195]), .B(p_input[13195]), .Z(n15124) );
  AND U22686 ( .A(p_input[33195]), .B(p_input[3195]), .Z(n15123) );
  AND U22687 ( .A(n15125), .B(n15126), .Z(o[3194]) );
  AND U22688 ( .A(p_input[23194]), .B(p_input[13194]), .Z(n15126) );
  AND U22689 ( .A(p_input[33194]), .B(p_input[3194]), .Z(n15125) );
  AND U22690 ( .A(n15127), .B(n15128), .Z(o[3193]) );
  AND U22691 ( .A(p_input[23193]), .B(p_input[13193]), .Z(n15128) );
  AND U22692 ( .A(p_input[33193]), .B(p_input[3193]), .Z(n15127) );
  AND U22693 ( .A(n15129), .B(n15130), .Z(o[3192]) );
  AND U22694 ( .A(p_input[23192]), .B(p_input[13192]), .Z(n15130) );
  AND U22695 ( .A(p_input[33192]), .B(p_input[3192]), .Z(n15129) );
  AND U22696 ( .A(n15131), .B(n15132), .Z(o[3191]) );
  AND U22697 ( .A(p_input[23191]), .B(p_input[13191]), .Z(n15132) );
  AND U22698 ( .A(p_input[33191]), .B(p_input[3191]), .Z(n15131) );
  AND U22699 ( .A(n15133), .B(n15134), .Z(o[3190]) );
  AND U22700 ( .A(p_input[23190]), .B(p_input[13190]), .Z(n15134) );
  AND U22701 ( .A(p_input[33190]), .B(p_input[3190]), .Z(n15133) );
  AND U22702 ( .A(n15135), .B(n15136), .Z(o[318]) );
  AND U22703 ( .A(p_input[20318]), .B(p_input[10318]), .Z(n15136) );
  AND U22704 ( .A(p_input[318]), .B(p_input[30318]), .Z(n15135) );
  AND U22705 ( .A(n15137), .B(n15138), .Z(o[3189]) );
  AND U22706 ( .A(p_input[23189]), .B(p_input[13189]), .Z(n15138) );
  AND U22707 ( .A(p_input[33189]), .B(p_input[3189]), .Z(n15137) );
  AND U22708 ( .A(n15139), .B(n15140), .Z(o[3188]) );
  AND U22709 ( .A(p_input[23188]), .B(p_input[13188]), .Z(n15140) );
  AND U22710 ( .A(p_input[33188]), .B(p_input[3188]), .Z(n15139) );
  AND U22711 ( .A(n15141), .B(n15142), .Z(o[3187]) );
  AND U22712 ( .A(p_input[23187]), .B(p_input[13187]), .Z(n15142) );
  AND U22713 ( .A(p_input[33187]), .B(p_input[3187]), .Z(n15141) );
  AND U22714 ( .A(n15143), .B(n15144), .Z(o[3186]) );
  AND U22715 ( .A(p_input[23186]), .B(p_input[13186]), .Z(n15144) );
  AND U22716 ( .A(p_input[33186]), .B(p_input[3186]), .Z(n15143) );
  AND U22717 ( .A(n15145), .B(n15146), .Z(o[3185]) );
  AND U22718 ( .A(p_input[23185]), .B(p_input[13185]), .Z(n15146) );
  AND U22719 ( .A(p_input[33185]), .B(p_input[3185]), .Z(n15145) );
  AND U22720 ( .A(n15147), .B(n15148), .Z(o[3184]) );
  AND U22721 ( .A(p_input[23184]), .B(p_input[13184]), .Z(n15148) );
  AND U22722 ( .A(p_input[33184]), .B(p_input[3184]), .Z(n15147) );
  AND U22723 ( .A(n15149), .B(n15150), .Z(o[3183]) );
  AND U22724 ( .A(p_input[23183]), .B(p_input[13183]), .Z(n15150) );
  AND U22725 ( .A(p_input[33183]), .B(p_input[3183]), .Z(n15149) );
  AND U22726 ( .A(n15151), .B(n15152), .Z(o[3182]) );
  AND U22727 ( .A(p_input[23182]), .B(p_input[13182]), .Z(n15152) );
  AND U22728 ( .A(p_input[33182]), .B(p_input[3182]), .Z(n15151) );
  AND U22729 ( .A(n15153), .B(n15154), .Z(o[3181]) );
  AND U22730 ( .A(p_input[23181]), .B(p_input[13181]), .Z(n15154) );
  AND U22731 ( .A(p_input[33181]), .B(p_input[3181]), .Z(n15153) );
  AND U22732 ( .A(n15155), .B(n15156), .Z(o[3180]) );
  AND U22733 ( .A(p_input[23180]), .B(p_input[13180]), .Z(n15156) );
  AND U22734 ( .A(p_input[33180]), .B(p_input[3180]), .Z(n15155) );
  AND U22735 ( .A(n15157), .B(n15158), .Z(o[317]) );
  AND U22736 ( .A(p_input[20317]), .B(p_input[10317]), .Z(n15158) );
  AND U22737 ( .A(p_input[317]), .B(p_input[30317]), .Z(n15157) );
  AND U22738 ( .A(n15159), .B(n15160), .Z(o[3179]) );
  AND U22739 ( .A(p_input[23179]), .B(p_input[13179]), .Z(n15160) );
  AND U22740 ( .A(p_input[33179]), .B(p_input[3179]), .Z(n15159) );
  AND U22741 ( .A(n15161), .B(n15162), .Z(o[3178]) );
  AND U22742 ( .A(p_input[23178]), .B(p_input[13178]), .Z(n15162) );
  AND U22743 ( .A(p_input[33178]), .B(p_input[3178]), .Z(n15161) );
  AND U22744 ( .A(n15163), .B(n15164), .Z(o[3177]) );
  AND U22745 ( .A(p_input[23177]), .B(p_input[13177]), .Z(n15164) );
  AND U22746 ( .A(p_input[33177]), .B(p_input[3177]), .Z(n15163) );
  AND U22747 ( .A(n15165), .B(n15166), .Z(o[3176]) );
  AND U22748 ( .A(p_input[23176]), .B(p_input[13176]), .Z(n15166) );
  AND U22749 ( .A(p_input[33176]), .B(p_input[3176]), .Z(n15165) );
  AND U22750 ( .A(n15167), .B(n15168), .Z(o[3175]) );
  AND U22751 ( .A(p_input[23175]), .B(p_input[13175]), .Z(n15168) );
  AND U22752 ( .A(p_input[33175]), .B(p_input[3175]), .Z(n15167) );
  AND U22753 ( .A(n15169), .B(n15170), .Z(o[3174]) );
  AND U22754 ( .A(p_input[23174]), .B(p_input[13174]), .Z(n15170) );
  AND U22755 ( .A(p_input[33174]), .B(p_input[3174]), .Z(n15169) );
  AND U22756 ( .A(n15171), .B(n15172), .Z(o[3173]) );
  AND U22757 ( .A(p_input[23173]), .B(p_input[13173]), .Z(n15172) );
  AND U22758 ( .A(p_input[33173]), .B(p_input[3173]), .Z(n15171) );
  AND U22759 ( .A(n15173), .B(n15174), .Z(o[3172]) );
  AND U22760 ( .A(p_input[23172]), .B(p_input[13172]), .Z(n15174) );
  AND U22761 ( .A(p_input[33172]), .B(p_input[3172]), .Z(n15173) );
  AND U22762 ( .A(n15175), .B(n15176), .Z(o[3171]) );
  AND U22763 ( .A(p_input[23171]), .B(p_input[13171]), .Z(n15176) );
  AND U22764 ( .A(p_input[33171]), .B(p_input[3171]), .Z(n15175) );
  AND U22765 ( .A(n15177), .B(n15178), .Z(o[3170]) );
  AND U22766 ( .A(p_input[23170]), .B(p_input[13170]), .Z(n15178) );
  AND U22767 ( .A(p_input[33170]), .B(p_input[3170]), .Z(n15177) );
  AND U22768 ( .A(n15179), .B(n15180), .Z(o[316]) );
  AND U22769 ( .A(p_input[20316]), .B(p_input[10316]), .Z(n15180) );
  AND U22770 ( .A(p_input[316]), .B(p_input[30316]), .Z(n15179) );
  AND U22771 ( .A(n15181), .B(n15182), .Z(o[3169]) );
  AND U22772 ( .A(p_input[23169]), .B(p_input[13169]), .Z(n15182) );
  AND U22773 ( .A(p_input[33169]), .B(p_input[3169]), .Z(n15181) );
  AND U22774 ( .A(n15183), .B(n15184), .Z(o[3168]) );
  AND U22775 ( .A(p_input[23168]), .B(p_input[13168]), .Z(n15184) );
  AND U22776 ( .A(p_input[33168]), .B(p_input[3168]), .Z(n15183) );
  AND U22777 ( .A(n15185), .B(n15186), .Z(o[3167]) );
  AND U22778 ( .A(p_input[23167]), .B(p_input[13167]), .Z(n15186) );
  AND U22779 ( .A(p_input[33167]), .B(p_input[3167]), .Z(n15185) );
  AND U22780 ( .A(n15187), .B(n15188), .Z(o[3166]) );
  AND U22781 ( .A(p_input[23166]), .B(p_input[13166]), .Z(n15188) );
  AND U22782 ( .A(p_input[33166]), .B(p_input[3166]), .Z(n15187) );
  AND U22783 ( .A(n15189), .B(n15190), .Z(o[3165]) );
  AND U22784 ( .A(p_input[23165]), .B(p_input[13165]), .Z(n15190) );
  AND U22785 ( .A(p_input[33165]), .B(p_input[3165]), .Z(n15189) );
  AND U22786 ( .A(n15191), .B(n15192), .Z(o[3164]) );
  AND U22787 ( .A(p_input[23164]), .B(p_input[13164]), .Z(n15192) );
  AND U22788 ( .A(p_input[33164]), .B(p_input[3164]), .Z(n15191) );
  AND U22789 ( .A(n15193), .B(n15194), .Z(o[3163]) );
  AND U22790 ( .A(p_input[23163]), .B(p_input[13163]), .Z(n15194) );
  AND U22791 ( .A(p_input[33163]), .B(p_input[3163]), .Z(n15193) );
  AND U22792 ( .A(n15195), .B(n15196), .Z(o[3162]) );
  AND U22793 ( .A(p_input[23162]), .B(p_input[13162]), .Z(n15196) );
  AND U22794 ( .A(p_input[33162]), .B(p_input[3162]), .Z(n15195) );
  AND U22795 ( .A(n15197), .B(n15198), .Z(o[3161]) );
  AND U22796 ( .A(p_input[23161]), .B(p_input[13161]), .Z(n15198) );
  AND U22797 ( .A(p_input[33161]), .B(p_input[3161]), .Z(n15197) );
  AND U22798 ( .A(n15199), .B(n15200), .Z(o[3160]) );
  AND U22799 ( .A(p_input[23160]), .B(p_input[13160]), .Z(n15200) );
  AND U22800 ( .A(p_input[33160]), .B(p_input[3160]), .Z(n15199) );
  AND U22801 ( .A(n15201), .B(n15202), .Z(o[315]) );
  AND U22802 ( .A(p_input[20315]), .B(p_input[10315]), .Z(n15202) );
  AND U22803 ( .A(p_input[315]), .B(p_input[30315]), .Z(n15201) );
  AND U22804 ( .A(n15203), .B(n15204), .Z(o[3159]) );
  AND U22805 ( .A(p_input[23159]), .B(p_input[13159]), .Z(n15204) );
  AND U22806 ( .A(p_input[33159]), .B(p_input[3159]), .Z(n15203) );
  AND U22807 ( .A(n15205), .B(n15206), .Z(o[3158]) );
  AND U22808 ( .A(p_input[23158]), .B(p_input[13158]), .Z(n15206) );
  AND U22809 ( .A(p_input[33158]), .B(p_input[3158]), .Z(n15205) );
  AND U22810 ( .A(n15207), .B(n15208), .Z(o[3157]) );
  AND U22811 ( .A(p_input[23157]), .B(p_input[13157]), .Z(n15208) );
  AND U22812 ( .A(p_input[33157]), .B(p_input[3157]), .Z(n15207) );
  AND U22813 ( .A(n15209), .B(n15210), .Z(o[3156]) );
  AND U22814 ( .A(p_input[23156]), .B(p_input[13156]), .Z(n15210) );
  AND U22815 ( .A(p_input[33156]), .B(p_input[3156]), .Z(n15209) );
  AND U22816 ( .A(n15211), .B(n15212), .Z(o[3155]) );
  AND U22817 ( .A(p_input[23155]), .B(p_input[13155]), .Z(n15212) );
  AND U22818 ( .A(p_input[33155]), .B(p_input[3155]), .Z(n15211) );
  AND U22819 ( .A(n15213), .B(n15214), .Z(o[3154]) );
  AND U22820 ( .A(p_input[23154]), .B(p_input[13154]), .Z(n15214) );
  AND U22821 ( .A(p_input[33154]), .B(p_input[3154]), .Z(n15213) );
  AND U22822 ( .A(n15215), .B(n15216), .Z(o[3153]) );
  AND U22823 ( .A(p_input[23153]), .B(p_input[13153]), .Z(n15216) );
  AND U22824 ( .A(p_input[33153]), .B(p_input[3153]), .Z(n15215) );
  AND U22825 ( .A(n15217), .B(n15218), .Z(o[3152]) );
  AND U22826 ( .A(p_input[23152]), .B(p_input[13152]), .Z(n15218) );
  AND U22827 ( .A(p_input[33152]), .B(p_input[3152]), .Z(n15217) );
  AND U22828 ( .A(n15219), .B(n15220), .Z(o[3151]) );
  AND U22829 ( .A(p_input[23151]), .B(p_input[13151]), .Z(n15220) );
  AND U22830 ( .A(p_input[33151]), .B(p_input[3151]), .Z(n15219) );
  AND U22831 ( .A(n15221), .B(n15222), .Z(o[3150]) );
  AND U22832 ( .A(p_input[23150]), .B(p_input[13150]), .Z(n15222) );
  AND U22833 ( .A(p_input[33150]), .B(p_input[3150]), .Z(n15221) );
  AND U22834 ( .A(n15223), .B(n15224), .Z(o[314]) );
  AND U22835 ( .A(p_input[20314]), .B(p_input[10314]), .Z(n15224) );
  AND U22836 ( .A(p_input[314]), .B(p_input[30314]), .Z(n15223) );
  AND U22837 ( .A(n15225), .B(n15226), .Z(o[3149]) );
  AND U22838 ( .A(p_input[23149]), .B(p_input[13149]), .Z(n15226) );
  AND U22839 ( .A(p_input[33149]), .B(p_input[3149]), .Z(n15225) );
  AND U22840 ( .A(n15227), .B(n15228), .Z(o[3148]) );
  AND U22841 ( .A(p_input[23148]), .B(p_input[13148]), .Z(n15228) );
  AND U22842 ( .A(p_input[33148]), .B(p_input[3148]), .Z(n15227) );
  AND U22843 ( .A(n15229), .B(n15230), .Z(o[3147]) );
  AND U22844 ( .A(p_input[23147]), .B(p_input[13147]), .Z(n15230) );
  AND U22845 ( .A(p_input[33147]), .B(p_input[3147]), .Z(n15229) );
  AND U22846 ( .A(n15231), .B(n15232), .Z(o[3146]) );
  AND U22847 ( .A(p_input[23146]), .B(p_input[13146]), .Z(n15232) );
  AND U22848 ( .A(p_input[33146]), .B(p_input[3146]), .Z(n15231) );
  AND U22849 ( .A(n15233), .B(n15234), .Z(o[3145]) );
  AND U22850 ( .A(p_input[23145]), .B(p_input[13145]), .Z(n15234) );
  AND U22851 ( .A(p_input[33145]), .B(p_input[3145]), .Z(n15233) );
  AND U22852 ( .A(n15235), .B(n15236), .Z(o[3144]) );
  AND U22853 ( .A(p_input[23144]), .B(p_input[13144]), .Z(n15236) );
  AND U22854 ( .A(p_input[33144]), .B(p_input[3144]), .Z(n15235) );
  AND U22855 ( .A(n15237), .B(n15238), .Z(o[3143]) );
  AND U22856 ( .A(p_input[23143]), .B(p_input[13143]), .Z(n15238) );
  AND U22857 ( .A(p_input[33143]), .B(p_input[3143]), .Z(n15237) );
  AND U22858 ( .A(n15239), .B(n15240), .Z(o[3142]) );
  AND U22859 ( .A(p_input[23142]), .B(p_input[13142]), .Z(n15240) );
  AND U22860 ( .A(p_input[33142]), .B(p_input[3142]), .Z(n15239) );
  AND U22861 ( .A(n15241), .B(n15242), .Z(o[3141]) );
  AND U22862 ( .A(p_input[23141]), .B(p_input[13141]), .Z(n15242) );
  AND U22863 ( .A(p_input[33141]), .B(p_input[3141]), .Z(n15241) );
  AND U22864 ( .A(n15243), .B(n15244), .Z(o[3140]) );
  AND U22865 ( .A(p_input[23140]), .B(p_input[13140]), .Z(n15244) );
  AND U22866 ( .A(p_input[33140]), .B(p_input[3140]), .Z(n15243) );
  AND U22867 ( .A(n15245), .B(n15246), .Z(o[313]) );
  AND U22868 ( .A(p_input[20313]), .B(p_input[10313]), .Z(n15246) );
  AND U22869 ( .A(p_input[313]), .B(p_input[30313]), .Z(n15245) );
  AND U22870 ( .A(n15247), .B(n15248), .Z(o[3139]) );
  AND U22871 ( .A(p_input[23139]), .B(p_input[13139]), .Z(n15248) );
  AND U22872 ( .A(p_input[33139]), .B(p_input[3139]), .Z(n15247) );
  AND U22873 ( .A(n15249), .B(n15250), .Z(o[3138]) );
  AND U22874 ( .A(p_input[23138]), .B(p_input[13138]), .Z(n15250) );
  AND U22875 ( .A(p_input[33138]), .B(p_input[3138]), .Z(n15249) );
  AND U22876 ( .A(n15251), .B(n15252), .Z(o[3137]) );
  AND U22877 ( .A(p_input[23137]), .B(p_input[13137]), .Z(n15252) );
  AND U22878 ( .A(p_input[33137]), .B(p_input[3137]), .Z(n15251) );
  AND U22879 ( .A(n15253), .B(n15254), .Z(o[3136]) );
  AND U22880 ( .A(p_input[23136]), .B(p_input[13136]), .Z(n15254) );
  AND U22881 ( .A(p_input[33136]), .B(p_input[3136]), .Z(n15253) );
  AND U22882 ( .A(n15255), .B(n15256), .Z(o[3135]) );
  AND U22883 ( .A(p_input[23135]), .B(p_input[13135]), .Z(n15256) );
  AND U22884 ( .A(p_input[33135]), .B(p_input[3135]), .Z(n15255) );
  AND U22885 ( .A(n15257), .B(n15258), .Z(o[3134]) );
  AND U22886 ( .A(p_input[23134]), .B(p_input[13134]), .Z(n15258) );
  AND U22887 ( .A(p_input[33134]), .B(p_input[3134]), .Z(n15257) );
  AND U22888 ( .A(n15259), .B(n15260), .Z(o[3133]) );
  AND U22889 ( .A(p_input[23133]), .B(p_input[13133]), .Z(n15260) );
  AND U22890 ( .A(p_input[33133]), .B(p_input[3133]), .Z(n15259) );
  AND U22891 ( .A(n15261), .B(n15262), .Z(o[3132]) );
  AND U22892 ( .A(p_input[23132]), .B(p_input[13132]), .Z(n15262) );
  AND U22893 ( .A(p_input[33132]), .B(p_input[3132]), .Z(n15261) );
  AND U22894 ( .A(n15263), .B(n15264), .Z(o[3131]) );
  AND U22895 ( .A(p_input[23131]), .B(p_input[13131]), .Z(n15264) );
  AND U22896 ( .A(p_input[33131]), .B(p_input[3131]), .Z(n15263) );
  AND U22897 ( .A(n15265), .B(n15266), .Z(o[3130]) );
  AND U22898 ( .A(p_input[23130]), .B(p_input[13130]), .Z(n15266) );
  AND U22899 ( .A(p_input[33130]), .B(p_input[3130]), .Z(n15265) );
  AND U22900 ( .A(n15267), .B(n15268), .Z(o[312]) );
  AND U22901 ( .A(p_input[20312]), .B(p_input[10312]), .Z(n15268) );
  AND U22902 ( .A(p_input[312]), .B(p_input[30312]), .Z(n15267) );
  AND U22903 ( .A(n15269), .B(n15270), .Z(o[3129]) );
  AND U22904 ( .A(p_input[23129]), .B(p_input[13129]), .Z(n15270) );
  AND U22905 ( .A(p_input[33129]), .B(p_input[3129]), .Z(n15269) );
  AND U22906 ( .A(n15271), .B(n15272), .Z(o[3128]) );
  AND U22907 ( .A(p_input[23128]), .B(p_input[13128]), .Z(n15272) );
  AND U22908 ( .A(p_input[33128]), .B(p_input[3128]), .Z(n15271) );
  AND U22909 ( .A(n15273), .B(n15274), .Z(o[3127]) );
  AND U22910 ( .A(p_input[23127]), .B(p_input[13127]), .Z(n15274) );
  AND U22911 ( .A(p_input[33127]), .B(p_input[3127]), .Z(n15273) );
  AND U22912 ( .A(n15275), .B(n15276), .Z(o[3126]) );
  AND U22913 ( .A(p_input[23126]), .B(p_input[13126]), .Z(n15276) );
  AND U22914 ( .A(p_input[33126]), .B(p_input[3126]), .Z(n15275) );
  AND U22915 ( .A(n15277), .B(n15278), .Z(o[3125]) );
  AND U22916 ( .A(p_input[23125]), .B(p_input[13125]), .Z(n15278) );
  AND U22917 ( .A(p_input[33125]), .B(p_input[3125]), .Z(n15277) );
  AND U22918 ( .A(n15279), .B(n15280), .Z(o[3124]) );
  AND U22919 ( .A(p_input[23124]), .B(p_input[13124]), .Z(n15280) );
  AND U22920 ( .A(p_input[33124]), .B(p_input[3124]), .Z(n15279) );
  AND U22921 ( .A(n15281), .B(n15282), .Z(o[3123]) );
  AND U22922 ( .A(p_input[23123]), .B(p_input[13123]), .Z(n15282) );
  AND U22923 ( .A(p_input[33123]), .B(p_input[3123]), .Z(n15281) );
  AND U22924 ( .A(n15283), .B(n15284), .Z(o[3122]) );
  AND U22925 ( .A(p_input[23122]), .B(p_input[13122]), .Z(n15284) );
  AND U22926 ( .A(p_input[33122]), .B(p_input[3122]), .Z(n15283) );
  AND U22927 ( .A(n15285), .B(n15286), .Z(o[3121]) );
  AND U22928 ( .A(p_input[23121]), .B(p_input[13121]), .Z(n15286) );
  AND U22929 ( .A(p_input[33121]), .B(p_input[3121]), .Z(n15285) );
  AND U22930 ( .A(n15287), .B(n15288), .Z(o[3120]) );
  AND U22931 ( .A(p_input[23120]), .B(p_input[13120]), .Z(n15288) );
  AND U22932 ( .A(p_input[33120]), .B(p_input[3120]), .Z(n15287) );
  AND U22933 ( .A(n15289), .B(n15290), .Z(o[311]) );
  AND U22934 ( .A(p_input[20311]), .B(p_input[10311]), .Z(n15290) );
  AND U22935 ( .A(p_input[311]), .B(p_input[30311]), .Z(n15289) );
  AND U22936 ( .A(n15291), .B(n15292), .Z(o[3119]) );
  AND U22937 ( .A(p_input[23119]), .B(p_input[13119]), .Z(n15292) );
  AND U22938 ( .A(p_input[33119]), .B(p_input[3119]), .Z(n15291) );
  AND U22939 ( .A(n15293), .B(n15294), .Z(o[3118]) );
  AND U22940 ( .A(p_input[23118]), .B(p_input[13118]), .Z(n15294) );
  AND U22941 ( .A(p_input[33118]), .B(p_input[3118]), .Z(n15293) );
  AND U22942 ( .A(n15295), .B(n15296), .Z(o[3117]) );
  AND U22943 ( .A(p_input[23117]), .B(p_input[13117]), .Z(n15296) );
  AND U22944 ( .A(p_input[33117]), .B(p_input[3117]), .Z(n15295) );
  AND U22945 ( .A(n15297), .B(n15298), .Z(o[3116]) );
  AND U22946 ( .A(p_input[23116]), .B(p_input[13116]), .Z(n15298) );
  AND U22947 ( .A(p_input[33116]), .B(p_input[3116]), .Z(n15297) );
  AND U22948 ( .A(n15299), .B(n15300), .Z(o[3115]) );
  AND U22949 ( .A(p_input[23115]), .B(p_input[13115]), .Z(n15300) );
  AND U22950 ( .A(p_input[33115]), .B(p_input[3115]), .Z(n15299) );
  AND U22951 ( .A(n15301), .B(n15302), .Z(o[3114]) );
  AND U22952 ( .A(p_input[23114]), .B(p_input[13114]), .Z(n15302) );
  AND U22953 ( .A(p_input[33114]), .B(p_input[3114]), .Z(n15301) );
  AND U22954 ( .A(n15303), .B(n15304), .Z(o[3113]) );
  AND U22955 ( .A(p_input[23113]), .B(p_input[13113]), .Z(n15304) );
  AND U22956 ( .A(p_input[33113]), .B(p_input[3113]), .Z(n15303) );
  AND U22957 ( .A(n15305), .B(n15306), .Z(o[3112]) );
  AND U22958 ( .A(p_input[23112]), .B(p_input[13112]), .Z(n15306) );
  AND U22959 ( .A(p_input[33112]), .B(p_input[3112]), .Z(n15305) );
  AND U22960 ( .A(n15307), .B(n15308), .Z(o[3111]) );
  AND U22961 ( .A(p_input[23111]), .B(p_input[13111]), .Z(n15308) );
  AND U22962 ( .A(p_input[33111]), .B(p_input[3111]), .Z(n15307) );
  AND U22963 ( .A(n15309), .B(n15310), .Z(o[3110]) );
  AND U22964 ( .A(p_input[23110]), .B(p_input[13110]), .Z(n15310) );
  AND U22965 ( .A(p_input[33110]), .B(p_input[3110]), .Z(n15309) );
  AND U22966 ( .A(n15311), .B(n15312), .Z(o[310]) );
  AND U22967 ( .A(p_input[20310]), .B(p_input[10310]), .Z(n15312) );
  AND U22968 ( .A(p_input[310]), .B(p_input[30310]), .Z(n15311) );
  AND U22969 ( .A(n15313), .B(n15314), .Z(o[3109]) );
  AND U22970 ( .A(p_input[23109]), .B(p_input[13109]), .Z(n15314) );
  AND U22971 ( .A(p_input[33109]), .B(p_input[3109]), .Z(n15313) );
  AND U22972 ( .A(n15315), .B(n15316), .Z(o[3108]) );
  AND U22973 ( .A(p_input[23108]), .B(p_input[13108]), .Z(n15316) );
  AND U22974 ( .A(p_input[33108]), .B(p_input[3108]), .Z(n15315) );
  AND U22975 ( .A(n15317), .B(n15318), .Z(o[3107]) );
  AND U22976 ( .A(p_input[23107]), .B(p_input[13107]), .Z(n15318) );
  AND U22977 ( .A(p_input[33107]), .B(p_input[3107]), .Z(n15317) );
  AND U22978 ( .A(n15319), .B(n15320), .Z(o[3106]) );
  AND U22979 ( .A(p_input[23106]), .B(p_input[13106]), .Z(n15320) );
  AND U22980 ( .A(p_input[33106]), .B(p_input[3106]), .Z(n15319) );
  AND U22981 ( .A(n15321), .B(n15322), .Z(o[3105]) );
  AND U22982 ( .A(p_input[23105]), .B(p_input[13105]), .Z(n15322) );
  AND U22983 ( .A(p_input[33105]), .B(p_input[3105]), .Z(n15321) );
  AND U22984 ( .A(n15323), .B(n15324), .Z(o[3104]) );
  AND U22985 ( .A(p_input[23104]), .B(p_input[13104]), .Z(n15324) );
  AND U22986 ( .A(p_input[33104]), .B(p_input[3104]), .Z(n15323) );
  AND U22987 ( .A(n15325), .B(n15326), .Z(o[3103]) );
  AND U22988 ( .A(p_input[23103]), .B(p_input[13103]), .Z(n15326) );
  AND U22989 ( .A(p_input[33103]), .B(p_input[3103]), .Z(n15325) );
  AND U22990 ( .A(n15327), .B(n15328), .Z(o[3102]) );
  AND U22991 ( .A(p_input[23102]), .B(p_input[13102]), .Z(n15328) );
  AND U22992 ( .A(p_input[33102]), .B(p_input[3102]), .Z(n15327) );
  AND U22993 ( .A(n15329), .B(n15330), .Z(o[3101]) );
  AND U22994 ( .A(p_input[23101]), .B(p_input[13101]), .Z(n15330) );
  AND U22995 ( .A(p_input[33101]), .B(p_input[3101]), .Z(n15329) );
  AND U22996 ( .A(n15331), .B(n15332), .Z(o[3100]) );
  AND U22997 ( .A(p_input[23100]), .B(p_input[13100]), .Z(n15332) );
  AND U22998 ( .A(p_input[33100]), .B(p_input[3100]), .Z(n15331) );
  AND U22999 ( .A(n15333), .B(n15334), .Z(o[30]) );
  AND U23000 ( .A(p_input[20030]), .B(p_input[10030]), .Z(n15334) );
  AND U23001 ( .A(p_input[30]), .B(p_input[30030]), .Z(n15333) );
  AND U23002 ( .A(n15335), .B(n15336), .Z(o[309]) );
  AND U23003 ( .A(p_input[20309]), .B(p_input[10309]), .Z(n15336) );
  AND U23004 ( .A(p_input[309]), .B(p_input[30309]), .Z(n15335) );
  AND U23005 ( .A(n15337), .B(n15338), .Z(o[3099]) );
  AND U23006 ( .A(p_input[23099]), .B(p_input[13099]), .Z(n15338) );
  AND U23007 ( .A(p_input[33099]), .B(p_input[3099]), .Z(n15337) );
  AND U23008 ( .A(n15339), .B(n15340), .Z(o[3098]) );
  AND U23009 ( .A(p_input[23098]), .B(p_input[13098]), .Z(n15340) );
  AND U23010 ( .A(p_input[33098]), .B(p_input[3098]), .Z(n15339) );
  AND U23011 ( .A(n15341), .B(n15342), .Z(o[3097]) );
  AND U23012 ( .A(p_input[23097]), .B(p_input[13097]), .Z(n15342) );
  AND U23013 ( .A(p_input[33097]), .B(p_input[3097]), .Z(n15341) );
  AND U23014 ( .A(n15343), .B(n15344), .Z(o[3096]) );
  AND U23015 ( .A(p_input[23096]), .B(p_input[13096]), .Z(n15344) );
  AND U23016 ( .A(p_input[33096]), .B(p_input[3096]), .Z(n15343) );
  AND U23017 ( .A(n15345), .B(n15346), .Z(o[3095]) );
  AND U23018 ( .A(p_input[23095]), .B(p_input[13095]), .Z(n15346) );
  AND U23019 ( .A(p_input[33095]), .B(p_input[3095]), .Z(n15345) );
  AND U23020 ( .A(n15347), .B(n15348), .Z(o[3094]) );
  AND U23021 ( .A(p_input[23094]), .B(p_input[13094]), .Z(n15348) );
  AND U23022 ( .A(p_input[33094]), .B(p_input[3094]), .Z(n15347) );
  AND U23023 ( .A(n15349), .B(n15350), .Z(o[3093]) );
  AND U23024 ( .A(p_input[23093]), .B(p_input[13093]), .Z(n15350) );
  AND U23025 ( .A(p_input[33093]), .B(p_input[3093]), .Z(n15349) );
  AND U23026 ( .A(n15351), .B(n15352), .Z(o[3092]) );
  AND U23027 ( .A(p_input[23092]), .B(p_input[13092]), .Z(n15352) );
  AND U23028 ( .A(p_input[33092]), .B(p_input[3092]), .Z(n15351) );
  AND U23029 ( .A(n15353), .B(n15354), .Z(o[3091]) );
  AND U23030 ( .A(p_input[23091]), .B(p_input[13091]), .Z(n15354) );
  AND U23031 ( .A(p_input[33091]), .B(p_input[3091]), .Z(n15353) );
  AND U23032 ( .A(n15355), .B(n15356), .Z(o[3090]) );
  AND U23033 ( .A(p_input[23090]), .B(p_input[13090]), .Z(n15356) );
  AND U23034 ( .A(p_input[33090]), .B(p_input[3090]), .Z(n15355) );
  AND U23035 ( .A(n15357), .B(n15358), .Z(o[308]) );
  AND U23036 ( .A(p_input[20308]), .B(p_input[10308]), .Z(n15358) );
  AND U23037 ( .A(p_input[308]), .B(p_input[30308]), .Z(n15357) );
  AND U23038 ( .A(n15359), .B(n15360), .Z(o[3089]) );
  AND U23039 ( .A(p_input[23089]), .B(p_input[13089]), .Z(n15360) );
  AND U23040 ( .A(p_input[33089]), .B(p_input[3089]), .Z(n15359) );
  AND U23041 ( .A(n15361), .B(n15362), .Z(o[3088]) );
  AND U23042 ( .A(p_input[23088]), .B(p_input[13088]), .Z(n15362) );
  AND U23043 ( .A(p_input[33088]), .B(p_input[3088]), .Z(n15361) );
  AND U23044 ( .A(n15363), .B(n15364), .Z(o[3087]) );
  AND U23045 ( .A(p_input[23087]), .B(p_input[13087]), .Z(n15364) );
  AND U23046 ( .A(p_input[33087]), .B(p_input[3087]), .Z(n15363) );
  AND U23047 ( .A(n15365), .B(n15366), .Z(o[3086]) );
  AND U23048 ( .A(p_input[23086]), .B(p_input[13086]), .Z(n15366) );
  AND U23049 ( .A(p_input[33086]), .B(p_input[3086]), .Z(n15365) );
  AND U23050 ( .A(n15367), .B(n15368), .Z(o[3085]) );
  AND U23051 ( .A(p_input[23085]), .B(p_input[13085]), .Z(n15368) );
  AND U23052 ( .A(p_input[33085]), .B(p_input[3085]), .Z(n15367) );
  AND U23053 ( .A(n15369), .B(n15370), .Z(o[3084]) );
  AND U23054 ( .A(p_input[23084]), .B(p_input[13084]), .Z(n15370) );
  AND U23055 ( .A(p_input[33084]), .B(p_input[3084]), .Z(n15369) );
  AND U23056 ( .A(n15371), .B(n15372), .Z(o[3083]) );
  AND U23057 ( .A(p_input[23083]), .B(p_input[13083]), .Z(n15372) );
  AND U23058 ( .A(p_input[33083]), .B(p_input[3083]), .Z(n15371) );
  AND U23059 ( .A(n15373), .B(n15374), .Z(o[3082]) );
  AND U23060 ( .A(p_input[23082]), .B(p_input[13082]), .Z(n15374) );
  AND U23061 ( .A(p_input[33082]), .B(p_input[3082]), .Z(n15373) );
  AND U23062 ( .A(n15375), .B(n15376), .Z(o[3081]) );
  AND U23063 ( .A(p_input[23081]), .B(p_input[13081]), .Z(n15376) );
  AND U23064 ( .A(p_input[33081]), .B(p_input[3081]), .Z(n15375) );
  AND U23065 ( .A(n15377), .B(n15378), .Z(o[3080]) );
  AND U23066 ( .A(p_input[23080]), .B(p_input[13080]), .Z(n15378) );
  AND U23067 ( .A(p_input[33080]), .B(p_input[3080]), .Z(n15377) );
  AND U23068 ( .A(n15379), .B(n15380), .Z(o[307]) );
  AND U23069 ( .A(p_input[20307]), .B(p_input[10307]), .Z(n15380) );
  AND U23070 ( .A(p_input[307]), .B(p_input[30307]), .Z(n15379) );
  AND U23071 ( .A(n15381), .B(n15382), .Z(o[3079]) );
  AND U23072 ( .A(p_input[23079]), .B(p_input[13079]), .Z(n15382) );
  AND U23073 ( .A(p_input[33079]), .B(p_input[3079]), .Z(n15381) );
  AND U23074 ( .A(n15383), .B(n15384), .Z(o[3078]) );
  AND U23075 ( .A(p_input[23078]), .B(p_input[13078]), .Z(n15384) );
  AND U23076 ( .A(p_input[33078]), .B(p_input[3078]), .Z(n15383) );
  AND U23077 ( .A(n15385), .B(n15386), .Z(o[3077]) );
  AND U23078 ( .A(p_input[23077]), .B(p_input[13077]), .Z(n15386) );
  AND U23079 ( .A(p_input[33077]), .B(p_input[3077]), .Z(n15385) );
  AND U23080 ( .A(n15387), .B(n15388), .Z(o[3076]) );
  AND U23081 ( .A(p_input[23076]), .B(p_input[13076]), .Z(n15388) );
  AND U23082 ( .A(p_input[33076]), .B(p_input[3076]), .Z(n15387) );
  AND U23083 ( .A(n15389), .B(n15390), .Z(o[3075]) );
  AND U23084 ( .A(p_input[23075]), .B(p_input[13075]), .Z(n15390) );
  AND U23085 ( .A(p_input[33075]), .B(p_input[3075]), .Z(n15389) );
  AND U23086 ( .A(n15391), .B(n15392), .Z(o[3074]) );
  AND U23087 ( .A(p_input[23074]), .B(p_input[13074]), .Z(n15392) );
  AND U23088 ( .A(p_input[33074]), .B(p_input[3074]), .Z(n15391) );
  AND U23089 ( .A(n15393), .B(n15394), .Z(o[3073]) );
  AND U23090 ( .A(p_input[23073]), .B(p_input[13073]), .Z(n15394) );
  AND U23091 ( .A(p_input[33073]), .B(p_input[3073]), .Z(n15393) );
  AND U23092 ( .A(n15395), .B(n15396), .Z(o[3072]) );
  AND U23093 ( .A(p_input[23072]), .B(p_input[13072]), .Z(n15396) );
  AND U23094 ( .A(p_input[33072]), .B(p_input[3072]), .Z(n15395) );
  AND U23095 ( .A(n15397), .B(n15398), .Z(o[3071]) );
  AND U23096 ( .A(p_input[23071]), .B(p_input[13071]), .Z(n15398) );
  AND U23097 ( .A(p_input[33071]), .B(p_input[3071]), .Z(n15397) );
  AND U23098 ( .A(n15399), .B(n15400), .Z(o[3070]) );
  AND U23099 ( .A(p_input[23070]), .B(p_input[13070]), .Z(n15400) );
  AND U23100 ( .A(p_input[33070]), .B(p_input[3070]), .Z(n15399) );
  AND U23101 ( .A(n15401), .B(n15402), .Z(o[306]) );
  AND U23102 ( .A(p_input[20306]), .B(p_input[10306]), .Z(n15402) );
  AND U23103 ( .A(p_input[306]), .B(p_input[30306]), .Z(n15401) );
  AND U23104 ( .A(n15403), .B(n15404), .Z(o[3069]) );
  AND U23105 ( .A(p_input[23069]), .B(p_input[13069]), .Z(n15404) );
  AND U23106 ( .A(p_input[33069]), .B(p_input[3069]), .Z(n15403) );
  AND U23107 ( .A(n15405), .B(n15406), .Z(o[3068]) );
  AND U23108 ( .A(p_input[23068]), .B(p_input[13068]), .Z(n15406) );
  AND U23109 ( .A(p_input[33068]), .B(p_input[3068]), .Z(n15405) );
  AND U23110 ( .A(n15407), .B(n15408), .Z(o[3067]) );
  AND U23111 ( .A(p_input[23067]), .B(p_input[13067]), .Z(n15408) );
  AND U23112 ( .A(p_input[33067]), .B(p_input[3067]), .Z(n15407) );
  AND U23113 ( .A(n15409), .B(n15410), .Z(o[3066]) );
  AND U23114 ( .A(p_input[23066]), .B(p_input[13066]), .Z(n15410) );
  AND U23115 ( .A(p_input[33066]), .B(p_input[3066]), .Z(n15409) );
  AND U23116 ( .A(n15411), .B(n15412), .Z(o[3065]) );
  AND U23117 ( .A(p_input[23065]), .B(p_input[13065]), .Z(n15412) );
  AND U23118 ( .A(p_input[33065]), .B(p_input[3065]), .Z(n15411) );
  AND U23119 ( .A(n15413), .B(n15414), .Z(o[3064]) );
  AND U23120 ( .A(p_input[23064]), .B(p_input[13064]), .Z(n15414) );
  AND U23121 ( .A(p_input[33064]), .B(p_input[3064]), .Z(n15413) );
  AND U23122 ( .A(n15415), .B(n15416), .Z(o[3063]) );
  AND U23123 ( .A(p_input[23063]), .B(p_input[13063]), .Z(n15416) );
  AND U23124 ( .A(p_input[33063]), .B(p_input[3063]), .Z(n15415) );
  AND U23125 ( .A(n15417), .B(n15418), .Z(o[3062]) );
  AND U23126 ( .A(p_input[23062]), .B(p_input[13062]), .Z(n15418) );
  AND U23127 ( .A(p_input[33062]), .B(p_input[3062]), .Z(n15417) );
  AND U23128 ( .A(n15419), .B(n15420), .Z(o[3061]) );
  AND U23129 ( .A(p_input[23061]), .B(p_input[13061]), .Z(n15420) );
  AND U23130 ( .A(p_input[33061]), .B(p_input[3061]), .Z(n15419) );
  AND U23131 ( .A(n15421), .B(n15422), .Z(o[3060]) );
  AND U23132 ( .A(p_input[23060]), .B(p_input[13060]), .Z(n15422) );
  AND U23133 ( .A(p_input[33060]), .B(p_input[3060]), .Z(n15421) );
  AND U23134 ( .A(n15423), .B(n15424), .Z(o[305]) );
  AND U23135 ( .A(p_input[20305]), .B(p_input[10305]), .Z(n15424) );
  AND U23136 ( .A(p_input[305]), .B(p_input[30305]), .Z(n15423) );
  AND U23137 ( .A(n15425), .B(n15426), .Z(o[3059]) );
  AND U23138 ( .A(p_input[23059]), .B(p_input[13059]), .Z(n15426) );
  AND U23139 ( .A(p_input[33059]), .B(p_input[3059]), .Z(n15425) );
  AND U23140 ( .A(n15427), .B(n15428), .Z(o[3058]) );
  AND U23141 ( .A(p_input[23058]), .B(p_input[13058]), .Z(n15428) );
  AND U23142 ( .A(p_input[33058]), .B(p_input[3058]), .Z(n15427) );
  AND U23143 ( .A(n15429), .B(n15430), .Z(o[3057]) );
  AND U23144 ( .A(p_input[23057]), .B(p_input[13057]), .Z(n15430) );
  AND U23145 ( .A(p_input[33057]), .B(p_input[3057]), .Z(n15429) );
  AND U23146 ( .A(n15431), .B(n15432), .Z(o[3056]) );
  AND U23147 ( .A(p_input[23056]), .B(p_input[13056]), .Z(n15432) );
  AND U23148 ( .A(p_input[33056]), .B(p_input[3056]), .Z(n15431) );
  AND U23149 ( .A(n15433), .B(n15434), .Z(o[3055]) );
  AND U23150 ( .A(p_input[23055]), .B(p_input[13055]), .Z(n15434) );
  AND U23151 ( .A(p_input[33055]), .B(p_input[3055]), .Z(n15433) );
  AND U23152 ( .A(n15435), .B(n15436), .Z(o[3054]) );
  AND U23153 ( .A(p_input[23054]), .B(p_input[13054]), .Z(n15436) );
  AND U23154 ( .A(p_input[33054]), .B(p_input[3054]), .Z(n15435) );
  AND U23155 ( .A(n15437), .B(n15438), .Z(o[3053]) );
  AND U23156 ( .A(p_input[23053]), .B(p_input[13053]), .Z(n15438) );
  AND U23157 ( .A(p_input[33053]), .B(p_input[3053]), .Z(n15437) );
  AND U23158 ( .A(n15439), .B(n15440), .Z(o[3052]) );
  AND U23159 ( .A(p_input[23052]), .B(p_input[13052]), .Z(n15440) );
  AND U23160 ( .A(p_input[33052]), .B(p_input[3052]), .Z(n15439) );
  AND U23161 ( .A(n15441), .B(n15442), .Z(o[3051]) );
  AND U23162 ( .A(p_input[23051]), .B(p_input[13051]), .Z(n15442) );
  AND U23163 ( .A(p_input[33051]), .B(p_input[3051]), .Z(n15441) );
  AND U23164 ( .A(n15443), .B(n15444), .Z(o[3050]) );
  AND U23165 ( .A(p_input[23050]), .B(p_input[13050]), .Z(n15444) );
  AND U23166 ( .A(p_input[33050]), .B(p_input[3050]), .Z(n15443) );
  AND U23167 ( .A(n15445), .B(n15446), .Z(o[304]) );
  AND U23168 ( .A(p_input[20304]), .B(p_input[10304]), .Z(n15446) );
  AND U23169 ( .A(p_input[304]), .B(p_input[30304]), .Z(n15445) );
  AND U23170 ( .A(n15447), .B(n15448), .Z(o[3049]) );
  AND U23171 ( .A(p_input[23049]), .B(p_input[13049]), .Z(n15448) );
  AND U23172 ( .A(p_input[33049]), .B(p_input[3049]), .Z(n15447) );
  AND U23173 ( .A(n15449), .B(n15450), .Z(o[3048]) );
  AND U23174 ( .A(p_input[23048]), .B(p_input[13048]), .Z(n15450) );
  AND U23175 ( .A(p_input[33048]), .B(p_input[3048]), .Z(n15449) );
  AND U23176 ( .A(n15451), .B(n15452), .Z(o[3047]) );
  AND U23177 ( .A(p_input[23047]), .B(p_input[13047]), .Z(n15452) );
  AND U23178 ( .A(p_input[33047]), .B(p_input[3047]), .Z(n15451) );
  AND U23179 ( .A(n15453), .B(n15454), .Z(o[3046]) );
  AND U23180 ( .A(p_input[23046]), .B(p_input[13046]), .Z(n15454) );
  AND U23181 ( .A(p_input[33046]), .B(p_input[3046]), .Z(n15453) );
  AND U23182 ( .A(n15455), .B(n15456), .Z(o[3045]) );
  AND U23183 ( .A(p_input[23045]), .B(p_input[13045]), .Z(n15456) );
  AND U23184 ( .A(p_input[33045]), .B(p_input[3045]), .Z(n15455) );
  AND U23185 ( .A(n15457), .B(n15458), .Z(o[3044]) );
  AND U23186 ( .A(p_input[23044]), .B(p_input[13044]), .Z(n15458) );
  AND U23187 ( .A(p_input[33044]), .B(p_input[3044]), .Z(n15457) );
  AND U23188 ( .A(n15459), .B(n15460), .Z(o[3043]) );
  AND U23189 ( .A(p_input[23043]), .B(p_input[13043]), .Z(n15460) );
  AND U23190 ( .A(p_input[33043]), .B(p_input[3043]), .Z(n15459) );
  AND U23191 ( .A(n15461), .B(n15462), .Z(o[3042]) );
  AND U23192 ( .A(p_input[23042]), .B(p_input[13042]), .Z(n15462) );
  AND U23193 ( .A(p_input[33042]), .B(p_input[3042]), .Z(n15461) );
  AND U23194 ( .A(n15463), .B(n15464), .Z(o[3041]) );
  AND U23195 ( .A(p_input[23041]), .B(p_input[13041]), .Z(n15464) );
  AND U23196 ( .A(p_input[33041]), .B(p_input[3041]), .Z(n15463) );
  AND U23197 ( .A(n15465), .B(n15466), .Z(o[3040]) );
  AND U23198 ( .A(p_input[23040]), .B(p_input[13040]), .Z(n15466) );
  AND U23199 ( .A(p_input[33040]), .B(p_input[3040]), .Z(n15465) );
  AND U23200 ( .A(n15467), .B(n15468), .Z(o[303]) );
  AND U23201 ( .A(p_input[20303]), .B(p_input[10303]), .Z(n15468) );
  AND U23202 ( .A(p_input[303]), .B(p_input[30303]), .Z(n15467) );
  AND U23203 ( .A(n15469), .B(n15470), .Z(o[3039]) );
  AND U23204 ( .A(p_input[23039]), .B(p_input[13039]), .Z(n15470) );
  AND U23205 ( .A(p_input[33039]), .B(p_input[3039]), .Z(n15469) );
  AND U23206 ( .A(n15471), .B(n15472), .Z(o[3038]) );
  AND U23207 ( .A(p_input[23038]), .B(p_input[13038]), .Z(n15472) );
  AND U23208 ( .A(p_input[33038]), .B(p_input[3038]), .Z(n15471) );
  AND U23209 ( .A(n15473), .B(n15474), .Z(o[3037]) );
  AND U23210 ( .A(p_input[23037]), .B(p_input[13037]), .Z(n15474) );
  AND U23211 ( .A(p_input[33037]), .B(p_input[3037]), .Z(n15473) );
  AND U23212 ( .A(n15475), .B(n15476), .Z(o[3036]) );
  AND U23213 ( .A(p_input[23036]), .B(p_input[13036]), .Z(n15476) );
  AND U23214 ( .A(p_input[33036]), .B(p_input[3036]), .Z(n15475) );
  AND U23215 ( .A(n15477), .B(n15478), .Z(o[3035]) );
  AND U23216 ( .A(p_input[23035]), .B(p_input[13035]), .Z(n15478) );
  AND U23217 ( .A(p_input[33035]), .B(p_input[3035]), .Z(n15477) );
  AND U23218 ( .A(n15479), .B(n15480), .Z(o[3034]) );
  AND U23219 ( .A(p_input[23034]), .B(p_input[13034]), .Z(n15480) );
  AND U23220 ( .A(p_input[33034]), .B(p_input[3034]), .Z(n15479) );
  AND U23221 ( .A(n15481), .B(n15482), .Z(o[3033]) );
  AND U23222 ( .A(p_input[23033]), .B(p_input[13033]), .Z(n15482) );
  AND U23223 ( .A(p_input[33033]), .B(p_input[3033]), .Z(n15481) );
  AND U23224 ( .A(n15483), .B(n15484), .Z(o[3032]) );
  AND U23225 ( .A(p_input[23032]), .B(p_input[13032]), .Z(n15484) );
  AND U23226 ( .A(p_input[33032]), .B(p_input[3032]), .Z(n15483) );
  AND U23227 ( .A(n15485), .B(n15486), .Z(o[3031]) );
  AND U23228 ( .A(p_input[23031]), .B(p_input[13031]), .Z(n15486) );
  AND U23229 ( .A(p_input[33031]), .B(p_input[3031]), .Z(n15485) );
  AND U23230 ( .A(n15487), .B(n15488), .Z(o[3030]) );
  AND U23231 ( .A(p_input[23030]), .B(p_input[13030]), .Z(n15488) );
  AND U23232 ( .A(p_input[33030]), .B(p_input[3030]), .Z(n15487) );
  AND U23233 ( .A(n15489), .B(n15490), .Z(o[302]) );
  AND U23234 ( .A(p_input[20302]), .B(p_input[10302]), .Z(n15490) );
  AND U23235 ( .A(p_input[30302]), .B(p_input[302]), .Z(n15489) );
  AND U23236 ( .A(n15491), .B(n15492), .Z(o[3029]) );
  AND U23237 ( .A(p_input[23029]), .B(p_input[13029]), .Z(n15492) );
  AND U23238 ( .A(p_input[33029]), .B(p_input[3029]), .Z(n15491) );
  AND U23239 ( .A(n15493), .B(n15494), .Z(o[3028]) );
  AND U23240 ( .A(p_input[23028]), .B(p_input[13028]), .Z(n15494) );
  AND U23241 ( .A(p_input[33028]), .B(p_input[3028]), .Z(n15493) );
  AND U23242 ( .A(n15495), .B(n15496), .Z(o[3027]) );
  AND U23243 ( .A(p_input[23027]), .B(p_input[13027]), .Z(n15496) );
  AND U23244 ( .A(p_input[33027]), .B(p_input[3027]), .Z(n15495) );
  AND U23245 ( .A(n15497), .B(n15498), .Z(o[3026]) );
  AND U23246 ( .A(p_input[23026]), .B(p_input[13026]), .Z(n15498) );
  AND U23247 ( .A(p_input[33026]), .B(p_input[3026]), .Z(n15497) );
  AND U23248 ( .A(n15499), .B(n15500), .Z(o[3025]) );
  AND U23249 ( .A(p_input[23025]), .B(p_input[13025]), .Z(n15500) );
  AND U23250 ( .A(p_input[33025]), .B(p_input[3025]), .Z(n15499) );
  AND U23251 ( .A(n15501), .B(n15502), .Z(o[3024]) );
  AND U23252 ( .A(p_input[23024]), .B(p_input[13024]), .Z(n15502) );
  AND U23253 ( .A(p_input[33024]), .B(p_input[3024]), .Z(n15501) );
  AND U23254 ( .A(n15503), .B(n15504), .Z(o[3023]) );
  AND U23255 ( .A(p_input[23023]), .B(p_input[13023]), .Z(n15504) );
  AND U23256 ( .A(p_input[33023]), .B(p_input[3023]), .Z(n15503) );
  AND U23257 ( .A(n15505), .B(n15506), .Z(o[3022]) );
  AND U23258 ( .A(p_input[23022]), .B(p_input[13022]), .Z(n15506) );
  AND U23259 ( .A(p_input[33022]), .B(p_input[3022]), .Z(n15505) );
  AND U23260 ( .A(n15507), .B(n15508), .Z(o[3021]) );
  AND U23261 ( .A(p_input[23021]), .B(p_input[13021]), .Z(n15508) );
  AND U23262 ( .A(p_input[33021]), .B(p_input[3021]), .Z(n15507) );
  AND U23263 ( .A(n15509), .B(n15510), .Z(o[3020]) );
  AND U23264 ( .A(p_input[23020]), .B(p_input[13020]), .Z(n15510) );
  AND U23265 ( .A(p_input[33020]), .B(p_input[3020]), .Z(n15509) );
  AND U23266 ( .A(n15511), .B(n15512), .Z(o[301]) );
  AND U23267 ( .A(p_input[20301]), .B(p_input[10301]), .Z(n15512) );
  AND U23268 ( .A(p_input[30301]), .B(p_input[301]), .Z(n15511) );
  AND U23269 ( .A(n15513), .B(n15514), .Z(o[3019]) );
  AND U23270 ( .A(p_input[23019]), .B(p_input[13019]), .Z(n15514) );
  AND U23271 ( .A(p_input[33019]), .B(p_input[3019]), .Z(n15513) );
  AND U23272 ( .A(n15515), .B(n15516), .Z(o[3018]) );
  AND U23273 ( .A(p_input[23018]), .B(p_input[13018]), .Z(n15516) );
  AND U23274 ( .A(p_input[33018]), .B(p_input[3018]), .Z(n15515) );
  AND U23275 ( .A(n15517), .B(n15518), .Z(o[3017]) );
  AND U23276 ( .A(p_input[23017]), .B(p_input[13017]), .Z(n15518) );
  AND U23277 ( .A(p_input[33017]), .B(p_input[3017]), .Z(n15517) );
  AND U23278 ( .A(n15519), .B(n15520), .Z(o[3016]) );
  AND U23279 ( .A(p_input[23016]), .B(p_input[13016]), .Z(n15520) );
  AND U23280 ( .A(p_input[33016]), .B(p_input[3016]), .Z(n15519) );
  AND U23281 ( .A(n15521), .B(n15522), .Z(o[3015]) );
  AND U23282 ( .A(p_input[23015]), .B(p_input[13015]), .Z(n15522) );
  AND U23283 ( .A(p_input[33015]), .B(p_input[3015]), .Z(n15521) );
  AND U23284 ( .A(n15523), .B(n15524), .Z(o[3014]) );
  AND U23285 ( .A(p_input[23014]), .B(p_input[13014]), .Z(n15524) );
  AND U23286 ( .A(p_input[33014]), .B(p_input[3014]), .Z(n15523) );
  AND U23287 ( .A(n15525), .B(n15526), .Z(o[3013]) );
  AND U23288 ( .A(p_input[23013]), .B(p_input[13013]), .Z(n15526) );
  AND U23289 ( .A(p_input[33013]), .B(p_input[3013]), .Z(n15525) );
  AND U23290 ( .A(n15527), .B(n15528), .Z(o[3012]) );
  AND U23291 ( .A(p_input[23012]), .B(p_input[13012]), .Z(n15528) );
  AND U23292 ( .A(p_input[33012]), .B(p_input[3012]), .Z(n15527) );
  AND U23293 ( .A(n15529), .B(n15530), .Z(o[3011]) );
  AND U23294 ( .A(p_input[23011]), .B(p_input[13011]), .Z(n15530) );
  AND U23295 ( .A(p_input[33011]), .B(p_input[3011]), .Z(n15529) );
  AND U23296 ( .A(n15531), .B(n15532), .Z(o[3010]) );
  AND U23297 ( .A(p_input[23010]), .B(p_input[13010]), .Z(n15532) );
  AND U23298 ( .A(p_input[33010]), .B(p_input[3010]), .Z(n15531) );
  AND U23299 ( .A(n15533), .B(n15534), .Z(o[300]) );
  AND U23300 ( .A(p_input[20300]), .B(p_input[10300]), .Z(n15534) );
  AND U23301 ( .A(p_input[30300]), .B(p_input[300]), .Z(n15533) );
  AND U23302 ( .A(n15535), .B(n15536), .Z(o[3009]) );
  AND U23303 ( .A(p_input[23009]), .B(p_input[13009]), .Z(n15536) );
  AND U23304 ( .A(p_input[33009]), .B(p_input[3009]), .Z(n15535) );
  AND U23305 ( .A(n15537), .B(n15538), .Z(o[3008]) );
  AND U23306 ( .A(p_input[23008]), .B(p_input[13008]), .Z(n15538) );
  AND U23307 ( .A(p_input[33008]), .B(p_input[3008]), .Z(n15537) );
  AND U23308 ( .A(n15539), .B(n15540), .Z(o[3007]) );
  AND U23309 ( .A(p_input[23007]), .B(p_input[13007]), .Z(n15540) );
  AND U23310 ( .A(p_input[33007]), .B(p_input[3007]), .Z(n15539) );
  AND U23311 ( .A(n15541), .B(n15542), .Z(o[3006]) );
  AND U23312 ( .A(p_input[23006]), .B(p_input[13006]), .Z(n15542) );
  AND U23313 ( .A(p_input[33006]), .B(p_input[3006]), .Z(n15541) );
  AND U23314 ( .A(n15543), .B(n15544), .Z(o[3005]) );
  AND U23315 ( .A(p_input[23005]), .B(p_input[13005]), .Z(n15544) );
  AND U23316 ( .A(p_input[33005]), .B(p_input[3005]), .Z(n15543) );
  AND U23317 ( .A(n15545), .B(n15546), .Z(o[3004]) );
  AND U23318 ( .A(p_input[23004]), .B(p_input[13004]), .Z(n15546) );
  AND U23319 ( .A(p_input[33004]), .B(p_input[3004]), .Z(n15545) );
  AND U23320 ( .A(n15547), .B(n15548), .Z(o[3003]) );
  AND U23321 ( .A(p_input[23003]), .B(p_input[13003]), .Z(n15548) );
  AND U23322 ( .A(p_input[33003]), .B(p_input[3003]), .Z(n15547) );
  AND U23323 ( .A(n15549), .B(n15550), .Z(o[3002]) );
  AND U23324 ( .A(p_input[23002]), .B(p_input[13002]), .Z(n15550) );
  AND U23325 ( .A(p_input[33002]), .B(p_input[3002]), .Z(n15549) );
  AND U23326 ( .A(n15551), .B(n15552), .Z(o[3001]) );
  AND U23327 ( .A(p_input[23001]), .B(p_input[13001]), .Z(n15552) );
  AND U23328 ( .A(p_input[33001]), .B(p_input[3001]), .Z(n15551) );
  AND U23329 ( .A(n15553), .B(n15554), .Z(o[3000]) );
  AND U23330 ( .A(p_input[23000]), .B(p_input[13000]), .Z(n15554) );
  AND U23331 ( .A(p_input[33000]), .B(p_input[3000]), .Z(n15553) );
  AND U23332 ( .A(n15555), .B(n15556), .Z(o[2]) );
  AND U23333 ( .A(p_input[20002]), .B(p_input[10002]), .Z(n15556) );
  AND U23334 ( .A(p_input[30002]), .B(p_input[2]), .Z(n15555) );
  AND U23335 ( .A(n15557), .B(n15558), .Z(o[29]) );
  AND U23336 ( .A(p_input[20029]), .B(p_input[10029]), .Z(n15558) );
  AND U23337 ( .A(p_input[30029]), .B(p_input[29]), .Z(n15557) );
  AND U23338 ( .A(n15559), .B(n15560), .Z(o[299]) );
  AND U23339 ( .A(p_input[20299]), .B(p_input[10299]), .Z(n15560) );
  AND U23340 ( .A(p_input[30299]), .B(p_input[299]), .Z(n15559) );
  AND U23341 ( .A(n15561), .B(n15562), .Z(o[2999]) );
  AND U23342 ( .A(p_input[22999]), .B(p_input[12999]), .Z(n15562) );
  AND U23343 ( .A(p_input[32999]), .B(p_input[2999]), .Z(n15561) );
  AND U23344 ( .A(n15563), .B(n15564), .Z(o[2998]) );
  AND U23345 ( .A(p_input[22998]), .B(p_input[12998]), .Z(n15564) );
  AND U23346 ( .A(p_input[32998]), .B(p_input[2998]), .Z(n15563) );
  AND U23347 ( .A(n15565), .B(n15566), .Z(o[2997]) );
  AND U23348 ( .A(p_input[22997]), .B(p_input[12997]), .Z(n15566) );
  AND U23349 ( .A(p_input[32997]), .B(p_input[2997]), .Z(n15565) );
  AND U23350 ( .A(n15567), .B(n15568), .Z(o[2996]) );
  AND U23351 ( .A(p_input[22996]), .B(p_input[12996]), .Z(n15568) );
  AND U23352 ( .A(p_input[32996]), .B(p_input[2996]), .Z(n15567) );
  AND U23353 ( .A(n15569), .B(n15570), .Z(o[2995]) );
  AND U23354 ( .A(p_input[22995]), .B(p_input[12995]), .Z(n15570) );
  AND U23355 ( .A(p_input[32995]), .B(p_input[2995]), .Z(n15569) );
  AND U23356 ( .A(n15571), .B(n15572), .Z(o[2994]) );
  AND U23357 ( .A(p_input[22994]), .B(p_input[12994]), .Z(n15572) );
  AND U23358 ( .A(p_input[32994]), .B(p_input[2994]), .Z(n15571) );
  AND U23359 ( .A(n15573), .B(n15574), .Z(o[2993]) );
  AND U23360 ( .A(p_input[22993]), .B(p_input[12993]), .Z(n15574) );
  AND U23361 ( .A(p_input[32993]), .B(p_input[2993]), .Z(n15573) );
  AND U23362 ( .A(n15575), .B(n15576), .Z(o[2992]) );
  AND U23363 ( .A(p_input[22992]), .B(p_input[12992]), .Z(n15576) );
  AND U23364 ( .A(p_input[32992]), .B(p_input[2992]), .Z(n15575) );
  AND U23365 ( .A(n15577), .B(n15578), .Z(o[2991]) );
  AND U23366 ( .A(p_input[22991]), .B(p_input[12991]), .Z(n15578) );
  AND U23367 ( .A(p_input[32991]), .B(p_input[2991]), .Z(n15577) );
  AND U23368 ( .A(n15579), .B(n15580), .Z(o[2990]) );
  AND U23369 ( .A(p_input[22990]), .B(p_input[12990]), .Z(n15580) );
  AND U23370 ( .A(p_input[32990]), .B(p_input[2990]), .Z(n15579) );
  AND U23371 ( .A(n15581), .B(n15582), .Z(o[298]) );
  AND U23372 ( .A(p_input[20298]), .B(p_input[10298]), .Z(n15582) );
  AND U23373 ( .A(p_input[30298]), .B(p_input[298]), .Z(n15581) );
  AND U23374 ( .A(n15583), .B(n15584), .Z(o[2989]) );
  AND U23375 ( .A(p_input[22989]), .B(p_input[12989]), .Z(n15584) );
  AND U23376 ( .A(p_input[32989]), .B(p_input[2989]), .Z(n15583) );
  AND U23377 ( .A(n15585), .B(n15586), .Z(o[2988]) );
  AND U23378 ( .A(p_input[22988]), .B(p_input[12988]), .Z(n15586) );
  AND U23379 ( .A(p_input[32988]), .B(p_input[2988]), .Z(n15585) );
  AND U23380 ( .A(n15587), .B(n15588), .Z(o[2987]) );
  AND U23381 ( .A(p_input[22987]), .B(p_input[12987]), .Z(n15588) );
  AND U23382 ( .A(p_input[32987]), .B(p_input[2987]), .Z(n15587) );
  AND U23383 ( .A(n15589), .B(n15590), .Z(o[2986]) );
  AND U23384 ( .A(p_input[22986]), .B(p_input[12986]), .Z(n15590) );
  AND U23385 ( .A(p_input[32986]), .B(p_input[2986]), .Z(n15589) );
  AND U23386 ( .A(n15591), .B(n15592), .Z(o[2985]) );
  AND U23387 ( .A(p_input[22985]), .B(p_input[12985]), .Z(n15592) );
  AND U23388 ( .A(p_input[32985]), .B(p_input[2985]), .Z(n15591) );
  AND U23389 ( .A(n15593), .B(n15594), .Z(o[2984]) );
  AND U23390 ( .A(p_input[22984]), .B(p_input[12984]), .Z(n15594) );
  AND U23391 ( .A(p_input[32984]), .B(p_input[2984]), .Z(n15593) );
  AND U23392 ( .A(n15595), .B(n15596), .Z(o[2983]) );
  AND U23393 ( .A(p_input[22983]), .B(p_input[12983]), .Z(n15596) );
  AND U23394 ( .A(p_input[32983]), .B(p_input[2983]), .Z(n15595) );
  AND U23395 ( .A(n15597), .B(n15598), .Z(o[2982]) );
  AND U23396 ( .A(p_input[22982]), .B(p_input[12982]), .Z(n15598) );
  AND U23397 ( .A(p_input[32982]), .B(p_input[2982]), .Z(n15597) );
  AND U23398 ( .A(n15599), .B(n15600), .Z(o[2981]) );
  AND U23399 ( .A(p_input[22981]), .B(p_input[12981]), .Z(n15600) );
  AND U23400 ( .A(p_input[32981]), .B(p_input[2981]), .Z(n15599) );
  AND U23401 ( .A(n15601), .B(n15602), .Z(o[2980]) );
  AND U23402 ( .A(p_input[22980]), .B(p_input[12980]), .Z(n15602) );
  AND U23403 ( .A(p_input[32980]), .B(p_input[2980]), .Z(n15601) );
  AND U23404 ( .A(n15603), .B(n15604), .Z(o[297]) );
  AND U23405 ( .A(p_input[20297]), .B(p_input[10297]), .Z(n15604) );
  AND U23406 ( .A(p_input[30297]), .B(p_input[297]), .Z(n15603) );
  AND U23407 ( .A(n15605), .B(n15606), .Z(o[2979]) );
  AND U23408 ( .A(p_input[22979]), .B(p_input[12979]), .Z(n15606) );
  AND U23409 ( .A(p_input[32979]), .B(p_input[2979]), .Z(n15605) );
  AND U23410 ( .A(n15607), .B(n15608), .Z(o[2978]) );
  AND U23411 ( .A(p_input[22978]), .B(p_input[12978]), .Z(n15608) );
  AND U23412 ( .A(p_input[32978]), .B(p_input[2978]), .Z(n15607) );
  AND U23413 ( .A(n15609), .B(n15610), .Z(o[2977]) );
  AND U23414 ( .A(p_input[22977]), .B(p_input[12977]), .Z(n15610) );
  AND U23415 ( .A(p_input[32977]), .B(p_input[2977]), .Z(n15609) );
  AND U23416 ( .A(n15611), .B(n15612), .Z(o[2976]) );
  AND U23417 ( .A(p_input[22976]), .B(p_input[12976]), .Z(n15612) );
  AND U23418 ( .A(p_input[32976]), .B(p_input[2976]), .Z(n15611) );
  AND U23419 ( .A(n15613), .B(n15614), .Z(o[2975]) );
  AND U23420 ( .A(p_input[22975]), .B(p_input[12975]), .Z(n15614) );
  AND U23421 ( .A(p_input[32975]), .B(p_input[2975]), .Z(n15613) );
  AND U23422 ( .A(n15615), .B(n15616), .Z(o[2974]) );
  AND U23423 ( .A(p_input[22974]), .B(p_input[12974]), .Z(n15616) );
  AND U23424 ( .A(p_input[32974]), .B(p_input[2974]), .Z(n15615) );
  AND U23425 ( .A(n15617), .B(n15618), .Z(o[2973]) );
  AND U23426 ( .A(p_input[22973]), .B(p_input[12973]), .Z(n15618) );
  AND U23427 ( .A(p_input[32973]), .B(p_input[2973]), .Z(n15617) );
  AND U23428 ( .A(n15619), .B(n15620), .Z(o[2972]) );
  AND U23429 ( .A(p_input[22972]), .B(p_input[12972]), .Z(n15620) );
  AND U23430 ( .A(p_input[32972]), .B(p_input[2972]), .Z(n15619) );
  AND U23431 ( .A(n15621), .B(n15622), .Z(o[2971]) );
  AND U23432 ( .A(p_input[22971]), .B(p_input[12971]), .Z(n15622) );
  AND U23433 ( .A(p_input[32971]), .B(p_input[2971]), .Z(n15621) );
  AND U23434 ( .A(n15623), .B(n15624), .Z(o[2970]) );
  AND U23435 ( .A(p_input[22970]), .B(p_input[12970]), .Z(n15624) );
  AND U23436 ( .A(p_input[32970]), .B(p_input[2970]), .Z(n15623) );
  AND U23437 ( .A(n15625), .B(n15626), .Z(o[296]) );
  AND U23438 ( .A(p_input[20296]), .B(p_input[10296]), .Z(n15626) );
  AND U23439 ( .A(p_input[30296]), .B(p_input[296]), .Z(n15625) );
  AND U23440 ( .A(n15627), .B(n15628), .Z(o[2969]) );
  AND U23441 ( .A(p_input[22969]), .B(p_input[12969]), .Z(n15628) );
  AND U23442 ( .A(p_input[32969]), .B(p_input[2969]), .Z(n15627) );
  AND U23443 ( .A(n15629), .B(n15630), .Z(o[2968]) );
  AND U23444 ( .A(p_input[22968]), .B(p_input[12968]), .Z(n15630) );
  AND U23445 ( .A(p_input[32968]), .B(p_input[2968]), .Z(n15629) );
  AND U23446 ( .A(n15631), .B(n15632), .Z(o[2967]) );
  AND U23447 ( .A(p_input[22967]), .B(p_input[12967]), .Z(n15632) );
  AND U23448 ( .A(p_input[32967]), .B(p_input[2967]), .Z(n15631) );
  AND U23449 ( .A(n15633), .B(n15634), .Z(o[2966]) );
  AND U23450 ( .A(p_input[22966]), .B(p_input[12966]), .Z(n15634) );
  AND U23451 ( .A(p_input[32966]), .B(p_input[2966]), .Z(n15633) );
  AND U23452 ( .A(n15635), .B(n15636), .Z(o[2965]) );
  AND U23453 ( .A(p_input[22965]), .B(p_input[12965]), .Z(n15636) );
  AND U23454 ( .A(p_input[32965]), .B(p_input[2965]), .Z(n15635) );
  AND U23455 ( .A(n15637), .B(n15638), .Z(o[2964]) );
  AND U23456 ( .A(p_input[22964]), .B(p_input[12964]), .Z(n15638) );
  AND U23457 ( .A(p_input[32964]), .B(p_input[2964]), .Z(n15637) );
  AND U23458 ( .A(n15639), .B(n15640), .Z(o[2963]) );
  AND U23459 ( .A(p_input[22963]), .B(p_input[12963]), .Z(n15640) );
  AND U23460 ( .A(p_input[32963]), .B(p_input[2963]), .Z(n15639) );
  AND U23461 ( .A(n15641), .B(n15642), .Z(o[2962]) );
  AND U23462 ( .A(p_input[22962]), .B(p_input[12962]), .Z(n15642) );
  AND U23463 ( .A(p_input[32962]), .B(p_input[2962]), .Z(n15641) );
  AND U23464 ( .A(n15643), .B(n15644), .Z(o[2961]) );
  AND U23465 ( .A(p_input[22961]), .B(p_input[12961]), .Z(n15644) );
  AND U23466 ( .A(p_input[32961]), .B(p_input[2961]), .Z(n15643) );
  AND U23467 ( .A(n15645), .B(n15646), .Z(o[2960]) );
  AND U23468 ( .A(p_input[22960]), .B(p_input[12960]), .Z(n15646) );
  AND U23469 ( .A(p_input[32960]), .B(p_input[2960]), .Z(n15645) );
  AND U23470 ( .A(n15647), .B(n15648), .Z(o[295]) );
  AND U23471 ( .A(p_input[20295]), .B(p_input[10295]), .Z(n15648) );
  AND U23472 ( .A(p_input[30295]), .B(p_input[295]), .Z(n15647) );
  AND U23473 ( .A(n15649), .B(n15650), .Z(o[2959]) );
  AND U23474 ( .A(p_input[22959]), .B(p_input[12959]), .Z(n15650) );
  AND U23475 ( .A(p_input[32959]), .B(p_input[2959]), .Z(n15649) );
  AND U23476 ( .A(n15651), .B(n15652), .Z(o[2958]) );
  AND U23477 ( .A(p_input[22958]), .B(p_input[12958]), .Z(n15652) );
  AND U23478 ( .A(p_input[32958]), .B(p_input[2958]), .Z(n15651) );
  AND U23479 ( .A(n15653), .B(n15654), .Z(o[2957]) );
  AND U23480 ( .A(p_input[22957]), .B(p_input[12957]), .Z(n15654) );
  AND U23481 ( .A(p_input[32957]), .B(p_input[2957]), .Z(n15653) );
  AND U23482 ( .A(n15655), .B(n15656), .Z(o[2956]) );
  AND U23483 ( .A(p_input[22956]), .B(p_input[12956]), .Z(n15656) );
  AND U23484 ( .A(p_input[32956]), .B(p_input[2956]), .Z(n15655) );
  AND U23485 ( .A(n15657), .B(n15658), .Z(o[2955]) );
  AND U23486 ( .A(p_input[22955]), .B(p_input[12955]), .Z(n15658) );
  AND U23487 ( .A(p_input[32955]), .B(p_input[2955]), .Z(n15657) );
  AND U23488 ( .A(n15659), .B(n15660), .Z(o[2954]) );
  AND U23489 ( .A(p_input[22954]), .B(p_input[12954]), .Z(n15660) );
  AND U23490 ( .A(p_input[32954]), .B(p_input[2954]), .Z(n15659) );
  AND U23491 ( .A(n15661), .B(n15662), .Z(o[2953]) );
  AND U23492 ( .A(p_input[22953]), .B(p_input[12953]), .Z(n15662) );
  AND U23493 ( .A(p_input[32953]), .B(p_input[2953]), .Z(n15661) );
  AND U23494 ( .A(n15663), .B(n15664), .Z(o[2952]) );
  AND U23495 ( .A(p_input[22952]), .B(p_input[12952]), .Z(n15664) );
  AND U23496 ( .A(p_input[32952]), .B(p_input[2952]), .Z(n15663) );
  AND U23497 ( .A(n15665), .B(n15666), .Z(o[2951]) );
  AND U23498 ( .A(p_input[22951]), .B(p_input[12951]), .Z(n15666) );
  AND U23499 ( .A(p_input[32951]), .B(p_input[2951]), .Z(n15665) );
  AND U23500 ( .A(n15667), .B(n15668), .Z(o[2950]) );
  AND U23501 ( .A(p_input[22950]), .B(p_input[12950]), .Z(n15668) );
  AND U23502 ( .A(p_input[32950]), .B(p_input[2950]), .Z(n15667) );
  AND U23503 ( .A(n15669), .B(n15670), .Z(o[294]) );
  AND U23504 ( .A(p_input[20294]), .B(p_input[10294]), .Z(n15670) );
  AND U23505 ( .A(p_input[30294]), .B(p_input[294]), .Z(n15669) );
  AND U23506 ( .A(n15671), .B(n15672), .Z(o[2949]) );
  AND U23507 ( .A(p_input[22949]), .B(p_input[12949]), .Z(n15672) );
  AND U23508 ( .A(p_input[32949]), .B(p_input[2949]), .Z(n15671) );
  AND U23509 ( .A(n15673), .B(n15674), .Z(o[2948]) );
  AND U23510 ( .A(p_input[22948]), .B(p_input[12948]), .Z(n15674) );
  AND U23511 ( .A(p_input[32948]), .B(p_input[2948]), .Z(n15673) );
  AND U23512 ( .A(n15675), .B(n15676), .Z(o[2947]) );
  AND U23513 ( .A(p_input[22947]), .B(p_input[12947]), .Z(n15676) );
  AND U23514 ( .A(p_input[32947]), .B(p_input[2947]), .Z(n15675) );
  AND U23515 ( .A(n15677), .B(n15678), .Z(o[2946]) );
  AND U23516 ( .A(p_input[22946]), .B(p_input[12946]), .Z(n15678) );
  AND U23517 ( .A(p_input[32946]), .B(p_input[2946]), .Z(n15677) );
  AND U23518 ( .A(n15679), .B(n15680), .Z(o[2945]) );
  AND U23519 ( .A(p_input[22945]), .B(p_input[12945]), .Z(n15680) );
  AND U23520 ( .A(p_input[32945]), .B(p_input[2945]), .Z(n15679) );
  AND U23521 ( .A(n15681), .B(n15682), .Z(o[2944]) );
  AND U23522 ( .A(p_input[22944]), .B(p_input[12944]), .Z(n15682) );
  AND U23523 ( .A(p_input[32944]), .B(p_input[2944]), .Z(n15681) );
  AND U23524 ( .A(n15683), .B(n15684), .Z(o[2943]) );
  AND U23525 ( .A(p_input[22943]), .B(p_input[12943]), .Z(n15684) );
  AND U23526 ( .A(p_input[32943]), .B(p_input[2943]), .Z(n15683) );
  AND U23527 ( .A(n15685), .B(n15686), .Z(o[2942]) );
  AND U23528 ( .A(p_input[22942]), .B(p_input[12942]), .Z(n15686) );
  AND U23529 ( .A(p_input[32942]), .B(p_input[2942]), .Z(n15685) );
  AND U23530 ( .A(n15687), .B(n15688), .Z(o[2941]) );
  AND U23531 ( .A(p_input[22941]), .B(p_input[12941]), .Z(n15688) );
  AND U23532 ( .A(p_input[32941]), .B(p_input[2941]), .Z(n15687) );
  AND U23533 ( .A(n15689), .B(n15690), .Z(o[2940]) );
  AND U23534 ( .A(p_input[22940]), .B(p_input[12940]), .Z(n15690) );
  AND U23535 ( .A(p_input[32940]), .B(p_input[2940]), .Z(n15689) );
  AND U23536 ( .A(n15691), .B(n15692), .Z(o[293]) );
  AND U23537 ( .A(p_input[20293]), .B(p_input[10293]), .Z(n15692) );
  AND U23538 ( .A(p_input[30293]), .B(p_input[293]), .Z(n15691) );
  AND U23539 ( .A(n15693), .B(n15694), .Z(o[2939]) );
  AND U23540 ( .A(p_input[22939]), .B(p_input[12939]), .Z(n15694) );
  AND U23541 ( .A(p_input[32939]), .B(p_input[2939]), .Z(n15693) );
  AND U23542 ( .A(n15695), .B(n15696), .Z(o[2938]) );
  AND U23543 ( .A(p_input[22938]), .B(p_input[12938]), .Z(n15696) );
  AND U23544 ( .A(p_input[32938]), .B(p_input[2938]), .Z(n15695) );
  AND U23545 ( .A(n15697), .B(n15698), .Z(o[2937]) );
  AND U23546 ( .A(p_input[22937]), .B(p_input[12937]), .Z(n15698) );
  AND U23547 ( .A(p_input[32937]), .B(p_input[2937]), .Z(n15697) );
  AND U23548 ( .A(n15699), .B(n15700), .Z(o[2936]) );
  AND U23549 ( .A(p_input[22936]), .B(p_input[12936]), .Z(n15700) );
  AND U23550 ( .A(p_input[32936]), .B(p_input[2936]), .Z(n15699) );
  AND U23551 ( .A(n15701), .B(n15702), .Z(o[2935]) );
  AND U23552 ( .A(p_input[22935]), .B(p_input[12935]), .Z(n15702) );
  AND U23553 ( .A(p_input[32935]), .B(p_input[2935]), .Z(n15701) );
  AND U23554 ( .A(n15703), .B(n15704), .Z(o[2934]) );
  AND U23555 ( .A(p_input[22934]), .B(p_input[12934]), .Z(n15704) );
  AND U23556 ( .A(p_input[32934]), .B(p_input[2934]), .Z(n15703) );
  AND U23557 ( .A(n15705), .B(n15706), .Z(o[2933]) );
  AND U23558 ( .A(p_input[22933]), .B(p_input[12933]), .Z(n15706) );
  AND U23559 ( .A(p_input[32933]), .B(p_input[2933]), .Z(n15705) );
  AND U23560 ( .A(n15707), .B(n15708), .Z(o[2932]) );
  AND U23561 ( .A(p_input[22932]), .B(p_input[12932]), .Z(n15708) );
  AND U23562 ( .A(p_input[32932]), .B(p_input[2932]), .Z(n15707) );
  AND U23563 ( .A(n15709), .B(n15710), .Z(o[2931]) );
  AND U23564 ( .A(p_input[22931]), .B(p_input[12931]), .Z(n15710) );
  AND U23565 ( .A(p_input[32931]), .B(p_input[2931]), .Z(n15709) );
  AND U23566 ( .A(n15711), .B(n15712), .Z(o[2930]) );
  AND U23567 ( .A(p_input[22930]), .B(p_input[12930]), .Z(n15712) );
  AND U23568 ( .A(p_input[32930]), .B(p_input[2930]), .Z(n15711) );
  AND U23569 ( .A(n15713), .B(n15714), .Z(o[292]) );
  AND U23570 ( .A(p_input[20292]), .B(p_input[10292]), .Z(n15714) );
  AND U23571 ( .A(p_input[30292]), .B(p_input[292]), .Z(n15713) );
  AND U23572 ( .A(n15715), .B(n15716), .Z(o[2929]) );
  AND U23573 ( .A(p_input[22929]), .B(p_input[12929]), .Z(n15716) );
  AND U23574 ( .A(p_input[32929]), .B(p_input[2929]), .Z(n15715) );
  AND U23575 ( .A(n15717), .B(n15718), .Z(o[2928]) );
  AND U23576 ( .A(p_input[22928]), .B(p_input[12928]), .Z(n15718) );
  AND U23577 ( .A(p_input[32928]), .B(p_input[2928]), .Z(n15717) );
  AND U23578 ( .A(n15719), .B(n15720), .Z(o[2927]) );
  AND U23579 ( .A(p_input[22927]), .B(p_input[12927]), .Z(n15720) );
  AND U23580 ( .A(p_input[32927]), .B(p_input[2927]), .Z(n15719) );
  AND U23581 ( .A(n15721), .B(n15722), .Z(o[2926]) );
  AND U23582 ( .A(p_input[22926]), .B(p_input[12926]), .Z(n15722) );
  AND U23583 ( .A(p_input[32926]), .B(p_input[2926]), .Z(n15721) );
  AND U23584 ( .A(n15723), .B(n15724), .Z(o[2925]) );
  AND U23585 ( .A(p_input[22925]), .B(p_input[12925]), .Z(n15724) );
  AND U23586 ( .A(p_input[32925]), .B(p_input[2925]), .Z(n15723) );
  AND U23587 ( .A(n15725), .B(n15726), .Z(o[2924]) );
  AND U23588 ( .A(p_input[22924]), .B(p_input[12924]), .Z(n15726) );
  AND U23589 ( .A(p_input[32924]), .B(p_input[2924]), .Z(n15725) );
  AND U23590 ( .A(n15727), .B(n15728), .Z(o[2923]) );
  AND U23591 ( .A(p_input[22923]), .B(p_input[12923]), .Z(n15728) );
  AND U23592 ( .A(p_input[32923]), .B(p_input[2923]), .Z(n15727) );
  AND U23593 ( .A(n15729), .B(n15730), .Z(o[2922]) );
  AND U23594 ( .A(p_input[22922]), .B(p_input[12922]), .Z(n15730) );
  AND U23595 ( .A(p_input[32922]), .B(p_input[2922]), .Z(n15729) );
  AND U23596 ( .A(n15731), .B(n15732), .Z(o[2921]) );
  AND U23597 ( .A(p_input[22921]), .B(p_input[12921]), .Z(n15732) );
  AND U23598 ( .A(p_input[32921]), .B(p_input[2921]), .Z(n15731) );
  AND U23599 ( .A(n15733), .B(n15734), .Z(o[2920]) );
  AND U23600 ( .A(p_input[22920]), .B(p_input[12920]), .Z(n15734) );
  AND U23601 ( .A(p_input[32920]), .B(p_input[2920]), .Z(n15733) );
  AND U23602 ( .A(n15735), .B(n15736), .Z(o[291]) );
  AND U23603 ( .A(p_input[20291]), .B(p_input[10291]), .Z(n15736) );
  AND U23604 ( .A(p_input[30291]), .B(p_input[291]), .Z(n15735) );
  AND U23605 ( .A(n15737), .B(n15738), .Z(o[2919]) );
  AND U23606 ( .A(p_input[22919]), .B(p_input[12919]), .Z(n15738) );
  AND U23607 ( .A(p_input[32919]), .B(p_input[2919]), .Z(n15737) );
  AND U23608 ( .A(n15739), .B(n15740), .Z(o[2918]) );
  AND U23609 ( .A(p_input[22918]), .B(p_input[12918]), .Z(n15740) );
  AND U23610 ( .A(p_input[32918]), .B(p_input[2918]), .Z(n15739) );
  AND U23611 ( .A(n15741), .B(n15742), .Z(o[2917]) );
  AND U23612 ( .A(p_input[22917]), .B(p_input[12917]), .Z(n15742) );
  AND U23613 ( .A(p_input[32917]), .B(p_input[2917]), .Z(n15741) );
  AND U23614 ( .A(n15743), .B(n15744), .Z(o[2916]) );
  AND U23615 ( .A(p_input[22916]), .B(p_input[12916]), .Z(n15744) );
  AND U23616 ( .A(p_input[32916]), .B(p_input[2916]), .Z(n15743) );
  AND U23617 ( .A(n15745), .B(n15746), .Z(o[2915]) );
  AND U23618 ( .A(p_input[22915]), .B(p_input[12915]), .Z(n15746) );
  AND U23619 ( .A(p_input[32915]), .B(p_input[2915]), .Z(n15745) );
  AND U23620 ( .A(n15747), .B(n15748), .Z(o[2914]) );
  AND U23621 ( .A(p_input[22914]), .B(p_input[12914]), .Z(n15748) );
  AND U23622 ( .A(p_input[32914]), .B(p_input[2914]), .Z(n15747) );
  AND U23623 ( .A(n15749), .B(n15750), .Z(o[2913]) );
  AND U23624 ( .A(p_input[22913]), .B(p_input[12913]), .Z(n15750) );
  AND U23625 ( .A(p_input[32913]), .B(p_input[2913]), .Z(n15749) );
  AND U23626 ( .A(n15751), .B(n15752), .Z(o[2912]) );
  AND U23627 ( .A(p_input[22912]), .B(p_input[12912]), .Z(n15752) );
  AND U23628 ( .A(p_input[32912]), .B(p_input[2912]), .Z(n15751) );
  AND U23629 ( .A(n15753), .B(n15754), .Z(o[2911]) );
  AND U23630 ( .A(p_input[22911]), .B(p_input[12911]), .Z(n15754) );
  AND U23631 ( .A(p_input[32911]), .B(p_input[2911]), .Z(n15753) );
  AND U23632 ( .A(n15755), .B(n15756), .Z(o[2910]) );
  AND U23633 ( .A(p_input[22910]), .B(p_input[12910]), .Z(n15756) );
  AND U23634 ( .A(p_input[32910]), .B(p_input[2910]), .Z(n15755) );
  AND U23635 ( .A(n15757), .B(n15758), .Z(o[290]) );
  AND U23636 ( .A(p_input[20290]), .B(p_input[10290]), .Z(n15758) );
  AND U23637 ( .A(p_input[30290]), .B(p_input[290]), .Z(n15757) );
  AND U23638 ( .A(n15759), .B(n15760), .Z(o[2909]) );
  AND U23639 ( .A(p_input[22909]), .B(p_input[12909]), .Z(n15760) );
  AND U23640 ( .A(p_input[32909]), .B(p_input[2909]), .Z(n15759) );
  AND U23641 ( .A(n15761), .B(n15762), .Z(o[2908]) );
  AND U23642 ( .A(p_input[22908]), .B(p_input[12908]), .Z(n15762) );
  AND U23643 ( .A(p_input[32908]), .B(p_input[2908]), .Z(n15761) );
  AND U23644 ( .A(n15763), .B(n15764), .Z(o[2907]) );
  AND U23645 ( .A(p_input[22907]), .B(p_input[12907]), .Z(n15764) );
  AND U23646 ( .A(p_input[32907]), .B(p_input[2907]), .Z(n15763) );
  AND U23647 ( .A(n15765), .B(n15766), .Z(o[2906]) );
  AND U23648 ( .A(p_input[22906]), .B(p_input[12906]), .Z(n15766) );
  AND U23649 ( .A(p_input[32906]), .B(p_input[2906]), .Z(n15765) );
  AND U23650 ( .A(n15767), .B(n15768), .Z(o[2905]) );
  AND U23651 ( .A(p_input[22905]), .B(p_input[12905]), .Z(n15768) );
  AND U23652 ( .A(p_input[32905]), .B(p_input[2905]), .Z(n15767) );
  AND U23653 ( .A(n15769), .B(n15770), .Z(o[2904]) );
  AND U23654 ( .A(p_input[22904]), .B(p_input[12904]), .Z(n15770) );
  AND U23655 ( .A(p_input[32904]), .B(p_input[2904]), .Z(n15769) );
  AND U23656 ( .A(n15771), .B(n15772), .Z(o[2903]) );
  AND U23657 ( .A(p_input[22903]), .B(p_input[12903]), .Z(n15772) );
  AND U23658 ( .A(p_input[32903]), .B(p_input[2903]), .Z(n15771) );
  AND U23659 ( .A(n15773), .B(n15774), .Z(o[2902]) );
  AND U23660 ( .A(p_input[22902]), .B(p_input[12902]), .Z(n15774) );
  AND U23661 ( .A(p_input[32902]), .B(p_input[2902]), .Z(n15773) );
  AND U23662 ( .A(n15775), .B(n15776), .Z(o[2901]) );
  AND U23663 ( .A(p_input[22901]), .B(p_input[12901]), .Z(n15776) );
  AND U23664 ( .A(p_input[32901]), .B(p_input[2901]), .Z(n15775) );
  AND U23665 ( .A(n15777), .B(n15778), .Z(o[2900]) );
  AND U23666 ( .A(p_input[22900]), .B(p_input[12900]), .Z(n15778) );
  AND U23667 ( .A(p_input[32900]), .B(p_input[2900]), .Z(n15777) );
  AND U23668 ( .A(n15779), .B(n15780), .Z(o[28]) );
  AND U23669 ( .A(p_input[20028]), .B(p_input[10028]), .Z(n15780) );
  AND U23670 ( .A(p_input[30028]), .B(p_input[28]), .Z(n15779) );
  AND U23671 ( .A(n15781), .B(n15782), .Z(o[289]) );
  AND U23672 ( .A(p_input[20289]), .B(p_input[10289]), .Z(n15782) );
  AND U23673 ( .A(p_input[30289]), .B(p_input[289]), .Z(n15781) );
  AND U23674 ( .A(n15783), .B(n15784), .Z(o[2899]) );
  AND U23675 ( .A(p_input[22899]), .B(p_input[12899]), .Z(n15784) );
  AND U23676 ( .A(p_input[32899]), .B(p_input[2899]), .Z(n15783) );
  AND U23677 ( .A(n15785), .B(n15786), .Z(o[2898]) );
  AND U23678 ( .A(p_input[22898]), .B(p_input[12898]), .Z(n15786) );
  AND U23679 ( .A(p_input[32898]), .B(p_input[2898]), .Z(n15785) );
  AND U23680 ( .A(n15787), .B(n15788), .Z(o[2897]) );
  AND U23681 ( .A(p_input[22897]), .B(p_input[12897]), .Z(n15788) );
  AND U23682 ( .A(p_input[32897]), .B(p_input[2897]), .Z(n15787) );
  AND U23683 ( .A(n15789), .B(n15790), .Z(o[2896]) );
  AND U23684 ( .A(p_input[22896]), .B(p_input[12896]), .Z(n15790) );
  AND U23685 ( .A(p_input[32896]), .B(p_input[2896]), .Z(n15789) );
  AND U23686 ( .A(n15791), .B(n15792), .Z(o[2895]) );
  AND U23687 ( .A(p_input[22895]), .B(p_input[12895]), .Z(n15792) );
  AND U23688 ( .A(p_input[32895]), .B(p_input[2895]), .Z(n15791) );
  AND U23689 ( .A(n15793), .B(n15794), .Z(o[2894]) );
  AND U23690 ( .A(p_input[22894]), .B(p_input[12894]), .Z(n15794) );
  AND U23691 ( .A(p_input[32894]), .B(p_input[2894]), .Z(n15793) );
  AND U23692 ( .A(n15795), .B(n15796), .Z(o[2893]) );
  AND U23693 ( .A(p_input[22893]), .B(p_input[12893]), .Z(n15796) );
  AND U23694 ( .A(p_input[32893]), .B(p_input[2893]), .Z(n15795) );
  AND U23695 ( .A(n15797), .B(n15798), .Z(o[2892]) );
  AND U23696 ( .A(p_input[22892]), .B(p_input[12892]), .Z(n15798) );
  AND U23697 ( .A(p_input[32892]), .B(p_input[2892]), .Z(n15797) );
  AND U23698 ( .A(n15799), .B(n15800), .Z(o[2891]) );
  AND U23699 ( .A(p_input[22891]), .B(p_input[12891]), .Z(n15800) );
  AND U23700 ( .A(p_input[32891]), .B(p_input[2891]), .Z(n15799) );
  AND U23701 ( .A(n15801), .B(n15802), .Z(o[2890]) );
  AND U23702 ( .A(p_input[22890]), .B(p_input[12890]), .Z(n15802) );
  AND U23703 ( .A(p_input[32890]), .B(p_input[2890]), .Z(n15801) );
  AND U23704 ( .A(n15803), .B(n15804), .Z(o[288]) );
  AND U23705 ( .A(p_input[20288]), .B(p_input[10288]), .Z(n15804) );
  AND U23706 ( .A(p_input[30288]), .B(p_input[288]), .Z(n15803) );
  AND U23707 ( .A(n15805), .B(n15806), .Z(o[2889]) );
  AND U23708 ( .A(p_input[22889]), .B(p_input[12889]), .Z(n15806) );
  AND U23709 ( .A(p_input[32889]), .B(p_input[2889]), .Z(n15805) );
  AND U23710 ( .A(n15807), .B(n15808), .Z(o[2888]) );
  AND U23711 ( .A(p_input[22888]), .B(p_input[12888]), .Z(n15808) );
  AND U23712 ( .A(p_input[32888]), .B(p_input[2888]), .Z(n15807) );
  AND U23713 ( .A(n15809), .B(n15810), .Z(o[2887]) );
  AND U23714 ( .A(p_input[22887]), .B(p_input[12887]), .Z(n15810) );
  AND U23715 ( .A(p_input[32887]), .B(p_input[2887]), .Z(n15809) );
  AND U23716 ( .A(n15811), .B(n15812), .Z(o[2886]) );
  AND U23717 ( .A(p_input[22886]), .B(p_input[12886]), .Z(n15812) );
  AND U23718 ( .A(p_input[32886]), .B(p_input[2886]), .Z(n15811) );
  AND U23719 ( .A(n15813), .B(n15814), .Z(o[2885]) );
  AND U23720 ( .A(p_input[22885]), .B(p_input[12885]), .Z(n15814) );
  AND U23721 ( .A(p_input[32885]), .B(p_input[2885]), .Z(n15813) );
  AND U23722 ( .A(n15815), .B(n15816), .Z(o[2884]) );
  AND U23723 ( .A(p_input[22884]), .B(p_input[12884]), .Z(n15816) );
  AND U23724 ( .A(p_input[32884]), .B(p_input[2884]), .Z(n15815) );
  AND U23725 ( .A(n15817), .B(n15818), .Z(o[2883]) );
  AND U23726 ( .A(p_input[22883]), .B(p_input[12883]), .Z(n15818) );
  AND U23727 ( .A(p_input[32883]), .B(p_input[2883]), .Z(n15817) );
  AND U23728 ( .A(n15819), .B(n15820), .Z(o[2882]) );
  AND U23729 ( .A(p_input[22882]), .B(p_input[12882]), .Z(n15820) );
  AND U23730 ( .A(p_input[32882]), .B(p_input[2882]), .Z(n15819) );
  AND U23731 ( .A(n15821), .B(n15822), .Z(o[2881]) );
  AND U23732 ( .A(p_input[22881]), .B(p_input[12881]), .Z(n15822) );
  AND U23733 ( .A(p_input[32881]), .B(p_input[2881]), .Z(n15821) );
  AND U23734 ( .A(n15823), .B(n15824), .Z(o[2880]) );
  AND U23735 ( .A(p_input[22880]), .B(p_input[12880]), .Z(n15824) );
  AND U23736 ( .A(p_input[32880]), .B(p_input[2880]), .Z(n15823) );
  AND U23737 ( .A(n15825), .B(n15826), .Z(o[287]) );
  AND U23738 ( .A(p_input[20287]), .B(p_input[10287]), .Z(n15826) );
  AND U23739 ( .A(p_input[30287]), .B(p_input[287]), .Z(n15825) );
  AND U23740 ( .A(n15827), .B(n15828), .Z(o[2879]) );
  AND U23741 ( .A(p_input[22879]), .B(p_input[12879]), .Z(n15828) );
  AND U23742 ( .A(p_input[32879]), .B(p_input[2879]), .Z(n15827) );
  AND U23743 ( .A(n15829), .B(n15830), .Z(o[2878]) );
  AND U23744 ( .A(p_input[22878]), .B(p_input[12878]), .Z(n15830) );
  AND U23745 ( .A(p_input[32878]), .B(p_input[2878]), .Z(n15829) );
  AND U23746 ( .A(n15831), .B(n15832), .Z(o[2877]) );
  AND U23747 ( .A(p_input[22877]), .B(p_input[12877]), .Z(n15832) );
  AND U23748 ( .A(p_input[32877]), .B(p_input[2877]), .Z(n15831) );
  AND U23749 ( .A(n15833), .B(n15834), .Z(o[2876]) );
  AND U23750 ( .A(p_input[22876]), .B(p_input[12876]), .Z(n15834) );
  AND U23751 ( .A(p_input[32876]), .B(p_input[2876]), .Z(n15833) );
  AND U23752 ( .A(n15835), .B(n15836), .Z(o[2875]) );
  AND U23753 ( .A(p_input[22875]), .B(p_input[12875]), .Z(n15836) );
  AND U23754 ( .A(p_input[32875]), .B(p_input[2875]), .Z(n15835) );
  AND U23755 ( .A(n15837), .B(n15838), .Z(o[2874]) );
  AND U23756 ( .A(p_input[22874]), .B(p_input[12874]), .Z(n15838) );
  AND U23757 ( .A(p_input[32874]), .B(p_input[2874]), .Z(n15837) );
  AND U23758 ( .A(n15839), .B(n15840), .Z(o[2873]) );
  AND U23759 ( .A(p_input[22873]), .B(p_input[12873]), .Z(n15840) );
  AND U23760 ( .A(p_input[32873]), .B(p_input[2873]), .Z(n15839) );
  AND U23761 ( .A(n15841), .B(n15842), .Z(o[2872]) );
  AND U23762 ( .A(p_input[22872]), .B(p_input[12872]), .Z(n15842) );
  AND U23763 ( .A(p_input[32872]), .B(p_input[2872]), .Z(n15841) );
  AND U23764 ( .A(n15843), .B(n15844), .Z(o[2871]) );
  AND U23765 ( .A(p_input[22871]), .B(p_input[12871]), .Z(n15844) );
  AND U23766 ( .A(p_input[32871]), .B(p_input[2871]), .Z(n15843) );
  AND U23767 ( .A(n15845), .B(n15846), .Z(o[2870]) );
  AND U23768 ( .A(p_input[22870]), .B(p_input[12870]), .Z(n15846) );
  AND U23769 ( .A(p_input[32870]), .B(p_input[2870]), .Z(n15845) );
  AND U23770 ( .A(n15847), .B(n15848), .Z(o[286]) );
  AND U23771 ( .A(p_input[20286]), .B(p_input[10286]), .Z(n15848) );
  AND U23772 ( .A(p_input[30286]), .B(p_input[286]), .Z(n15847) );
  AND U23773 ( .A(n15849), .B(n15850), .Z(o[2869]) );
  AND U23774 ( .A(p_input[22869]), .B(p_input[12869]), .Z(n15850) );
  AND U23775 ( .A(p_input[32869]), .B(p_input[2869]), .Z(n15849) );
  AND U23776 ( .A(n15851), .B(n15852), .Z(o[2868]) );
  AND U23777 ( .A(p_input[22868]), .B(p_input[12868]), .Z(n15852) );
  AND U23778 ( .A(p_input[32868]), .B(p_input[2868]), .Z(n15851) );
  AND U23779 ( .A(n15853), .B(n15854), .Z(o[2867]) );
  AND U23780 ( .A(p_input[22867]), .B(p_input[12867]), .Z(n15854) );
  AND U23781 ( .A(p_input[32867]), .B(p_input[2867]), .Z(n15853) );
  AND U23782 ( .A(n15855), .B(n15856), .Z(o[2866]) );
  AND U23783 ( .A(p_input[22866]), .B(p_input[12866]), .Z(n15856) );
  AND U23784 ( .A(p_input[32866]), .B(p_input[2866]), .Z(n15855) );
  AND U23785 ( .A(n15857), .B(n15858), .Z(o[2865]) );
  AND U23786 ( .A(p_input[22865]), .B(p_input[12865]), .Z(n15858) );
  AND U23787 ( .A(p_input[32865]), .B(p_input[2865]), .Z(n15857) );
  AND U23788 ( .A(n15859), .B(n15860), .Z(o[2864]) );
  AND U23789 ( .A(p_input[22864]), .B(p_input[12864]), .Z(n15860) );
  AND U23790 ( .A(p_input[32864]), .B(p_input[2864]), .Z(n15859) );
  AND U23791 ( .A(n15861), .B(n15862), .Z(o[2863]) );
  AND U23792 ( .A(p_input[22863]), .B(p_input[12863]), .Z(n15862) );
  AND U23793 ( .A(p_input[32863]), .B(p_input[2863]), .Z(n15861) );
  AND U23794 ( .A(n15863), .B(n15864), .Z(o[2862]) );
  AND U23795 ( .A(p_input[22862]), .B(p_input[12862]), .Z(n15864) );
  AND U23796 ( .A(p_input[32862]), .B(p_input[2862]), .Z(n15863) );
  AND U23797 ( .A(n15865), .B(n15866), .Z(o[2861]) );
  AND U23798 ( .A(p_input[22861]), .B(p_input[12861]), .Z(n15866) );
  AND U23799 ( .A(p_input[32861]), .B(p_input[2861]), .Z(n15865) );
  AND U23800 ( .A(n15867), .B(n15868), .Z(o[2860]) );
  AND U23801 ( .A(p_input[22860]), .B(p_input[12860]), .Z(n15868) );
  AND U23802 ( .A(p_input[32860]), .B(p_input[2860]), .Z(n15867) );
  AND U23803 ( .A(n15869), .B(n15870), .Z(o[285]) );
  AND U23804 ( .A(p_input[20285]), .B(p_input[10285]), .Z(n15870) );
  AND U23805 ( .A(p_input[30285]), .B(p_input[285]), .Z(n15869) );
  AND U23806 ( .A(n15871), .B(n15872), .Z(o[2859]) );
  AND U23807 ( .A(p_input[22859]), .B(p_input[12859]), .Z(n15872) );
  AND U23808 ( .A(p_input[32859]), .B(p_input[2859]), .Z(n15871) );
  AND U23809 ( .A(n15873), .B(n15874), .Z(o[2858]) );
  AND U23810 ( .A(p_input[22858]), .B(p_input[12858]), .Z(n15874) );
  AND U23811 ( .A(p_input[32858]), .B(p_input[2858]), .Z(n15873) );
  AND U23812 ( .A(n15875), .B(n15876), .Z(o[2857]) );
  AND U23813 ( .A(p_input[22857]), .B(p_input[12857]), .Z(n15876) );
  AND U23814 ( .A(p_input[32857]), .B(p_input[2857]), .Z(n15875) );
  AND U23815 ( .A(n15877), .B(n15878), .Z(o[2856]) );
  AND U23816 ( .A(p_input[22856]), .B(p_input[12856]), .Z(n15878) );
  AND U23817 ( .A(p_input[32856]), .B(p_input[2856]), .Z(n15877) );
  AND U23818 ( .A(n15879), .B(n15880), .Z(o[2855]) );
  AND U23819 ( .A(p_input[22855]), .B(p_input[12855]), .Z(n15880) );
  AND U23820 ( .A(p_input[32855]), .B(p_input[2855]), .Z(n15879) );
  AND U23821 ( .A(n15881), .B(n15882), .Z(o[2854]) );
  AND U23822 ( .A(p_input[22854]), .B(p_input[12854]), .Z(n15882) );
  AND U23823 ( .A(p_input[32854]), .B(p_input[2854]), .Z(n15881) );
  AND U23824 ( .A(n15883), .B(n15884), .Z(o[2853]) );
  AND U23825 ( .A(p_input[22853]), .B(p_input[12853]), .Z(n15884) );
  AND U23826 ( .A(p_input[32853]), .B(p_input[2853]), .Z(n15883) );
  AND U23827 ( .A(n15885), .B(n15886), .Z(o[2852]) );
  AND U23828 ( .A(p_input[22852]), .B(p_input[12852]), .Z(n15886) );
  AND U23829 ( .A(p_input[32852]), .B(p_input[2852]), .Z(n15885) );
  AND U23830 ( .A(n15887), .B(n15888), .Z(o[2851]) );
  AND U23831 ( .A(p_input[22851]), .B(p_input[12851]), .Z(n15888) );
  AND U23832 ( .A(p_input[32851]), .B(p_input[2851]), .Z(n15887) );
  AND U23833 ( .A(n15889), .B(n15890), .Z(o[2850]) );
  AND U23834 ( .A(p_input[22850]), .B(p_input[12850]), .Z(n15890) );
  AND U23835 ( .A(p_input[32850]), .B(p_input[2850]), .Z(n15889) );
  AND U23836 ( .A(n15891), .B(n15892), .Z(o[284]) );
  AND U23837 ( .A(p_input[20284]), .B(p_input[10284]), .Z(n15892) );
  AND U23838 ( .A(p_input[30284]), .B(p_input[284]), .Z(n15891) );
  AND U23839 ( .A(n15893), .B(n15894), .Z(o[2849]) );
  AND U23840 ( .A(p_input[22849]), .B(p_input[12849]), .Z(n15894) );
  AND U23841 ( .A(p_input[32849]), .B(p_input[2849]), .Z(n15893) );
  AND U23842 ( .A(n15895), .B(n15896), .Z(o[2848]) );
  AND U23843 ( .A(p_input[22848]), .B(p_input[12848]), .Z(n15896) );
  AND U23844 ( .A(p_input[32848]), .B(p_input[2848]), .Z(n15895) );
  AND U23845 ( .A(n15897), .B(n15898), .Z(o[2847]) );
  AND U23846 ( .A(p_input[22847]), .B(p_input[12847]), .Z(n15898) );
  AND U23847 ( .A(p_input[32847]), .B(p_input[2847]), .Z(n15897) );
  AND U23848 ( .A(n15899), .B(n15900), .Z(o[2846]) );
  AND U23849 ( .A(p_input[22846]), .B(p_input[12846]), .Z(n15900) );
  AND U23850 ( .A(p_input[32846]), .B(p_input[2846]), .Z(n15899) );
  AND U23851 ( .A(n15901), .B(n15902), .Z(o[2845]) );
  AND U23852 ( .A(p_input[22845]), .B(p_input[12845]), .Z(n15902) );
  AND U23853 ( .A(p_input[32845]), .B(p_input[2845]), .Z(n15901) );
  AND U23854 ( .A(n15903), .B(n15904), .Z(o[2844]) );
  AND U23855 ( .A(p_input[22844]), .B(p_input[12844]), .Z(n15904) );
  AND U23856 ( .A(p_input[32844]), .B(p_input[2844]), .Z(n15903) );
  AND U23857 ( .A(n15905), .B(n15906), .Z(o[2843]) );
  AND U23858 ( .A(p_input[22843]), .B(p_input[12843]), .Z(n15906) );
  AND U23859 ( .A(p_input[32843]), .B(p_input[2843]), .Z(n15905) );
  AND U23860 ( .A(n15907), .B(n15908), .Z(o[2842]) );
  AND U23861 ( .A(p_input[22842]), .B(p_input[12842]), .Z(n15908) );
  AND U23862 ( .A(p_input[32842]), .B(p_input[2842]), .Z(n15907) );
  AND U23863 ( .A(n15909), .B(n15910), .Z(o[2841]) );
  AND U23864 ( .A(p_input[22841]), .B(p_input[12841]), .Z(n15910) );
  AND U23865 ( .A(p_input[32841]), .B(p_input[2841]), .Z(n15909) );
  AND U23866 ( .A(n15911), .B(n15912), .Z(o[2840]) );
  AND U23867 ( .A(p_input[22840]), .B(p_input[12840]), .Z(n15912) );
  AND U23868 ( .A(p_input[32840]), .B(p_input[2840]), .Z(n15911) );
  AND U23869 ( .A(n15913), .B(n15914), .Z(o[283]) );
  AND U23870 ( .A(p_input[20283]), .B(p_input[10283]), .Z(n15914) );
  AND U23871 ( .A(p_input[30283]), .B(p_input[283]), .Z(n15913) );
  AND U23872 ( .A(n15915), .B(n15916), .Z(o[2839]) );
  AND U23873 ( .A(p_input[22839]), .B(p_input[12839]), .Z(n15916) );
  AND U23874 ( .A(p_input[32839]), .B(p_input[2839]), .Z(n15915) );
  AND U23875 ( .A(n15917), .B(n15918), .Z(o[2838]) );
  AND U23876 ( .A(p_input[22838]), .B(p_input[12838]), .Z(n15918) );
  AND U23877 ( .A(p_input[32838]), .B(p_input[2838]), .Z(n15917) );
  AND U23878 ( .A(n15919), .B(n15920), .Z(o[2837]) );
  AND U23879 ( .A(p_input[22837]), .B(p_input[12837]), .Z(n15920) );
  AND U23880 ( .A(p_input[32837]), .B(p_input[2837]), .Z(n15919) );
  AND U23881 ( .A(n15921), .B(n15922), .Z(o[2836]) );
  AND U23882 ( .A(p_input[22836]), .B(p_input[12836]), .Z(n15922) );
  AND U23883 ( .A(p_input[32836]), .B(p_input[2836]), .Z(n15921) );
  AND U23884 ( .A(n15923), .B(n15924), .Z(o[2835]) );
  AND U23885 ( .A(p_input[22835]), .B(p_input[12835]), .Z(n15924) );
  AND U23886 ( .A(p_input[32835]), .B(p_input[2835]), .Z(n15923) );
  AND U23887 ( .A(n15925), .B(n15926), .Z(o[2834]) );
  AND U23888 ( .A(p_input[22834]), .B(p_input[12834]), .Z(n15926) );
  AND U23889 ( .A(p_input[32834]), .B(p_input[2834]), .Z(n15925) );
  AND U23890 ( .A(n15927), .B(n15928), .Z(o[2833]) );
  AND U23891 ( .A(p_input[22833]), .B(p_input[12833]), .Z(n15928) );
  AND U23892 ( .A(p_input[32833]), .B(p_input[2833]), .Z(n15927) );
  AND U23893 ( .A(n15929), .B(n15930), .Z(o[2832]) );
  AND U23894 ( .A(p_input[22832]), .B(p_input[12832]), .Z(n15930) );
  AND U23895 ( .A(p_input[32832]), .B(p_input[2832]), .Z(n15929) );
  AND U23896 ( .A(n15931), .B(n15932), .Z(o[2831]) );
  AND U23897 ( .A(p_input[22831]), .B(p_input[12831]), .Z(n15932) );
  AND U23898 ( .A(p_input[32831]), .B(p_input[2831]), .Z(n15931) );
  AND U23899 ( .A(n15933), .B(n15934), .Z(o[2830]) );
  AND U23900 ( .A(p_input[22830]), .B(p_input[12830]), .Z(n15934) );
  AND U23901 ( .A(p_input[32830]), .B(p_input[2830]), .Z(n15933) );
  AND U23902 ( .A(n15935), .B(n15936), .Z(o[282]) );
  AND U23903 ( .A(p_input[20282]), .B(p_input[10282]), .Z(n15936) );
  AND U23904 ( .A(p_input[30282]), .B(p_input[282]), .Z(n15935) );
  AND U23905 ( .A(n15937), .B(n15938), .Z(o[2829]) );
  AND U23906 ( .A(p_input[22829]), .B(p_input[12829]), .Z(n15938) );
  AND U23907 ( .A(p_input[32829]), .B(p_input[2829]), .Z(n15937) );
  AND U23908 ( .A(n15939), .B(n15940), .Z(o[2828]) );
  AND U23909 ( .A(p_input[22828]), .B(p_input[12828]), .Z(n15940) );
  AND U23910 ( .A(p_input[32828]), .B(p_input[2828]), .Z(n15939) );
  AND U23911 ( .A(n15941), .B(n15942), .Z(o[2827]) );
  AND U23912 ( .A(p_input[22827]), .B(p_input[12827]), .Z(n15942) );
  AND U23913 ( .A(p_input[32827]), .B(p_input[2827]), .Z(n15941) );
  AND U23914 ( .A(n15943), .B(n15944), .Z(o[2826]) );
  AND U23915 ( .A(p_input[22826]), .B(p_input[12826]), .Z(n15944) );
  AND U23916 ( .A(p_input[32826]), .B(p_input[2826]), .Z(n15943) );
  AND U23917 ( .A(n15945), .B(n15946), .Z(o[2825]) );
  AND U23918 ( .A(p_input[22825]), .B(p_input[12825]), .Z(n15946) );
  AND U23919 ( .A(p_input[32825]), .B(p_input[2825]), .Z(n15945) );
  AND U23920 ( .A(n15947), .B(n15948), .Z(o[2824]) );
  AND U23921 ( .A(p_input[22824]), .B(p_input[12824]), .Z(n15948) );
  AND U23922 ( .A(p_input[32824]), .B(p_input[2824]), .Z(n15947) );
  AND U23923 ( .A(n15949), .B(n15950), .Z(o[2823]) );
  AND U23924 ( .A(p_input[22823]), .B(p_input[12823]), .Z(n15950) );
  AND U23925 ( .A(p_input[32823]), .B(p_input[2823]), .Z(n15949) );
  AND U23926 ( .A(n15951), .B(n15952), .Z(o[2822]) );
  AND U23927 ( .A(p_input[22822]), .B(p_input[12822]), .Z(n15952) );
  AND U23928 ( .A(p_input[32822]), .B(p_input[2822]), .Z(n15951) );
  AND U23929 ( .A(n15953), .B(n15954), .Z(o[2821]) );
  AND U23930 ( .A(p_input[22821]), .B(p_input[12821]), .Z(n15954) );
  AND U23931 ( .A(p_input[32821]), .B(p_input[2821]), .Z(n15953) );
  AND U23932 ( .A(n15955), .B(n15956), .Z(o[2820]) );
  AND U23933 ( .A(p_input[22820]), .B(p_input[12820]), .Z(n15956) );
  AND U23934 ( .A(p_input[32820]), .B(p_input[2820]), .Z(n15955) );
  AND U23935 ( .A(n15957), .B(n15958), .Z(o[281]) );
  AND U23936 ( .A(p_input[20281]), .B(p_input[10281]), .Z(n15958) );
  AND U23937 ( .A(p_input[30281]), .B(p_input[281]), .Z(n15957) );
  AND U23938 ( .A(n15959), .B(n15960), .Z(o[2819]) );
  AND U23939 ( .A(p_input[22819]), .B(p_input[12819]), .Z(n15960) );
  AND U23940 ( .A(p_input[32819]), .B(p_input[2819]), .Z(n15959) );
  AND U23941 ( .A(n15961), .B(n15962), .Z(o[2818]) );
  AND U23942 ( .A(p_input[22818]), .B(p_input[12818]), .Z(n15962) );
  AND U23943 ( .A(p_input[32818]), .B(p_input[2818]), .Z(n15961) );
  AND U23944 ( .A(n15963), .B(n15964), .Z(o[2817]) );
  AND U23945 ( .A(p_input[22817]), .B(p_input[12817]), .Z(n15964) );
  AND U23946 ( .A(p_input[32817]), .B(p_input[2817]), .Z(n15963) );
  AND U23947 ( .A(n15965), .B(n15966), .Z(o[2816]) );
  AND U23948 ( .A(p_input[22816]), .B(p_input[12816]), .Z(n15966) );
  AND U23949 ( .A(p_input[32816]), .B(p_input[2816]), .Z(n15965) );
  AND U23950 ( .A(n15967), .B(n15968), .Z(o[2815]) );
  AND U23951 ( .A(p_input[22815]), .B(p_input[12815]), .Z(n15968) );
  AND U23952 ( .A(p_input[32815]), .B(p_input[2815]), .Z(n15967) );
  AND U23953 ( .A(n15969), .B(n15970), .Z(o[2814]) );
  AND U23954 ( .A(p_input[22814]), .B(p_input[12814]), .Z(n15970) );
  AND U23955 ( .A(p_input[32814]), .B(p_input[2814]), .Z(n15969) );
  AND U23956 ( .A(n15971), .B(n15972), .Z(o[2813]) );
  AND U23957 ( .A(p_input[22813]), .B(p_input[12813]), .Z(n15972) );
  AND U23958 ( .A(p_input[32813]), .B(p_input[2813]), .Z(n15971) );
  AND U23959 ( .A(n15973), .B(n15974), .Z(o[2812]) );
  AND U23960 ( .A(p_input[22812]), .B(p_input[12812]), .Z(n15974) );
  AND U23961 ( .A(p_input[32812]), .B(p_input[2812]), .Z(n15973) );
  AND U23962 ( .A(n15975), .B(n15976), .Z(o[2811]) );
  AND U23963 ( .A(p_input[22811]), .B(p_input[12811]), .Z(n15976) );
  AND U23964 ( .A(p_input[32811]), .B(p_input[2811]), .Z(n15975) );
  AND U23965 ( .A(n15977), .B(n15978), .Z(o[2810]) );
  AND U23966 ( .A(p_input[22810]), .B(p_input[12810]), .Z(n15978) );
  AND U23967 ( .A(p_input[32810]), .B(p_input[2810]), .Z(n15977) );
  AND U23968 ( .A(n15979), .B(n15980), .Z(o[280]) );
  AND U23969 ( .A(p_input[20280]), .B(p_input[10280]), .Z(n15980) );
  AND U23970 ( .A(p_input[30280]), .B(p_input[280]), .Z(n15979) );
  AND U23971 ( .A(n15981), .B(n15982), .Z(o[2809]) );
  AND U23972 ( .A(p_input[22809]), .B(p_input[12809]), .Z(n15982) );
  AND U23973 ( .A(p_input[32809]), .B(p_input[2809]), .Z(n15981) );
  AND U23974 ( .A(n15983), .B(n15984), .Z(o[2808]) );
  AND U23975 ( .A(p_input[22808]), .B(p_input[12808]), .Z(n15984) );
  AND U23976 ( .A(p_input[32808]), .B(p_input[2808]), .Z(n15983) );
  AND U23977 ( .A(n15985), .B(n15986), .Z(o[2807]) );
  AND U23978 ( .A(p_input[22807]), .B(p_input[12807]), .Z(n15986) );
  AND U23979 ( .A(p_input[32807]), .B(p_input[2807]), .Z(n15985) );
  AND U23980 ( .A(n15987), .B(n15988), .Z(o[2806]) );
  AND U23981 ( .A(p_input[22806]), .B(p_input[12806]), .Z(n15988) );
  AND U23982 ( .A(p_input[32806]), .B(p_input[2806]), .Z(n15987) );
  AND U23983 ( .A(n15989), .B(n15990), .Z(o[2805]) );
  AND U23984 ( .A(p_input[22805]), .B(p_input[12805]), .Z(n15990) );
  AND U23985 ( .A(p_input[32805]), .B(p_input[2805]), .Z(n15989) );
  AND U23986 ( .A(n15991), .B(n15992), .Z(o[2804]) );
  AND U23987 ( .A(p_input[22804]), .B(p_input[12804]), .Z(n15992) );
  AND U23988 ( .A(p_input[32804]), .B(p_input[2804]), .Z(n15991) );
  AND U23989 ( .A(n15993), .B(n15994), .Z(o[2803]) );
  AND U23990 ( .A(p_input[22803]), .B(p_input[12803]), .Z(n15994) );
  AND U23991 ( .A(p_input[32803]), .B(p_input[2803]), .Z(n15993) );
  AND U23992 ( .A(n15995), .B(n15996), .Z(o[2802]) );
  AND U23993 ( .A(p_input[22802]), .B(p_input[12802]), .Z(n15996) );
  AND U23994 ( .A(p_input[32802]), .B(p_input[2802]), .Z(n15995) );
  AND U23995 ( .A(n15997), .B(n15998), .Z(o[2801]) );
  AND U23996 ( .A(p_input[22801]), .B(p_input[12801]), .Z(n15998) );
  AND U23997 ( .A(p_input[32801]), .B(p_input[2801]), .Z(n15997) );
  AND U23998 ( .A(n15999), .B(n16000), .Z(o[2800]) );
  AND U23999 ( .A(p_input[22800]), .B(p_input[12800]), .Z(n16000) );
  AND U24000 ( .A(p_input[32800]), .B(p_input[2800]), .Z(n15999) );
  AND U24001 ( .A(n16001), .B(n16002), .Z(o[27]) );
  AND U24002 ( .A(p_input[20027]), .B(p_input[10027]), .Z(n16002) );
  AND U24003 ( .A(p_input[30027]), .B(p_input[27]), .Z(n16001) );
  AND U24004 ( .A(n16003), .B(n16004), .Z(o[279]) );
  AND U24005 ( .A(p_input[20279]), .B(p_input[10279]), .Z(n16004) );
  AND U24006 ( .A(p_input[30279]), .B(p_input[279]), .Z(n16003) );
  AND U24007 ( .A(n16005), .B(n16006), .Z(o[2799]) );
  AND U24008 ( .A(p_input[22799]), .B(p_input[12799]), .Z(n16006) );
  AND U24009 ( .A(p_input[32799]), .B(p_input[2799]), .Z(n16005) );
  AND U24010 ( .A(n16007), .B(n16008), .Z(o[2798]) );
  AND U24011 ( .A(p_input[22798]), .B(p_input[12798]), .Z(n16008) );
  AND U24012 ( .A(p_input[32798]), .B(p_input[2798]), .Z(n16007) );
  AND U24013 ( .A(n16009), .B(n16010), .Z(o[2797]) );
  AND U24014 ( .A(p_input[22797]), .B(p_input[12797]), .Z(n16010) );
  AND U24015 ( .A(p_input[32797]), .B(p_input[2797]), .Z(n16009) );
  AND U24016 ( .A(n16011), .B(n16012), .Z(o[2796]) );
  AND U24017 ( .A(p_input[22796]), .B(p_input[12796]), .Z(n16012) );
  AND U24018 ( .A(p_input[32796]), .B(p_input[2796]), .Z(n16011) );
  AND U24019 ( .A(n16013), .B(n16014), .Z(o[2795]) );
  AND U24020 ( .A(p_input[22795]), .B(p_input[12795]), .Z(n16014) );
  AND U24021 ( .A(p_input[32795]), .B(p_input[2795]), .Z(n16013) );
  AND U24022 ( .A(n16015), .B(n16016), .Z(o[2794]) );
  AND U24023 ( .A(p_input[22794]), .B(p_input[12794]), .Z(n16016) );
  AND U24024 ( .A(p_input[32794]), .B(p_input[2794]), .Z(n16015) );
  AND U24025 ( .A(n16017), .B(n16018), .Z(o[2793]) );
  AND U24026 ( .A(p_input[22793]), .B(p_input[12793]), .Z(n16018) );
  AND U24027 ( .A(p_input[32793]), .B(p_input[2793]), .Z(n16017) );
  AND U24028 ( .A(n16019), .B(n16020), .Z(o[2792]) );
  AND U24029 ( .A(p_input[22792]), .B(p_input[12792]), .Z(n16020) );
  AND U24030 ( .A(p_input[32792]), .B(p_input[2792]), .Z(n16019) );
  AND U24031 ( .A(n16021), .B(n16022), .Z(o[2791]) );
  AND U24032 ( .A(p_input[22791]), .B(p_input[12791]), .Z(n16022) );
  AND U24033 ( .A(p_input[32791]), .B(p_input[2791]), .Z(n16021) );
  AND U24034 ( .A(n16023), .B(n16024), .Z(o[2790]) );
  AND U24035 ( .A(p_input[22790]), .B(p_input[12790]), .Z(n16024) );
  AND U24036 ( .A(p_input[32790]), .B(p_input[2790]), .Z(n16023) );
  AND U24037 ( .A(n16025), .B(n16026), .Z(o[278]) );
  AND U24038 ( .A(p_input[20278]), .B(p_input[10278]), .Z(n16026) );
  AND U24039 ( .A(p_input[30278]), .B(p_input[278]), .Z(n16025) );
  AND U24040 ( .A(n16027), .B(n16028), .Z(o[2789]) );
  AND U24041 ( .A(p_input[22789]), .B(p_input[12789]), .Z(n16028) );
  AND U24042 ( .A(p_input[32789]), .B(p_input[2789]), .Z(n16027) );
  AND U24043 ( .A(n16029), .B(n16030), .Z(o[2788]) );
  AND U24044 ( .A(p_input[22788]), .B(p_input[12788]), .Z(n16030) );
  AND U24045 ( .A(p_input[32788]), .B(p_input[2788]), .Z(n16029) );
  AND U24046 ( .A(n16031), .B(n16032), .Z(o[2787]) );
  AND U24047 ( .A(p_input[22787]), .B(p_input[12787]), .Z(n16032) );
  AND U24048 ( .A(p_input[32787]), .B(p_input[2787]), .Z(n16031) );
  AND U24049 ( .A(n16033), .B(n16034), .Z(o[2786]) );
  AND U24050 ( .A(p_input[22786]), .B(p_input[12786]), .Z(n16034) );
  AND U24051 ( .A(p_input[32786]), .B(p_input[2786]), .Z(n16033) );
  AND U24052 ( .A(n16035), .B(n16036), .Z(o[2785]) );
  AND U24053 ( .A(p_input[22785]), .B(p_input[12785]), .Z(n16036) );
  AND U24054 ( .A(p_input[32785]), .B(p_input[2785]), .Z(n16035) );
  AND U24055 ( .A(n16037), .B(n16038), .Z(o[2784]) );
  AND U24056 ( .A(p_input[22784]), .B(p_input[12784]), .Z(n16038) );
  AND U24057 ( .A(p_input[32784]), .B(p_input[2784]), .Z(n16037) );
  AND U24058 ( .A(n16039), .B(n16040), .Z(o[2783]) );
  AND U24059 ( .A(p_input[22783]), .B(p_input[12783]), .Z(n16040) );
  AND U24060 ( .A(p_input[32783]), .B(p_input[2783]), .Z(n16039) );
  AND U24061 ( .A(n16041), .B(n16042), .Z(o[2782]) );
  AND U24062 ( .A(p_input[22782]), .B(p_input[12782]), .Z(n16042) );
  AND U24063 ( .A(p_input[32782]), .B(p_input[2782]), .Z(n16041) );
  AND U24064 ( .A(n16043), .B(n16044), .Z(o[2781]) );
  AND U24065 ( .A(p_input[22781]), .B(p_input[12781]), .Z(n16044) );
  AND U24066 ( .A(p_input[32781]), .B(p_input[2781]), .Z(n16043) );
  AND U24067 ( .A(n16045), .B(n16046), .Z(o[2780]) );
  AND U24068 ( .A(p_input[22780]), .B(p_input[12780]), .Z(n16046) );
  AND U24069 ( .A(p_input[32780]), .B(p_input[2780]), .Z(n16045) );
  AND U24070 ( .A(n16047), .B(n16048), .Z(o[277]) );
  AND U24071 ( .A(p_input[20277]), .B(p_input[10277]), .Z(n16048) );
  AND U24072 ( .A(p_input[30277]), .B(p_input[277]), .Z(n16047) );
  AND U24073 ( .A(n16049), .B(n16050), .Z(o[2779]) );
  AND U24074 ( .A(p_input[22779]), .B(p_input[12779]), .Z(n16050) );
  AND U24075 ( .A(p_input[32779]), .B(p_input[2779]), .Z(n16049) );
  AND U24076 ( .A(n16051), .B(n16052), .Z(o[2778]) );
  AND U24077 ( .A(p_input[22778]), .B(p_input[12778]), .Z(n16052) );
  AND U24078 ( .A(p_input[32778]), .B(p_input[2778]), .Z(n16051) );
  AND U24079 ( .A(n16053), .B(n16054), .Z(o[2777]) );
  AND U24080 ( .A(p_input[22777]), .B(p_input[12777]), .Z(n16054) );
  AND U24081 ( .A(p_input[32777]), .B(p_input[2777]), .Z(n16053) );
  AND U24082 ( .A(n16055), .B(n16056), .Z(o[2776]) );
  AND U24083 ( .A(p_input[22776]), .B(p_input[12776]), .Z(n16056) );
  AND U24084 ( .A(p_input[32776]), .B(p_input[2776]), .Z(n16055) );
  AND U24085 ( .A(n16057), .B(n16058), .Z(o[2775]) );
  AND U24086 ( .A(p_input[22775]), .B(p_input[12775]), .Z(n16058) );
  AND U24087 ( .A(p_input[32775]), .B(p_input[2775]), .Z(n16057) );
  AND U24088 ( .A(n16059), .B(n16060), .Z(o[2774]) );
  AND U24089 ( .A(p_input[22774]), .B(p_input[12774]), .Z(n16060) );
  AND U24090 ( .A(p_input[32774]), .B(p_input[2774]), .Z(n16059) );
  AND U24091 ( .A(n16061), .B(n16062), .Z(o[2773]) );
  AND U24092 ( .A(p_input[22773]), .B(p_input[12773]), .Z(n16062) );
  AND U24093 ( .A(p_input[32773]), .B(p_input[2773]), .Z(n16061) );
  AND U24094 ( .A(n16063), .B(n16064), .Z(o[2772]) );
  AND U24095 ( .A(p_input[22772]), .B(p_input[12772]), .Z(n16064) );
  AND U24096 ( .A(p_input[32772]), .B(p_input[2772]), .Z(n16063) );
  AND U24097 ( .A(n16065), .B(n16066), .Z(o[2771]) );
  AND U24098 ( .A(p_input[22771]), .B(p_input[12771]), .Z(n16066) );
  AND U24099 ( .A(p_input[32771]), .B(p_input[2771]), .Z(n16065) );
  AND U24100 ( .A(n16067), .B(n16068), .Z(o[2770]) );
  AND U24101 ( .A(p_input[22770]), .B(p_input[12770]), .Z(n16068) );
  AND U24102 ( .A(p_input[32770]), .B(p_input[2770]), .Z(n16067) );
  AND U24103 ( .A(n16069), .B(n16070), .Z(o[276]) );
  AND U24104 ( .A(p_input[20276]), .B(p_input[10276]), .Z(n16070) );
  AND U24105 ( .A(p_input[30276]), .B(p_input[276]), .Z(n16069) );
  AND U24106 ( .A(n16071), .B(n16072), .Z(o[2769]) );
  AND U24107 ( .A(p_input[22769]), .B(p_input[12769]), .Z(n16072) );
  AND U24108 ( .A(p_input[32769]), .B(p_input[2769]), .Z(n16071) );
  AND U24109 ( .A(n16073), .B(n16074), .Z(o[2768]) );
  AND U24110 ( .A(p_input[22768]), .B(p_input[12768]), .Z(n16074) );
  AND U24111 ( .A(p_input[32768]), .B(p_input[2768]), .Z(n16073) );
  AND U24112 ( .A(n16075), .B(n16076), .Z(o[2767]) );
  AND U24113 ( .A(p_input[22767]), .B(p_input[12767]), .Z(n16076) );
  AND U24114 ( .A(p_input[32767]), .B(p_input[2767]), .Z(n16075) );
  AND U24115 ( .A(n16077), .B(n16078), .Z(o[2766]) );
  AND U24116 ( .A(p_input[22766]), .B(p_input[12766]), .Z(n16078) );
  AND U24117 ( .A(p_input[32766]), .B(p_input[2766]), .Z(n16077) );
  AND U24118 ( .A(n16079), .B(n16080), .Z(o[2765]) );
  AND U24119 ( .A(p_input[22765]), .B(p_input[12765]), .Z(n16080) );
  AND U24120 ( .A(p_input[32765]), .B(p_input[2765]), .Z(n16079) );
  AND U24121 ( .A(n16081), .B(n16082), .Z(o[2764]) );
  AND U24122 ( .A(p_input[22764]), .B(p_input[12764]), .Z(n16082) );
  AND U24123 ( .A(p_input[32764]), .B(p_input[2764]), .Z(n16081) );
  AND U24124 ( .A(n16083), .B(n16084), .Z(o[2763]) );
  AND U24125 ( .A(p_input[22763]), .B(p_input[12763]), .Z(n16084) );
  AND U24126 ( .A(p_input[32763]), .B(p_input[2763]), .Z(n16083) );
  AND U24127 ( .A(n16085), .B(n16086), .Z(o[2762]) );
  AND U24128 ( .A(p_input[22762]), .B(p_input[12762]), .Z(n16086) );
  AND U24129 ( .A(p_input[32762]), .B(p_input[2762]), .Z(n16085) );
  AND U24130 ( .A(n16087), .B(n16088), .Z(o[2761]) );
  AND U24131 ( .A(p_input[22761]), .B(p_input[12761]), .Z(n16088) );
  AND U24132 ( .A(p_input[32761]), .B(p_input[2761]), .Z(n16087) );
  AND U24133 ( .A(n16089), .B(n16090), .Z(o[2760]) );
  AND U24134 ( .A(p_input[22760]), .B(p_input[12760]), .Z(n16090) );
  AND U24135 ( .A(p_input[32760]), .B(p_input[2760]), .Z(n16089) );
  AND U24136 ( .A(n16091), .B(n16092), .Z(o[275]) );
  AND U24137 ( .A(p_input[20275]), .B(p_input[10275]), .Z(n16092) );
  AND U24138 ( .A(p_input[30275]), .B(p_input[275]), .Z(n16091) );
  AND U24139 ( .A(n16093), .B(n16094), .Z(o[2759]) );
  AND U24140 ( .A(p_input[22759]), .B(p_input[12759]), .Z(n16094) );
  AND U24141 ( .A(p_input[32759]), .B(p_input[2759]), .Z(n16093) );
  AND U24142 ( .A(n16095), .B(n16096), .Z(o[2758]) );
  AND U24143 ( .A(p_input[22758]), .B(p_input[12758]), .Z(n16096) );
  AND U24144 ( .A(p_input[32758]), .B(p_input[2758]), .Z(n16095) );
  AND U24145 ( .A(n16097), .B(n16098), .Z(o[2757]) );
  AND U24146 ( .A(p_input[22757]), .B(p_input[12757]), .Z(n16098) );
  AND U24147 ( .A(p_input[32757]), .B(p_input[2757]), .Z(n16097) );
  AND U24148 ( .A(n16099), .B(n16100), .Z(o[2756]) );
  AND U24149 ( .A(p_input[22756]), .B(p_input[12756]), .Z(n16100) );
  AND U24150 ( .A(p_input[32756]), .B(p_input[2756]), .Z(n16099) );
  AND U24151 ( .A(n16101), .B(n16102), .Z(o[2755]) );
  AND U24152 ( .A(p_input[22755]), .B(p_input[12755]), .Z(n16102) );
  AND U24153 ( .A(p_input[32755]), .B(p_input[2755]), .Z(n16101) );
  AND U24154 ( .A(n16103), .B(n16104), .Z(o[2754]) );
  AND U24155 ( .A(p_input[22754]), .B(p_input[12754]), .Z(n16104) );
  AND U24156 ( .A(p_input[32754]), .B(p_input[2754]), .Z(n16103) );
  AND U24157 ( .A(n16105), .B(n16106), .Z(o[2753]) );
  AND U24158 ( .A(p_input[22753]), .B(p_input[12753]), .Z(n16106) );
  AND U24159 ( .A(p_input[32753]), .B(p_input[2753]), .Z(n16105) );
  AND U24160 ( .A(n16107), .B(n16108), .Z(o[2752]) );
  AND U24161 ( .A(p_input[22752]), .B(p_input[12752]), .Z(n16108) );
  AND U24162 ( .A(p_input[32752]), .B(p_input[2752]), .Z(n16107) );
  AND U24163 ( .A(n16109), .B(n16110), .Z(o[2751]) );
  AND U24164 ( .A(p_input[22751]), .B(p_input[12751]), .Z(n16110) );
  AND U24165 ( .A(p_input[32751]), .B(p_input[2751]), .Z(n16109) );
  AND U24166 ( .A(n16111), .B(n16112), .Z(o[2750]) );
  AND U24167 ( .A(p_input[22750]), .B(p_input[12750]), .Z(n16112) );
  AND U24168 ( .A(p_input[32750]), .B(p_input[2750]), .Z(n16111) );
  AND U24169 ( .A(n16113), .B(n16114), .Z(o[274]) );
  AND U24170 ( .A(p_input[20274]), .B(p_input[10274]), .Z(n16114) );
  AND U24171 ( .A(p_input[30274]), .B(p_input[274]), .Z(n16113) );
  AND U24172 ( .A(n16115), .B(n16116), .Z(o[2749]) );
  AND U24173 ( .A(p_input[22749]), .B(p_input[12749]), .Z(n16116) );
  AND U24174 ( .A(p_input[32749]), .B(p_input[2749]), .Z(n16115) );
  AND U24175 ( .A(n16117), .B(n16118), .Z(o[2748]) );
  AND U24176 ( .A(p_input[22748]), .B(p_input[12748]), .Z(n16118) );
  AND U24177 ( .A(p_input[32748]), .B(p_input[2748]), .Z(n16117) );
  AND U24178 ( .A(n16119), .B(n16120), .Z(o[2747]) );
  AND U24179 ( .A(p_input[22747]), .B(p_input[12747]), .Z(n16120) );
  AND U24180 ( .A(p_input[32747]), .B(p_input[2747]), .Z(n16119) );
  AND U24181 ( .A(n16121), .B(n16122), .Z(o[2746]) );
  AND U24182 ( .A(p_input[22746]), .B(p_input[12746]), .Z(n16122) );
  AND U24183 ( .A(p_input[32746]), .B(p_input[2746]), .Z(n16121) );
  AND U24184 ( .A(n16123), .B(n16124), .Z(o[2745]) );
  AND U24185 ( .A(p_input[22745]), .B(p_input[12745]), .Z(n16124) );
  AND U24186 ( .A(p_input[32745]), .B(p_input[2745]), .Z(n16123) );
  AND U24187 ( .A(n16125), .B(n16126), .Z(o[2744]) );
  AND U24188 ( .A(p_input[22744]), .B(p_input[12744]), .Z(n16126) );
  AND U24189 ( .A(p_input[32744]), .B(p_input[2744]), .Z(n16125) );
  AND U24190 ( .A(n16127), .B(n16128), .Z(o[2743]) );
  AND U24191 ( .A(p_input[22743]), .B(p_input[12743]), .Z(n16128) );
  AND U24192 ( .A(p_input[32743]), .B(p_input[2743]), .Z(n16127) );
  AND U24193 ( .A(n16129), .B(n16130), .Z(o[2742]) );
  AND U24194 ( .A(p_input[22742]), .B(p_input[12742]), .Z(n16130) );
  AND U24195 ( .A(p_input[32742]), .B(p_input[2742]), .Z(n16129) );
  AND U24196 ( .A(n16131), .B(n16132), .Z(o[2741]) );
  AND U24197 ( .A(p_input[22741]), .B(p_input[12741]), .Z(n16132) );
  AND U24198 ( .A(p_input[32741]), .B(p_input[2741]), .Z(n16131) );
  AND U24199 ( .A(n16133), .B(n16134), .Z(o[2740]) );
  AND U24200 ( .A(p_input[22740]), .B(p_input[12740]), .Z(n16134) );
  AND U24201 ( .A(p_input[32740]), .B(p_input[2740]), .Z(n16133) );
  AND U24202 ( .A(n16135), .B(n16136), .Z(o[273]) );
  AND U24203 ( .A(p_input[20273]), .B(p_input[10273]), .Z(n16136) );
  AND U24204 ( .A(p_input[30273]), .B(p_input[273]), .Z(n16135) );
  AND U24205 ( .A(n16137), .B(n16138), .Z(o[2739]) );
  AND U24206 ( .A(p_input[22739]), .B(p_input[12739]), .Z(n16138) );
  AND U24207 ( .A(p_input[32739]), .B(p_input[2739]), .Z(n16137) );
  AND U24208 ( .A(n16139), .B(n16140), .Z(o[2738]) );
  AND U24209 ( .A(p_input[22738]), .B(p_input[12738]), .Z(n16140) );
  AND U24210 ( .A(p_input[32738]), .B(p_input[2738]), .Z(n16139) );
  AND U24211 ( .A(n16141), .B(n16142), .Z(o[2737]) );
  AND U24212 ( .A(p_input[22737]), .B(p_input[12737]), .Z(n16142) );
  AND U24213 ( .A(p_input[32737]), .B(p_input[2737]), .Z(n16141) );
  AND U24214 ( .A(n16143), .B(n16144), .Z(o[2736]) );
  AND U24215 ( .A(p_input[22736]), .B(p_input[12736]), .Z(n16144) );
  AND U24216 ( .A(p_input[32736]), .B(p_input[2736]), .Z(n16143) );
  AND U24217 ( .A(n16145), .B(n16146), .Z(o[2735]) );
  AND U24218 ( .A(p_input[22735]), .B(p_input[12735]), .Z(n16146) );
  AND U24219 ( .A(p_input[32735]), .B(p_input[2735]), .Z(n16145) );
  AND U24220 ( .A(n16147), .B(n16148), .Z(o[2734]) );
  AND U24221 ( .A(p_input[22734]), .B(p_input[12734]), .Z(n16148) );
  AND U24222 ( .A(p_input[32734]), .B(p_input[2734]), .Z(n16147) );
  AND U24223 ( .A(n16149), .B(n16150), .Z(o[2733]) );
  AND U24224 ( .A(p_input[22733]), .B(p_input[12733]), .Z(n16150) );
  AND U24225 ( .A(p_input[32733]), .B(p_input[2733]), .Z(n16149) );
  AND U24226 ( .A(n16151), .B(n16152), .Z(o[2732]) );
  AND U24227 ( .A(p_input[22732]), .B(p_input[12732]), .Z(n16152) );
  AND U24228 ( .A(p_input[32732]), .B(p_input[2732]), .Z(n16151) );
  AND U24229 ( .A(n16153), .B(n16154), .Z(o[2731]) );
  AND U24230 ( .A(p_input[22731]), .B(p_input[12731]), .Z(n16154) );
  AND U24231 ( .A(p_input[32731]), .B(p_input[2731]), .Z(n16153) );
  AND U24232 ( .A(n16155), .B(n16156), .Z(o[2730]) );
  AND U24233 ( .A(p_input[22730]), .B(p_input[12730]), .Z(n16156) );
  AND U24234 ( .A(p_input[32730]), .B(p_input[2730]), .Z(n16155) );
  AND U24235 ( .A(n16157), .B(n16158), .Z(o[272]) );
  AND U24236 ( .A(p_input[20272]), .B(p_input[10272]), .Z(n16158) );
  AND U24237 ( .A(p_input[30272]), .B(p_input[272]), .Z(n16157) );
  AND U24238 ( .A(n16159), .B(n16160), .Z(o[2729]) );
  AND U24239 ( .A(p_input[22729]), .B(p_input[12729]), .Z(n16160) );
  AND U24240 ( .A(p_input[32729]), .B(p_input[2729]), .Z(n16159) );
  AND U24241 ( .A(n16161), .B(n16162), .Z(o[2728]) );
  AND U24242 ( .A(p_input[22728]), .B(p_input[12728]), .Z(n16162) );
  AND U24243 ( .A(p_input[32728]), .B(p_input[2728]), .Z(n16161) );
  AND U24244 ( .A(n16163), .B(n16164), .Z(o[2727]) );
  AND U24245 ( .A(p_input[22727]), .B(p_input[12727]), .Z(n16164) );
  AND U24246 ( .A(p_input[32727]), .B(p_input[2727]), .Z(n16163) );
  AND U24247 ( .A(n16165), .B(n16166), .Z(o[2726]) );
  AND U24248 ( .A(p_input[22726]), .B(p_input[12726]), .Z(n16166) );
  AND U24249 ( .A(p_input[32726]), .B(p_input[2726]), .Z(n16165) );
  AND U24250 ( .A(n16167), .B(n16168), .Z(o[2725]) );
  AND U24251 ( .A(p_input[22725]), .B(p_input[12725]), .Z(n16168) );
  AND U24252 ( .A(p_input[32725]), .B(p_input[2725]), .Z(n16167) );
  AND U24253 ( .A(n16169), .B(n16170), .Z(o[2724]) );
  AND U24254 ( .A(p_input[22724]), .B(p_input[12724]), .Z(n16170) );
  AND U24255 ( .A(p_input[32724]), .B(p_input[2724]), .Z(n16169) );
  AND U24256 ( .A(n16171), .B(n16172), .Z(o[2723]) );
  AND U24257 ( .A(p_input[22723]), .B(p_input[12723]), .Z(n16172) );
  AND U24258 ( .A(p_input[32723]), .B(p_input[2723]), .Z(n16171) );
  AND U24259 ( .A(n16173), .B(n16174), .Z(o[2722]) );
  AND U24260 ( .A(p_input[22722]), .B(p_input[12722]), .Z(n16174) );
  AND U24261 ( .A(p_input[32722]), .B(p_input[2722]), .Z(n16173) );
  AND U24262 ( .A(n16175), .B(n16176), .Z(o[2721]) );
  AND U24263 ( .A(p_input[22721]), .B(p_input[12721]), .Z(n16176) );
  AND U24264 ( .A(p_input[32721]), .B(p_input[2721]), .Z(n16175) );
  AND U24265 ( .A(n16177), .B(n16178), .Z(o[2720]) );
  AND U24266 ( .A(p_input[22720]), .B(p_input[12720]), .Z(n16178) );
  AND U24267 ( .A(p_input[32720]), .B(p_input[2720]), .Z(n16177) );
  AND U24268 ( .A(n16179), .B(n16180), .Z(o[271]) );
  AND U24269 ( .A(p_input[20271]), .B(p_input[10271]), .Z(n16180) );
  AND U24270 ( .A(p_input[30271]), .B(p_input[271]), .Z(n16179) );
  AND U24271 ( .A(n16181), .B(n16182), .Z(o[2719]) );
  AND U24272 ( .A(p_input[22719]), .B(p_input[12719]), .Z(n16182) );
  AND U24273 ( .A(p_input[32719]), .B(p_input[2719]), .Z(n16181) );
  AND U24274 ( .A(n16183), .B(n16184), .Z(o[2718]) );
  AND U24275 ( .A(p_input[22718]), .B(p_input[12718]), .Z(n16184) );
  AND U24276 ( .A(p_input[32718]), .B(p_input[2718]), .Z(n16183) );
  AND U24277 ( .A(n16185), .B(n16186), .Z(o[2717]) );
  AND U24278 ( .A(p_input[22717]), .B(p_input[12717]), .Z(n16186) );
  AND U24279 ( .A(p_input[32717]), .B(p_input[2717]), .Z(n16185) );
  AND U24280 ( .A(n16187), .B(n16188), .Z(o[2716]) );
  AND U24281 ( .A(p_input[22716]), .B(p_input[12716]), .Z(n16188) );
  AND U24282 ( .A(p_input[32716]), .B(p_input[2716]), .Z(n16187) );
  AND U24283 ( .A(n16189), .B(n16190), .Z(o[2715]) );
  AND U24284 ( .A(p_input[22715]), .B(p_input[12715]), .Z(n16190) );
  AND U24285 ( .A(p_input[32715]), .B(p_input[2715]), .Z(n16189) );
  AND U24286 ( .A(n16191), .B(n16192), .Z(o[2714]) );
  AND U24287 ( .A(p_input[22714]), .B(p_input[12714]), .Z(n16192) );
  AND U24288 ( .A(p_input[32714]), .B(p_input[2714]), .Z(n16191) );
  AND U24289 ( .A(n16193), .B(n16194), .Z(o[2713]) );
  AND U24290 ( .A(p_input[22713]), .B(p_input[12713]), .Z(n16194) );
  AND U24291 ( .A(p_input[32713]), .B(p_input[2713]), .Z(n16193) );
  AND U24292 ( .A(n16195), .B(n16196), .Z(o[2712]) );
  AND U24293 ( .A(p_input[22712]), .B(p_input[12712]), .Z(n16196) );
  AND U24294 ( .A(p_input[32712]), .B(p_input[2712]), .Z(n16195) );
  AND U24295 ( .A(n16197), .B(n16198), .Z(o[2711]) );
  AND U24296 ( .A(p_input[22711]), .B(p_input[12711]), .Z(n16198) );
  AND U24297 ( .A(p_input[32711]), .B(p_input[2711]), .Z(n16197) );
  AND U24298 ( .A(n16199), .B(n16200), .Z(o[2710]) );
  AND U24299 ( .A(p_input[22710]), .B(p_input[12710]), .Z(n16200) );
  AND U24300 ( .A(p_input[32710]), .B(p_input[2710]), .Z(n16199) );
  AND U24301 ( .A(n16201), .B(n16202), .Z(o[270]) );
  AND U24302 ( .A(p_input[20270]), .B(p_input[10270]), .Z(n16202) );
  AND U24303 ( .A(p_input[30270]), .B(p_input[270]), .Z(n16201) );
  AND U24304 ( .A(n16203), .B(n16204), .Z(o[2709]) );
  AND U24305 ( .A(p_input[22709]), .B(p_input[12709]), .Z(n16204) );
  AND U24306 ( .A(p_input[32709]), .B(p_input[2709]), .Z(n16203) );
  AND U24307 ( .A(n16205), .B(n16206), .Z(o[2708]) );
  AND U24308 ( .A(p_input[22708]), .B(p_input[12708]), .Z(n16206) );
  AND U24309 ( .A(p_input[32708]), .B(p_input[2708]), .Z(n16205) );
  AND U24310 ( .A(n16207), .B(n16208), .Z(o[2707]) );
  AND U24311 ( .A(p_input[22707]), .B(p_input[12707]), .Z(n16208) );
  AND U24312 ( .A(p_input[32707]), .B(p_input[2707]), .Z(n16207) );
  AND U24313 ( .A(n16209), .B(n16210), .Z(o[2706]) );
  AND U24314 ( .A(p_input[22706]), .B(p_input[12706]), .Z(n16210) );
  AND U24315 ( .A(p_input[32706]), .B(p_input[2706]), .Z(n16209) );
  AND U24316 ( .A(n16211), .B(n16212), .Z(o[2705]) );
  AND U24317 ( .A(p_input[22705]), .B(p_input[12705]), .Z(n16212) );
  AND U24318 ( .A(p_input[32705]), .B(p_input[2705]), .Z(n16211) );
  AND U24319 ( .A(n16213), .B(n16214), .Z(o[2704]) );
  AND U24320 ( .A(p_input[22704]), .B(p_input[12704]), .Z(n16214) );
  AND U24321 ( .A(p_input[32704]), .B(p_input[2704]), .Z(n16213) );
  AND U24322 ( .A(n16215), .B(n16216), .Z(o[2703]) );
  AND U24323 ( .A(p_input[22703]), .B(p_input[12703]), .Z(n16216) );
  AND U24324 ( .A(p_input[32703]), .B(p_input[2703]), .Z(n16215) );
  AND U24325 ( .A(n16217), .B(n16218), .Z(o[2702]) );
  AND U24326 ( .A(p_input[22702]), .B(p_input[12702]), .Z(n16218) );
  AND U24327 ( .A(p_input[32702]), .B(p_input[2702]), .Z(n16217) );
  AND U24328 ( .A(n16219), .B(n16220), .Z(o[2701]) );
  AND U24329 ( .A(p_input[22701]), .B(p_input[12701]), .Z(n16220) );
  AND U24330 ( .A(p_input[32701]), .B(p_input[2701]), .Z(n16219) );
  AND U24331 ( .A(n16221), .B(n16222), .Z(o[2700]) );
  AND U24332 ( .A(p_input[22700]), .B(p_input[12700]), .Z(n16222) );
  AND U24333 ( .A(p_input[32700]), .B(p_input[2700]), .Z(n16221) );
  AND U24334 ( .A(n16223), .B(n16224), .Z(o[26]) );
  AND U24335 ( .A(p_input[20026]), .B(p_input[10026]), .Z(n16224) );
  AND U24336 ( .A(p_input[30026]), .B(p_input[26]), .Z(n16223) );
  AND U24337 ( .A(n16225), .B(n16226), .Z(o[269]) );
  AND U24338 ( .A(p_input[20269]), .B(p_input[10269]), .Z(n16226) );
  AND U24339 ( .A(p_input[30269]), .B(p_input[269]), .Z(n16225) );
  AND U24340 ( .A(n16227), .B(n16228), .Z(o[2699]) );
  AND U24341 ( .A(p_input[22699]), .B(p_input[12699]), .Z(n16228) );
  AND U24342 ( .A(p_input[32699]), .B(p_input[2699]), .Z(n16227) );
  AND U24343 ( .A(n16229), .B(n16230), .Z(o[2698]) );
  AND U24344 ( .A(p_input[22698]), .B(p_input[12698]), .Z(n16230) );
  AND U24345 ( .A(p_input[32698]), .B(p_input[2698]), .Z(n16229) );
  AND U24346 ( .A(n16231), .B(n16232), .Z(o[2697]) );
  AND U24347 ( .A(p_input[22697]), .B(p_input[12697]), .Z(n16232) );
  AND U24348 ( .A(p_input[32697]), .B(p_input[2697]), .Z(n16231) );
  AND U24349 ( .A(n16233), .B(n16234), .Z(o[2696]) );
  AND U24350 ( .A(p_input[22696]), .B(p_input[12696]), .Z(n16234) );
  AND U24351 ( .A(p_input[32696]), .B(p_input[2696]), .Z(n16233) );
  AND U24352 ( .A(n16235), .B(n16236), .Z(o[2695]) );
  AND U24353 ( .A(p_input[22695]), .B(p_input[12695]), .Z(n16236) );
  AND U24354 ( .A(p_input[32695]), .B(p_input[2695]), .Z(n16235) );
  AND U24355 ( .A(n16237), .B(n16238), .Z(o[2694]) );
  AND U24356 ( .A(p_input[22694]), .B(p_input[12694]), .Z(n16238) );
  AND U24357 ( .A(p_input[32694]), .B(p_input[2694]), .Z(n16237) );
  AND U24358 ( .A(n16239), .B(n16240), .Z(o[2693]) );
  AND U24359 ( .A(p_input[22693]), .B(p_input[12693]), .Z(n16240) );
  AND U24360 ( .A(p_input[32693]), .B(p_input[2693]), .Z(n16239) );
  AND U24361 ( .A(n16241), .B(n16242), .Z(o[2692]) );
  AND U24362 ( .A(p_input[22692]), .B(p_input[12692]), .Z(n16242) );
  AND U24363 ( .A(p_input[32692]), .B(p_input[2692]), .Z(n16241) );
  AND U24364 ( .A(n16243), .B(n16244), .Z(o[2691]) );
  AND U24365 ( .A(p_input[22691]), .B(p_input[12691]), .Z(n16244) );
  AND U24366 ( .A(p_input[32691]), .B(p_input[2691]), .Z(n16243) );
  AND U24367 ( .A(n16245), .B(n16246), .Z(o[2690]) );
  AND U24368 ( .A(p_input[22690]), .B(p_input[12690]), .Z(n16246) );
  AND U24369 ( .A(p_input[32690]), .B(p_input[2690]), .Z(n16245) );
  AND U24370 ( .A(n16247), .B(n16248), .Z(o[268]) );
  AND U24371 ( .A(p_input[20268]), .B(p_input[10268]), .Z(n16248) );
  AND U24372 ( .A(p_input[30268]), .B(p_input[268]), .Z(n16247) );
  AND U24373 ( .A(n16249), .B(n16250), .Z(o[2689]) );
  AND U24374 ( .A(p_input[22689]), .B(p_input[12689]), .Z(n16250) );
  AND U24375 ( .A(p_input[32689]), .B(p_input[2689]), .Z(n16249) );
  AND U24376 ( .A(n16251), .B(n16252), .Z(o[2688]) );
  AND U24377 ( .A(p_input[22688]), .B(p_input[12688]), .Z(n16252) );
  AND U24378 ( .A(p_input[32688]), .B(p_input[2688]), .Z(n16251) );
  AND U24379 ( .A(n16253), .B(n16254), .Z(o[2687]) );
  AND U24380 ( .A(p_input[22687]), .B(p_input[12687]), .Z(n16254) );
  AND U24381 ( .A(p_input[32687]), .B(p_input[2687]), .Z(n16253) );
  AND U24382 ( .A(n16255), .B(n16256), .Z(o[2686]) );
  AND U24383 ( .A(p_input[22686]), .B(p_input[12686]), .Z(n16256) );
  AND U24384 ( .A(p_input[32686]), .B(p_input[2686]), .Z(n16255) );
  AND U24385 ( .A(n16257), .B(n16258), .Z(o[2685]) );
  AND U24386 ( .A(p_input[22685]), .B(p_input[12685]), .Z(n16258) );
  AND U24387 ( .A(p_input[32685]), .B(p_input[2685]), .Z(n16257) );
  AND U24388 ( .A(n16259), .B(n16260), .Z(o[2684]) );
  AND U24389 ( .A(p_input[22684]), .B(p_input[12684]), .Z(n16260) );
  AND U24390 ( .A(p_input[32684]), .B(p_input[2684]), .Z(n16259) );
  AND U24391 ( .A(n16261), .B(n16262), .Z(o[2683]) );
  AND U24392 ( .A(p_input[22683]), .B(p_input[12683]), .Z(n16262) );
  AND U24393 ( .A(p_input[32683]), .B(p_input[2683]), .Z(n16261) );
  AND U24394 ( .A(n16263), .B(n16264), .Z(o[2682]) );
  AND U24395 ( .A(p_input[22682]), .B(p_input[12682]), .Z(n16264) );
  AND U24396 ( .A(p_input[32682]), .B(p_input[2682]), .Z(n16263) );
  AND U24397 ( .A(n16265), .B(n16266), .Z(o[2681]) );
  AND U24398 ( .A(p_input[22681]), .B(p_input[12681]), .Z(n16266) );
  AND U24399 ( .A(p_input[32681]), .B(p_input[2681]), .Z(n16265) );
  AND U24400 ( .A(n16267), .B(n16268), .Z(o[2680]) );
  AND U24401 ( .A(p_input[22680]), .B(p_input[12680]), .Z(n16268) );
  AND U24402 ( .A(p_input[32680]), .B(p_input[2680]), .Z(n16267) );
  AND U24403 ( .A(n16269), .B(n16270), .Z(o[267]) );
  AND U24404 ( .A(p_input[20267]), .B(p_input[10267]), .Z(n16270) );
  AND U24405 ( .A(p_input[30267]), .B(p_input[267]), .Z(n16269) );
  AND U24406 ( .A(n16271), .B(n16272), .Z(o[2679]) );
  AND U24407 ( .A(p_input[22679]), .B(p_input[12679]), .Z(n16272) );
  AND U24408 ( .A(p_input[32679]), .B(p_input[2679]), .Z(n16271) );
  AND U24409 ( .A(n16273), .B(n16274), .Z(o[2678]) );
  AND U24410 ( .A(p_input[22678]), .B(p_input[12678]), .Z(n16274) );
  AND U24411 ( .A(p_input[32678]), .B(p_input[2678]), .Z(n16273) );
  AND U24412 ( .A(n16275), .B(n16276), .Z(o[2677]) );
  AND U24413 ( .A(p_input[22677]), .B(p_input[12677]), .Z(n16276) );
  AND U24414 ( .A(p_input[32677]), .B(p_input[2677]), .Z(n16275) );
  AND U24415 ( .A(n16277), .B(n16278), .Z(o[2676]) );
  AND U24416 ( .A(p_input[22676]), .B(p_input[12676]), .Z(n16278) );
  AND U24417 ( .A(p_input[32676]), .B(p_input[2676]), .Z(n16277) );
  AND U24418 ( .A(n16279), .B(n16280), .Z(o[2675]) );
  AND U24419 ( .A(p_input[22675]), .B(p_input[12675]), .Z(n16280) );
  AND U24420 ( .A(p_input[32675]), .B(p_input[2675]), .Z(n16279) );
  AND U24421 ( .A(n16281), .B(n16282), .Z(o[2674]) );
  AND U24422 ( .A(p_input[22674]), .B(p_input[12674]), .Z(n16282) );
  AND U24423 ( .A(p_input[32674]), .B(p_input[2674]), .Z(n16281) );
  AND U24424 ( .A(n16283), .B(n16284), .Z(o[2673]) );
  AND U24425 ( .A(p_input[22673]), .B(p_input[12673]), .Z(n16284) );
  AND U24426 ( .A(p_input[32673]), .B(p_input[2673]), .Z(n16283) );
  AND U24427 ( .A(n16285), .B(n16286), .Z(o[2672]) );
  AND U24428 ( .A(p_input[22672]), .B(p_input[12672]), .Z(n16286) );
  AND U24429 ( .A(p_input[32672]), .B(p_input[2672]), .Z(n16285) );
  AND U24430 ( .A(n16287), .B(n16288), .Z(o[2671]) );
  AND U24431 ( .A(p_input[22671]), .B(p_input[12671]), .Z(n16288) );
  AND U24432 ( .A(p_input[32671]), .B(p_input[2671]), .Z(n16287) );
  AND U24433 ( .A(n16289), .B(n16290), .Z(o[2670]) );
  AND U24434 ( .A(p_input[22670]), .B(p_input[12670]), .Z(n16290) );
  AND U24435 ( .A(p_input[32670]), .B(p_input[2670]), .Z(n16289) );
  AND U24436 ( .A(n16291), .B(n16292), .Z(o[266]) );
  AND U24437 ( .A(p_input[20266]), .B(p_input[10266]), .Z(n16292) );
  AND U24438 ( .A(p_input[30266]), .B(p_input[266]), .Z(n16291) );
  AND U24439 ( .A(n16293), .B(n16294), .Z(o[2669]) );
  AND U24440 ( .A(p_input[22669]), .B(p_input[12669]), .Z(n16294) );
  AND U24441 ( .A(p_input[32669]), .B(p_input[2669]), .Z(n16293) );
  AND U24442 ( .A(n16295), .B(n16296), .Z(o[2668]) );
  AND U24443 ( .A(p_input[22668]), .B(p_input[12668]), .Z(n16296) );
  AND U24444 ( .A(p_input[32668]), .B(p_input[2668]), .Z(n16295) );
  AND U24445 ( .A(n16297), .B(n16298), .Z(o[2667]) );
  AND U24446 ( .A(p_input[22667]), .B(p_input[12667]), .Z(n16298) );
  AND U24447 ( .A(p_input[32667]), .B(p_input[2667]), .Z(n16297) );
  AND U24448 ( .A(n16299), .B(n16300), .Z(o[2666]) );
  AND U24449 ( .A(p_input[22666]), .B(p_input[12666]), .Z(n16300) );
  AND U24450 ( .A(p_input[32666]), .B(p_input[2666]), .Z(n16299) );
  AND U24451 ( .A(n16301), .B(n16302), .Z(o[2665]) );
  AND U24452 ( .A(p_input[22665]), .B(p_input[12665]), .Z(n16302) );
  AND U24453 ( .A(p_input[32665]), .B(p_input[2665]), .Z(n16301) );
  AND U24454 ( .A(n16303), .B(n16304), .Z(o[2664]) );
  AND U24455 ( .A(p_input[22664]), .B(p_input[12664]), .Z(n16304) );
  AND U24456 ( .A(p_input[32664]), .B(p_input[2664]), .Z(n16303) );
  AND U24457 ( .A(n16305), .B(n16306), .Z(o[2663]) );
  AND U24458 ( .A(p_input[22663]), .B(p_input[12663]), .Z(n16306) );
  AND U24459 ( .A(p_input[32663]), .B(p_input[2663]), .Z(n16305) );
  AND U24460 ( .A(n16307), .B(n16308), .Z(o[2662]) );
  AND U24461 ( .A(p_input[22662]), .B(p_input[12662]), .Z(n16308) );
  AND U24462 ( .A(p_input[32662]), .B(p_input[2662]), .Z(n16307) );
  AND U24463 ( .A(n16309), .B(n16310), .Z(o[2661]) );
  AND U24464 ( .A(p_input[22661]), .B(p_input[12661]), .Z(n16310) );
  AND U24465 ( .A(p_input[32661]), .B(p_input[2661]), .Z(n16309) );
  AND U24466 ( .A(n16311), .B(n16312), .Z(o[2660]) );
  AND U24467 ( .A(p_input[22660]), .B(p_input[12660]), .Z(n16312) );
  AND U24468 ( .A(p_input[32660]), .B(p_input[2660]), .Z(n16311) );
  AND U24469 ( .A(n16313), .B(n16314), .Z(o[265]) );
  AND U24470 ( .A(p_input[20265]), .B(p_input[10265]), .Z(n16314) );
  AND U24471 ( .A(p_input[30265]), .B(p_input[265]), .Z(n16313) );
  AND U24472 ( .A(n16315), .B(n16316), .Z(o[2659]) );
  AND U24473 ( .A(p_input[22659]), .B(p_input[12659]), .Z(n16316) );
  AND U24474 ( .A(p_input[32659]), .B(p_input[2659]), .Z(n16315) );
  AND U24475 ( .A(n16317), .B(n16318), .Z(o[2658]) );
  AND U24476 ( .A(p_input[22658]), .B(p_input[12658]), .Z(n16318) );
  AND U24477 ( .A(p_input[32658]), .B(p_input[2658]), .Z(n16317) );
  AND U24478 ( .A(n16319), .B(n16320), .Z(o[2657]) );
  AND U24479 ( .A(p_input[22657]), .B(p_input[12657]), .Z(n16320) );
  AND U24480 ( .A(p_input[32657]), .B(p_input[2657]), .Z(n16319) );
  AND U24481 ( .A(n16321), .B(n16322), .Z(o[2656]) );
  AND U24482 ( .A(p_input[22656]), .B(p_input[12656]), .Z(n16322) );
  AND U24483 ( .A(p_input[32656]), .B(p_input[2656]), .Z(n16321) );
  AND U24484 ( .A(n16323), .B(n16324), .Z(o[2655]) );
  AND U24485 ( .A(p_input[22655]), .B(p_input[12655]), .Z(n16324) );
  AND U24486 ( .A(p_input[32655]), .B(p_input[2655]), .Z(n16323) );
  AND U24487 ( .A(n16325), .B(n16326), .Z(o[2654]) );
  AND U24488 ( .A(p_input[22654]), .B(p_input[12654]), .Z(n16326) );
  AND U24489 ( .A(p_input[32654]), .B(p_input[2654]), .Z(n16325) );
  AND U24490 ( .A(n16327), .B(n16328), .Z(o[2653]) );
  AND U24491 ( .A(p_input[22653]), .B(p_input[12653]), .Z(n16328) );
  AND U24492 ( .A(p_input[32653]), .B(p_input[2653]), .Z(n16327) );
  AND U24493 ( .A(n16329), .B(n16330), .Z(o[2652]) );
  AND U24494 ( .A(p_input[22652]), .B(p_input[12652]), .Z(n16330) );
  AND U24495 ( .A(p_input[32652]), .B(p_input[2652]), .Z(n16329) );
  AND U24496 ( .A(n16331), .B(n16332), .Z(o[2651]) );
  AND U24497 ( .A(p_input[22651]), .B(p_input[12651]), .Z(n16332) );
  AND U24498 ( .A(p_input[32651]), .B(p_input[2651]), .Z(n16331) );
  AND U24499 ( .A(n16333), .B(n16334), .Z(o[2650]) );
  AND U24500 ( .A(p_input[22650]), .B(p_input[12650]), .Z(n16334) );
  AND U24501 ( .A(p_input[32650]), .B(p_input[2650]), .Z(n16333) );
  AND U24502 ( .A(n16335), .B(n16336), .Z(o[264]) );
  AND U24503 ( .A(p_input[20264]), .B(p_input[10264]), .Z(n16336) );
  AND U24504 ( .A(p_input[30264]), .B(p_input[264]), .Z(n16335) );
  AND U24505 ( .A(n16337), .B(n16338), .Z(o[2649]) );
  AND U24506 ( .A(p_input[22649]), .B(p_input[12649]), .Z(n16338) );
  AND U24507 ( .A(p_input[32649]), .B(p_input[2649]), .Z(n16337) );
  AND U24508 ( .A(n16339), .B(n16340), .Z(o[2648]) );
  AND U24509 ( .A(p_input[22648]), .B(p_input[12648]), .Z(n16340) );
  AND U24510 ( .A(p_input[32648]), .B(p_input[2648]), .Z(n16339) );
  AND U24511 ( .A(n16341), .B(n16342), .Z(o[2647]) );
  AND U24512 ( .A(p_input[22647]), .B(p_input[12647]), .Z(n16342) );
  AND U24513 ( .A(p_input[32647]), .B(p_input[2647]), .Z(n16341) );
  AND U24514 ( .A(n16343), .B(n16344), .Z(o[2646]) );
  AND U24515 ( .A(p_input[22646]), .B(p_input[12646]), .Z(n16344) );
  AND U24516 ( .A(p_input[32646]), .B(p_input[2646]), .Z(n16343) );
  AND U24517 ( .A(n16345), .B(n16346), .Z(o[2645]) );
  AND U24518 ( .A(p_input[22645]), .B(p_input[12645]), .Z(n16346) );
  AND U24519 ( .A(p_input[32645]), .B(p_input[2645]), .Z(n16345) );
  AND U24520 ( .A(n16347), .B(n16348), .Z(o[2644]) );
  AND U24521 ( .A(p_input[22644]), .B(p_input[12644]), .Z(n16348) );
  AND U24522 ( .A(p_input[32644]), .B(p_input[2644]), .Z(n16347) );
  AND U24523 ( .A(n16349), .B(n16350), .Z(o[2643]) );
  AND U24524 ( .A(p_input[22643]), .B(p_input[12643]), .Z(n16350) );
  AND U24525 ( .A(p_input[32643]), .B(p_input[2643]), .Z(n16349) );
  AND U24526 ( .A(n16351), .B(n16352), .Z(o[2642]) );
  AND U24527 ( .A(p_input[22642]), .B(p_input[12642]), .Z(n16352) );
  AND U24528 ( .A(p_input[32642]), .B(p_input[2642]), .Z(n16351) );
  AND U24529 ( .A(n16353), .B(n16354), .Z(o[2641]) );
  AND U24530 ( .A(p_input[22641]), .B(p_input[12641]), .Z(n16354) );
  AND U24531 ( .A(p_input[32641]), .B(p_input[2641]), .Z(n16353) );
  AND U24532 ( .A(n16355), .B(n16356), .Z(o[2640]) );
  AND U24533 ( .A(p_input[22640]), .B(p_input[12640]), .Z(n16356) );
  AND U24534 ( .A(p_input[32640]), .B(p_input[2640]), .Z(n16355) );
  AND U24535 ( .A(n16357), .B(n16358), .Z(o[263]) );
  AND U24536 ( .A(p_input[20263]), .B(p_input[10263]), .Z(n16358) );
  AND U24537 ( .A(p_input[30263]), .B(p_input[263]), .Z(n16357) );
  AND U24538 ( .A(n16359), .B(n16360), .Z(o[2639]) );
  AND U24539 ( .A(p_input[22639]), .B(p_input[12639]), .Z(n16360) );
  AND U24540 ( .A(p_input[32639]), .B(p_input[2639]), .Z(n16359) );
  AND U24541 ( .A(n16361), .B(n16362), .Z(o[2638]) );
  AND U24542 ( .A(p_input[22638]), .B(p_input[12638]), .Z(n16362) );
  AND U24543 ( .A(p_input[32638]), .B(p_input[2638]), .Z(n16361) );
  AND U24544 ( .A(n16363), .B(n16364), .Z(o[2637]) );
  AND U24545 ( .A(p_input[22637]), .B(p_input[12637]), .Z(n16364) );
  AND U24546 ( .A(p_input[32637]), .B(p_input[2637]), .Z(n16363) );
  AND U24547 ( .A(n16365), .B(n16366), .Z(o[2636]) );
  AND U24548 ( .A(p_input[22636]), .B(p_input[12636]), .Z(n16366) );
  AND U24549 ( .A(p_input[32636]), .B(p_input[2636]), .Z(n16365) );
  AND U24550 ( .A(n16367), .B(n16368), .Z(o[2635]) );
  AND U24551 ( .A(p_input[22635]), .B(p_input[12635]), .Z(n16368) );
  AND U24552 ( .A(p_input[32635]), .B(p_input[2635]), .Z(n16367) );
  AND U24553 ( .A(n16369), .B(n16370), .Z(o[2634]) );
  AND U24554 ( .A(p_input[22634]), .B(p_input[12634]), .Z(n16370) );
  AND U24555 ( .A(p_input[32634]), .B(p_input[2634]), .Z(n16369) );
  AND U24556 ( .A(n16371), .B(n16372), .Z(o[2633]) );
  AND U24557 ( .A(p_input[22633]), .B(p_input[12633]), .Z(n16372) );
  AND U24558 ( .A(p_input[32633]), .B(p_input[2633]), .Z(n16371) );
  AND U24559 ( .A(n16373), .B(n16374), .Z(o[2632]) );
  AND U24560 ( .A(p_input[22632]), .B(p_input[12632]), .Z(n16374) );
  AND U24561 ( .A(p_input[32632]), .B(p_input[2632]), .Z(n16373) );
  AND U24562 ( .A(n16375), .B(n16376), .Z(o[2631]) );
  AND U24563 ( .A(p_input[22631]), .B(p_input[12631]), .Z(n16376) );
  AND U24564 ( .A(p_input[32631]), .B(p_input[2631]), .Z(n16375) );
  AND U24565 ( .A(n16377), .B(n16378), .Z(o[2630]) );
  AND U24566 ( .A(p_input[22630]), .B(p_input[12630]), .Z(n16378) );
  AND U24567 ( .A(p_input[32630]), .B(p_input[2630]), .Z(n16377) );
  AND U24568 ( .A(n16379), .B(n16380), .Z(o[262]) );
  AND U24569 ( .A(p_input[20262]), .B(p_input[10262]), .Z(n16380) );
  AND U24570 ( .A(p_input[30262]), .B(p_input[262]), .Z(n16379) );
  AND U24571 ( .A(n16381), .B(n16382), .Z(o[2629]) );
  AND U24572 ( .A(p_input[22629]), .B(p_input[12629]), .Z(n16382) );
  AND U24573 ( .A(p_input[32629]), .B(p_input[2629]), .Z(n16381) );
  AND U24574 ( .A(n16383), .B(n16384), .Z(o[2628]) );
  AND U24575 ( .A(p_input[22628]), .B(p_input[12628]), .Z(n16384) );
  AND U24576 ( .A(p_input[32628]), .B(p_input[2628]), .Z(n16383) );
  AND U24577 ( .A(n16385), .B(n16386), .Z(o[2627]) );
  AND U24578 ( .A(p_input[22627]), .B(p_input[12627]), .Z(n16386) );
  AND U24579 ( .A(p_input[32627]), .B(p_input[2627]), .Z(n16385) );
  AND U24580 ( .A(n16387), .B(n16388), .Z(o[2626]) );
  AND U24581 ( .A(p_input[22626]), .B(p_input[12626]), .Z(n16388) );
  AND U24582 ( .A(p_input[32626]), .B(p_input[2626]), .Z(n16387) );
  AND U24583 ( .A(n16389), .B(n16390), .Z(o[2625]) );
  AND U24584 ( .A(p_input[22625]), .B(p_input[12625]), .Z(n16390) );
  AND U24585 ( .A(p_input[32625]), .B(p_input[2625]), .Z(n16389) );
  AND U24586 ( .A(n16391), .B(n16392), .Z(o[2624]) );
  AND U24587 ( .A(p_input[22624]), .B(p_input[12624]), .Z(n16392) );
  AND U24588 ( .A(p_input[32624]), .B(p_input[2624]), .Z(n16391) );
  AND U24589 ( .A(n16393), .B(n16394), .Z(o[2623]) );
  AND U24590 ( .A(p_input[22623]), .B(p_input[12623]), .Z(n16394) );
  AND U24591 ( .A(p_input[32623]), .B(p_input[2623]), .Z(n16393) );
  AND U24592 ( .A(n16395), .B(n16396), .Z(o[2622]) );
  AND U24593 ( .A(p_input[22622]), .B(p_input[12622]), .Z(n16396) );
  AND U24594 ( .A(p_input[32622]), .B(p_input[2622]), .Z(n16395) );
  AND U24595 ( .A(n16397), .B(n16398), .Z(o[2621]) );
  AND U24596 ( .A(p_input[22621]), .B(p_input[12621]), .Z(n16398) );
  AND U24597 ( .A(p_input[32621]), .B(p_input[2621]), .Z(n16397) );
  AND U24598 ( .A(n16399), .B(n16400), .Z(o[2620]) );
  AND U24599 ( .A(p_input[22620]), .B(p_input[12620]), .Z(n16400) );
  AND U24600 ( .A(p_input[32620]), .B(p_input[2620]), .Z(n16399) );
  AND U24601 ( .A(n16401), .B(n16402), .Z(o[261]) );
  AND U24602 ( .A(p_input[20261]), .B(p_input[10261]), .Z(n16402) );
  AND U24603 ( .A(p_input[30261]), .B(p_input[261]), .Z(n16401) );
  AND U24604 ( .A(n16403), .B(n16404), .Z(o[2619]) );
  AND U24605 ( .A(p_input[22619]), .B(p_input[12619]), .Z(n16404) );
  AND U24606 ( .A(p_input[32619]), .B(p_input[2619]), .Z(n16403) );
  AND U24607 ( .A(n16405), .B(n16406), .Z(o[2618]) );
  AND U24608 ( .A(p_input[22618]), .B(p_input[12618]), .Z(n16406) );
  AND U24609 ( .A(p_input[32618]), .B(p_input[2618]), .Z(n16405) );
  AND U24610 ( .A(n16407), .B(n16408), .Z(o[2617]) );
  AND U24611 ( .A(p_input[22617]), .B(p_input[12617]), .Z(n16408) );
  AND U24612 ( .A(p_input[32617]), .B(p_input[2617]), .Z(n16407) );
  AND U24613 ( .A(n16409), .B(n16410), .Z(o[2616]) );
  AND U24614 ( .A(p_input[22616]), .B(p_input[12616]), .Z(n16410) );
  AND U24615 ( .A(p_input[32616]), .B(p_input[2616]), .Z(n16409) );
  AND U24616 ( .A(n16411), .B(n16412), .Z(o[2615]) );
  AND U24617 ( .A(p_input[22615]), .B(p_input[12615]), .Z(n16412) );
  AND U24618 ( .A(p_input[32615]), .B(p_input[2615]), .Z(n16411) );
  AND U24619 ( .A(n16413), .B(n16414), .Z(o[2614]) );
  AND U24620 ( .A(p_input[22614]), .B(p_input[12614]), .Z(n16414) );
  AND U24621 ( .A(p_input[32614]), .B(p_input[2614]), .Z(n16413) );
  AND U24622 ( .A(n16415), .B(n16416), .Z(o[2613]) );
  AND U24623 ( .A(p_input[22613]), .B(p_input[12613]), .Z(n16416) );
  AND U24624 ( .A(p_input[32613]), .B(p_input[2613]), .Z(n16415) );
  AND U24625 ( .A(n16417), .B(n16418), .Z(o[2612]) );
  AND U24626 ( .A(p_input[22612]), .B(p_input[12612]), .Z(n16418) );
  AND U24627 ( .A(p_input[32612]), .B(p_input[2612]), .Z(n16417) );
  AND U24628 ( .A(n16419), .B(n16420), .Z(o[2611]) );
  AND U24629 ( .A(p_input[22611]), .B(p_input[12611]), .Z(n16420) );
  AND U24630 ( .A(p_input[32611]), .B(p_input[2611]), .Z(n16419) );
  AND U24631 ( .A(n16421), .B(n16422), .Z(o[2610]) );
  AND U24632 ( .A(p_input[22610]), .B(p_input[12610]), .Z(n16422) );
  AND U24633 ( .A(p_input[32610]), .B(p_input[2610]), .Z(n16421) );
  AND U24634 ( .A(n16423), .B(n16424), .Z(o[260]) );
  AND U24635 ( .A(p_input[20260]), .B(p_input[10260]), .Z(n16424) );
  AND U24636 ( .A(p_input[30260]), .B(p_input[260]), .Z(n16423) );
  AND U24637 ( .A(n16425), .B(n16426), .Z(o[2609]) );
  AND U24638 ( .A(p_input[22609]), .B(p_input[12609]), .Z(n16426) );
  AND U24639 ( .A(p_input[32609]), .B(p_input[2609]), .Z(n16425) );
  AND U24640 ( .A(n16427), .B(n16428), .Z(o[2608]) );
  AND U24641 ( .A(p_input[22608]), .B(p_input[12608]), .Z(n16428) );
  AND U24642 ( .A(p_input[32608]), .B(p_input[2608]), .Z(n16427) );
  AND U24643 ( .A(n16429), .B(n16430), .Z(o[2607]) );
  AND U24644 ( .A(p_input[22607]), .B(p_input[12607]), .Z(n16430) );
  AND U24645 ( .A(p_input[32607]), .B(p_input[2607]), .Z(n16429) );
  AND U24646 ( .A(n16431), .B(n16432), .Z(o[2606]) );
  AND U24647 ( .A(p_input[22606]), .B(p_input[12606]), .Z(n16432) );
  AND U24648 ( .A(p_input[32606]), .B(p_input[2606]), .Z(n16431) );
  AND U24649 ( .A(n16433), .B(n16434), .Z(o[2605]) );
  AND U24650 ( .A(p_input[22605]), .B(p_input[12605]), .Z(n16434) );
  AND U24651 ( .A(p_input[32605]), .B(p_input[2605]), .Z(n16433) );
  AND U24652 ( .A(n16435), .B(n16436), .Z(o[2604]) );
  AND U24653 ( .A(p_input[22604]), .B(p_input[12604]), .Z(n16436) );
  AND U24654 ( .A(p_input[32604]), .B(p_input[2604]), .Z(n16435) );
  AND U24655 ( .A(n16437), .B(n16438), .Z(o[2603]) );
  AND U24656 ( .A(p_input[22603]), .B(p_input[12603]), .Z(n16438) );
  AND U24657 ( .A(p_input[32603]), .B(p_input[2603]), .Z(n16437) );
  AND U24658 ( .A(n16439), .B(n16440), .Z(o[2602]) );
  AND U24659 ( .A(p_input[22602]), .B(p_input[12602]), .Z(n16440) );
  AND U24660 ( .A(p_input[32602]), .B(p_input[2602]), .Z(n16439) );
  AND U24661 ( .A(n16441), .B(n16442), .Z(o[2601]) );
  AND U24662 ( .A(p_input[22601]), .B(p_input[12601]), .Z(n16442) );
  AND U24663 ( .A(p_input[32601]), .B(p_input[2601]), .Z(n16441) );
  AND U24664 ( .A(n16443), .B(n16444), .Z(o[2600]) );
  AND U24665 ( .A(p_input[22600]), .B(p_input[12600]), .Z(n16444) );
  AND U24666 ( .A(p_input[32600]), .B(p_input[2600]), .Z(n16443) );
  AND U24667 ( .A(n16445), .B(n16446), .Z(o[25]) );
  AND U24668 ( .A(p_input[20025]), .B(p_input[10025]), .Z(n16446) );
  AND U24669 ( .A(p_input[30025]), .B(p_input[25]), .Z(n16445) );
  AND U24670 ( .A(n16447), .B(n16448), .Z(o[259]) );
  AND U24671 ( .A(p_input[20259]), .B(p_input[10259]), .Z(n16448) );
  AND U24672 ( .A(p_input[30259]), .B(p_input[259]), .Z(n16447) );
  AND U24673 ( .A(n16449), .B(n16450), .Z(o[2599]) );
  AND U24674 ( .A(p_input[22599]), .B(p_input[12599]), .Z(n16450) );
  AND U24675 ( .A(p_input[32599]), .B(p_input[2599]), .Z(n16449) );
  AND U24676 ( .A(n16451), .B(n16452), .Z(o[2598]) );
  AND U24677 ( .A(p_input[22598]), .B(p_input[12598]), .Z(n16452) );
  AND U24678 ( .A(p_input[32598]), .B(p_input[2598]), .Z(n16451) );
  AND U24679 ( .A(n16453), .B(n16454), .Z(o[2597]) );
  AND U24680 ( .A(p_input[22597]), .B(p_input[12597]), .Z(n16454) );
  AND U24681 ( .A(p_input[32597]), .B(p_input[2597]), .Z(n16453) );
  AND U24682 ( .A(n16455), .B(n16456), .Z(o[2596]) );
  AND U24683 ( .A(p_input[22596]), .B(p_input[12596]), .Z(n16456) );
  AND U24684 ( .A(p_input[32596]), .B(p_input[2596]), .Z(n16455) );
  AND U24685 ( .A(n16457), .B(n16458), .Z(o[2595]) );
  AND U24686 ( .A(p_input[22595]), .B(p_input[12595]), .Z(n16458) );
  AND U24687 ( .A(p_input[32595]), .B(p_input[2595]), .Z(n16457) );
  AND U24688 ( .A(n16459), .B(n16460), .Z(o[2594]) );
  AND U24689 ( .A(p_input[22594]), .B(p_input[12594]), .Z(n16460) );
  AND U24690 ( .A(p_input[32594]), .B(p_input[2594]), .Z(n16459) );
  AND U24691 ( .A(n16461), .B(n16462), .Z(o[2593]) );
  AND U24692 ( .A(p_input[22593]), .B(p_input[12593]), .Z(n16462) );
  AND U24693 ( .A(p_input[32593]), .B(p_input[2593]), .Z(n16461) );
  AND U24694 ( .A(n16463), .B(n16464), .Z(o[2592]) );
  AND U24695 ( .A(p_input[22592]), .B(p_input[12592]), .Z(n16464) );
  AND U24696 ( .A(p_input[32592]), .B(p_input[2592]), .Z(n16463) );
  AND U24697 ( .A(n16465), .B(n16466), .Z(o[2591]) );
  AND U24698 ( .A(p_input[22591]), .B(p_input[12591]), .Z(n16466) );
  AND U24699 ( .A(p_input[32591]), .B(p_input[2591]), .Z(n16465) );
  AND U24700 ( .A(n16467), .B(n16468), .Z(o[2590]) );
  AND U24701 ( .A(p_input[22590]), .B(p_input[12590]), .Z(n16468) );
  AND U24702 ( .A(p_input[32590]), .B(p_input[2590]), .Z(n16467) );
  AND U24703 ( .A(n16469), .B(n16470), .Z(o[258]) );
  AND U24704 ( .A(p_input[20258]), .B(p_input[10258]), .Z(n16470) );
  AND U24705 ( .A(p_input[30258]), .B(p_input[258]), .Z(n16469) );
  AND U24706 ( .A(n16471), .B(n16472), .Z(o[2589]) );
  AND U24707 ( .A(p_input[22589]), .B(p_input[12589]), .Z(n16472) );
  AND U24708 ( .A(p_input[32589]), .B(p_input[2589]), .Z(n16471) );
  AND U24709 ( .A(n16473), .B(n16474), .Z(o[2588]) );
  AND U24710 ( .A(p_input[22588]), .B(p_input[12588]), .Z(n16474) );
  AND U24711 ( .A(p_input[32588]), .B(p_input[2588]), .Z(n16473) );
  AND U24712 ( .A(n16475), .B(n16476), .Z(o[2587]) );
  AND U24713 ( .A(p_input[22587]), .B(p_input[12587]), .Z(n16476) );
  AND U24714 ( .A(p_input[32587]), .B(p_input[2587]), .Z(n16475) );
  AND U24715 ( .A(n16477), .B(n16478), .Z(o[2586]) );
  AND U24716 ( .A(p_input[22586]), .B(p_input[12586]), .Z(n16478) );
  AND U24717 ( .A(p_input[32586]), .B(p_input[2586]), .Z(n16477) );
  AND U24718 ( .A(n16479), .B(n16480), .Z(o[2585]) );
  AND U24719 ( .A(p_input[22585]), .B(p_input[12585]), .Z(n16480) );
  AND U24720 ( .A(p_input[32585]), .B(p_input[2585]), .Z(n16479) );
  AND U24721 ( .A(n16481), .B(n16482), .Z(o[2584]) );
  AND U24722 ( .A(p_input[22584]), .B(p_input[12584]), .Z(n16482) );
  AND U24723 ( .A(p_input[32584]), .B(p_input[2584]), .Z(n16481) );
  AND U24724 ( .A(n16483), .B(n16484), .Z(o[2583]) );
  AND U24725 ( .A(p_input[22583]), .B(p_input[12583]), .Z(n16484) );
  AND U24726 ( .A(p_input[32583]), .B(p_input[2583]), .Z(n16483) );
  AND U24727 ( .A(n16485), .B(n16486), .Z(o[2582]) );
  AND U24728 ( .A(p_input[22582]), .B(p_input[12582]), .Z(n16486) );
  AND U24729 ( .A(p_input[32582]), .B(p_input[2582]), .Z(n16485) );
  AND U24730 ( .A(n16487), .B(n16488), .Z(o[2581]) );
  AND U24731 ( .A(p_input[22581]), .B(p_input[12581]), .Z(n16488) );
  AND U24732 ( .A(p_input[32581]), .B(p_input[2581]), .Z(n16487) );
  AND U24733 ( .A(n16489), .B(n16490), .Z(o[2580]) );
  AND U24734 ( .A(p_input[22580]), .B(p_input[12580]), .Z(n16490) );
  AND U24735 ( .A(p_input[32580]), .B(p_input[2580]), .Z(n16489) );
  AND U24736 ( .A(n16491), .B(n16492), .Z(o[257]) );
  AND U24737 ( .A(p_input[20257]), .B(p_input[10257]), .Z(n16492) );
  AND U24738 ( .A(p_input[30257]), .B(p_input[257]), .Z(n16491) );
  AND U24739 ( .A(n16493), .B(n16494), .Z(o[2579]) );
  AND U24740 ( .A(p_input[22579]), .B(p_input[12579]), .Z(n16494) );
  AND U24741 ( .A(p_input[32579]), .B(p_input[2579]), .Z(n16493) );
  AND U24742 ( .A(n16495), .B(n16496), .Z(o[2578]) );
  AND U24743 ( .A(p_input[22578]), .B(p_input[12578]), .Z(n16496) );
  AND U24744 ( .A(p_input[32578]), .B(p_input[2578]), .Z(n16495) );
  AND U24745 ( .A(n16497), .B(n16498), .Z(o[2577]) );
  AND U24746 ( .A(p_input[22577]), .B(p_input[12577]), .Z(n16498) );
  AND U24747 ( .A(p_input[32577]), .B(p_input[2577]), .Z(n16497) );
  AND U24748 ( .A(n16499), .B(n16500), .Z(o[2576]) );
  AND U24749 ( .A(p_input[22576]), .B(p_input[12576]), .Z(n16500) );
  AND U24750 ( .A(p_input[32576]), .B(p_input[2576]), .Z(n16499) );
  AND U24751 ( .A(n16501), .B(n16502), .Z(o[2575]) );
  AND U24752 ( .A(p_input[22575]), .B(p_input[12575]), .Z(n16502) );
  AND U24753 ( .A(p_input[32575]), .B(p_input[2575]), .Z(n16501) );
  AND U24754 ( .A(n16503), .B(n16504), .Z(o[2574]) );
  AND U24755 ( .A(p_input[22574]), .B(p_input[12574]), .Z(n16504) );
  AND U24756 ( .A(p_input[32574]), .B(p_input[2574]), .Z(n16503) );
  AND U24757 ( .A(n16505), .B(n16506), .Z(o[2573]) );
  AND U24758 ( .A(p_input[22573]), .B(p_input[12573]), .Z(n16506) );
  AND U24759 ( .A(p_input[32573]), .B(p_input[2573]), .Z(n16505) );
  AND U24760 ( .A(n16507), .B(n16508), .Z(o[2572]) );
  AND U24761 ( .A(p_input[22572]), .B(p_input[12572]), .Z(n16508) );
  AND U24762 ( .A(p_input[32572]), .B(p_input[2572]), .Z(n16507) );
  AND U24763 ( .A(n16509), .B(n16510), .Z(o[2571]) );
  AND U24764 ( .A(p_input[22571]), .B(p_input[12571]), .Z(n16510) );
  AND U24765 ( .A(p_input[32571]), .B(p_input[2571]), .Z(n16509) );
  AND U24766 ( .A(n16511), .B(n16512), .Z(o[2570]) );
  AND U24767 ( .A(p_input[22570]), .B(p_input[12570]), .Z(n16512) );
  AND U24768 ( .A(p_input[32570]), .B(p_input[2570]), .Z(n16511) );
  AND U24769 ( .A(n16513), .B(n16514), .Z(o[256]) );
  AND U24770 ( .A(p_input[20256]), .B(p_input[10256]), .Z(n16514) );
  AND U24771 ( .A(p_input[30256]), .B(p_input[256]), .Z(n16513) );
  AND U24772 ( .A(n16515), .B(n16516), .Z(o[2569]) );
  AND U24773 ( .A(p_input[22569]), .B(p_input[12569]), .Z(n16516) );
  AND U24774 ( .A(p_input[32569]), .B(p_input[2569]), .Z(n16515) );
  AND U24775 ( .A(n16517), .B(n16518), .Z(o[2568]) );
  AND U24776 ( .A(p_input[22568]), .B(p_input[12568]), .Z(n16518) );
  AND U24777 ( .A(p_input[32568]), .B(p_input[2568]), .Z(n16517) );
  AND U24778 ( .A(n16519), .B(n16520), .Z(o[2567]) );
  AND U24779 ( .A(p_input[22567]), .B(p_input[12567]), .Z(n16520) );
  AND U24780 ( .A(p_input[32567]), .B(p_input[2567]), .Z(n16519) );
  AND U24781 ( .A(n16521), .B(n16522), .Z(o[2566]) );
  AND U24782 ( .A(p_input[22566]), .B(p_input[12566]), .Z(n16522) );
  AND U24783 ( .A(p_input[32566]), .B(p_input[2566]), .Z(n16521) );
  AND U24784 ( .A(n16523), .B(n16524), .Z(o[2565]) );
  AND U24785 ( .A(p_input[22565]), .B(p_input[12565]), .Z(n16524) );
  AND U24786 ( .A(p_input[32565]), .B(p_input[2565]), .Z(n16523) );
  AND U24787 ( .A(n16525), .B(n16526), .Z(o[2564]) );
  AND U24788 ( .A(p_input[22564]), .B(p_input[12564]), .Z(n16526) );
  AND U24789 ( .A(p_input[32564]), .B(p_input[2564]), .Z(n16525) );
  AND U24790 ( .A(n16527), .B(n16528), .Z(o[2563]) );
  AND U24791 ( .A(p_input[22563]), .B(p_input[12563]), .Z(n16528) );
  AND U24792 ( .A(p_input[32563]), .B(p_input[2563]), .Z(n16527) );
  AND U24793 ( .A(n16529), .B(n16530), .Z(o[2562]) );
  AND U24794 ( .A(p_input[22562]), .B(p_input[12562]), .Z(n16530) );
  AND U24795 ( .A(p_input[32562]), .B(p_input[2562]), .Z(n16529) );
  AND U24796 ( .A(n16531), .B(n16532), .Z(o[2561]) );
  AND U24797 ( .A(p_input[22561]), .B(p_input[12561]), .Z(n16532) );
  AND U24798 ( .A(p_input[32561]), .B(p_input[2561]), .Z(n16531) );
  AND U24799 ( .A(n16533), .B(n16534), .Z(o[2560]) );
  AND U24800 ( .A(p_input[22560]), .B(p_input[12560]), .Z(n16534) );
  AND U24801 ( .A(p_input[32560]), .B(p_input[2560]), .Z(n16533) );
  AND U24802 ( .A(n16535), .B(n16536), .Z(o[255]) );
  AND U24803 ( .A(p_input[20255]), .B(p_input[10255]), .Z(n16536) );
  AND U24804 ( .A(p_input[30255]), .B(p_input[255]), .Z(n16535) );
  AND U24805 ( .A(n16537), .B(n16538), .Z(o[2559]) );
  AND U24806 ( .A(p_input[22559]), .B(p_input[12559]), .Z(n16538) );
  AND U24807 ( .A(p_input[32559]), .B(p_input[2559]), .Z(n16537) );
  AND U24808 ( .A(n16539), .B(n16540), .Z(o[2558]) );
  AND U24809 ( .A(p_input[22558]), .B(p_input[12558]), .Z(n16540) );
  AND U24810 ( .A(p_input[32558]), .B(p_input[2558]), .Z(n16539) );
  AND U24811 ( .A(n16541), .B(n16542), .Z(o[2557]) );
  AND U24812 ( .A(p_input[22557]), .B(p_input[12557]), .Z(n16542) );
  AND U24813 ( .A(p_input[32557]), .B(p_input[2557]), .Z(n16541) );
  AND U24814 ( .A(n16543), .B(n16544), .Z(o[2556]) );
  AND U24815 ( .A(p_input[22556]), .B(p_input[12556]), .Z(n16544) );
  AND U24816 ( .A(p_input[32556]), .B(p_input[2556]), .Z(n16543) );
  AND U24817 ( .A(n16545), .B(n16546), .Z(o[2555]) );
  AND U24818 ( .A(p_input[22555]), .B(p_input[12555]), .Z(n16546) );
  AND U24819 ( .A(p_input[32555]), .B(p_input[2555]), .Z(n16545) );
  AND U24820 ( .A(n16547), .B(n16548), .Z(o[2554]) );
  AND U24821 ( .A(p_input[22554]), .B(p_input[12554]), .Z(n16548) );
  AND U24822 ( .A(p_input[32554]), .B(p_input[2554]), .Z(n16547) );
  AND U24823 ( .A(n16549), .B(n16550), .Z(o[2553]) );
  AND U24824 ( .A(p_input[22553]), .B(p_input[12553]), .Z(n16550) );
  AND U24825 ( .A(p_input[32553]), .B(p_input[2553]), .Z(n16549) );
  AND U24826 ( .A(n16551), .B(n16552), .Z(o[2552]) );
  AND U24827 ( .A(p_input[22552]), .B(p_input[12552]), .Z(n16552) );
  AND U24828 ( .A(p_input[32552]), .B(p_input[2552]), .Z(n16551) );
  AND U24829 ( .A(n16553), .B(n16554), .Z(o[2551]) );
  AND U24830 ( .A(p_input[22551]), .B(p_input[12551]), .Z(n16554) );
  AND U24831 ( .A(p_input[32551]), .B(p_input[2551]), .Z(n16553) );
  AND U24832 ( .A(n16555), .B(n16556), .Z(o[2550]) );
  AND U24833 ( .A(p_input[22550]), .B(p_input[12550]), .Z(n16556) );
  AND U24834 ( .A(p_input[32550]), .B(p_input[2550]), .Z(n16555) );
  AND U24835 ( .A(n16557), .B(n16558), .Z(o[254]) );
  AND U24836 ( .A(p_input[20254]), .B(p_input[10254]), .Z(n16558) );
  AND U24837 ( .A(p_input[30254]), .B(p_input[254]), .Z(n16557) );
  AND U24838 ( .A(n16559), .B(n16560), .Z(o[2549]) );
  AND U24839 ( .A(p_input[22549]), .B(p_input[12549]), .Z(n16560) );
  AND U24840 ( .A(p_input[32549]), .B(p_input[2549]), .Z(n16559) );
  AND U24841 ( .A(n16561), .B(n16562), .Z(o[2548]) );
  AND U24842 ( .A(p_input[22548]), .B(p_input[12548]), .Z(n16562) );
  AND U24843 ( .A(p_input[32548]), .B(p_input[2548]), .Z(n16561) );
  AND U24844 ( .A(n16563), .B(n16564), .Z(o[2547]) );
  AND U24845 ( .A(p_input[22547]), .B(p_input[12547]), .Z(n16564) );
  AND U24846 ( .A(p_input[32547]), .B(p_input[2547]), .Z(n16563) );
  AND U24847 ( .A(n16565), .B(n16566), .Z(o[2546]) );
  AND U24848 ( .A(p_input[22546]), .B(p_input[12546]), .Z(n16566) );
  AND U24849 ( .A(p_input[32546]), .B(p_input[2546]), .Z(n16565) );
  AND U24850 ( .A(n16567), .B(n16568), .Z(o[2545]) );
  AND U24851 ( .A(p_input[22545]), .B(p_input[12545]), .Z(n16568) );
  AND U24852 ( .A(p_input[32545]), .B(p_input[2545]), .Z(n16567) );
  AND U24853 ( .A(n16569), .B(n16570), .Z(o[2544]) );
  AND U24854 ( .A(p_input[22544]), .B(p_input[12544]), .Z(n16570) );
  AND U24855 ( .A(p_input[32544]), .B(p_input[2544]), .Z(n16569) );
  AND U24856 ( .A(n16571), .B(n16572), .Z(o[2543]) );
  AND U24857 ( .A(p_input[22543]), .B(p_input[12543]), .Z(n16572) );
  AND U24858 ( .A(p_input[32543]), .B(p_input[2543]), .Z(n16571) );
  AND U24859 ( .A(n16573), .B(n16574), .Z(o[2542]) );
  AND U24860 ( .A(p_input[22542]), .B(p_input[12542]), .Z(n16574) );
  AND U24861 ( .A(p_input[32542]), .B(p_input[2542]), .Z(n16573) );
  AND U24862 ( .A(n16575), .B(n16576), .Z(o[2541]) );
  AND U24863 ( .A(p_input[22541]), .B(p_input[12541]), .Z(n16576) );
  AND U24864 ( .A(p_input[32541]), .B(p_input[2541]), .Z(n16575) );
  AND U24865 ( .A(n16577), .B(n16578), .Z(o[2540]) );
  AND U24866 ( .A(p_input[22540]), .B(p_input[12540]), .Z(n16578) );
  AND U24867 ( .A(p_input[32540]), .B(p_input[2540]), .Z(n16577) );
  AND U24868 ( .A(n16579), .B(n16580), .Z(o[253]) );
  AND U24869 ( .A(p_input[20253]), .B(p_input[10253]), .Z(n16580) );
  AND U24870 ( .A(p_input[30253]), .B(p_input[253]), .Z(n16579) );
  AND U24871 ( .A(n16581), .B(n16582), .Z(o[2539]) );
  AND U24872 ( .A(p_input[22539]), .B(p_input[12539]), .Z(n16582) );
  AND U24873 ( .A(p_input[32539]), .B(p_input[2539]), .Z(n16581) );
  AND U24874 ( .A(n16583), .B(n16584), .Z(o[2538]) );
  AND U24875 ( .A(p_input[22538]), .B(p_input[12538]), .Z(n16584) );
  AND U24876 ( .A(p_input[32538]), .B(p_input[2538]), .Z(n16583) );
  AND U24877 ( .A(n16585), .B(n16586), .Z(o[2537]) );
  AND U24878 ( .A(p_input[22537]), .B(p_input[12537]), .Z(n16586) );
  AND U24879 ( .A(p_input[32537]), .B(p_input[2537]), .Z(n16585) );
  AND U24880 ( .A(n16587), .B(n16588), .Z(o[2536]) );
  AND U24881 ( .A(p_input[22536]), .B(p_input[12536]), .Z(n16588) );
  AND U24882 ( .A(p_input[32536]), .B(p_input[2536]), .Z(n16587) );
  AND U24883 ( .A(n16589), .B(n16590), .Z(o[2535]) );
  AND U24884 ( .A(p_input[22535]), .B(p_input[12535]), .Z(n16590) );
  AND U24885 ( .A(p_input[32535]), .B(p_input[2535]), .Z(n16589) );
  AND U24886 ( .A(n16591), .B(n16592), .Z(o[2534]) );
  AND U24887 ( .A(p_input[22534]), .B(p_input[12534]), .Z(n16592) );
  AND U24888 ( .A(p_input[32534]), .B(p_input[2534]), .Z(n16591) );
  AND U24889 ( .A(n16593), .B(n16594), .Z(o[2533]) );
  AND U24890 ( .A(p_input[22533]), .B(p_input[12533]), .Z(n16594) );
  AND U24891 ( .A(p_input[32533]), .B(p_input[2533]), .Z(n16593) );
  AND U24892 ( .A(n16595), .B(n16596), .Z(o[2532]) );
  AND U24893 ( .A(p_input[22532]), .B(p_input[12532]), .Z(n16596) );
  AND U24894 ( .A(p_input[32532]), .B(p_input[2532]), .Z(n16595) );
  AND U24895 ( .A(n16597), .B(n16598), .Z(o[2531]) );
  AND U24896 ( .A(p_input[22531]), .B(p_input[12531]), .Z(n16598) );
  AND U24897 ( .A(p_input[32531]), .B(p_input[2531]), .Z(n16597) );
  AND U24898 ( .A(n16599), .B(n16600), .Z(o[2530]) );
  AND U24899 ( .A(p_input[22530]), .B(p_input[12530]), .Z(n16600) );
  AND U24900 ( .A(p_input[32530]), .B(p_input[2530]), .Z(n16599) );
  AND U24901 ( .A(n16601), .B(n16602), .Z(o[252]) );
  AND U24902 ( .A(p_input[20252]), .B(p_input[10252]), .Z(n16602) );
  AND U24903 ( .A(p_input[30252]), .B(p_input[252]), .Z(n16601) );
  AND U24904 ( .A(n16603), .B(n16604), .Z(o[2529]) );
  AND U24905 ( .A(p_input[22529]), .B(p_input[12529]), .Z(n16604) );
  AND U24906 ( .A(p_input[32529]), .B(p_input[2529]), .Z(n16603) );
  AND U24907 ( .A(n16605), .B(n16606), .Z(o[2528]) );
  AND U24908 ( .A(p_input[22528]), .B(p_input[12528]), .Z(n16606) );
  AND U24909 ( .A(p_input[32528]), .B(p_input[2528]), .Z(n16605) );
  AND U24910 ( .A(n16607), .B(n16608), .Z(o[2527]) );
  AND U24911 ( .A(p_input[22527]), .B(p_input[12527]), .Z(n16608) );
  AND U24912 ( .A(p_input[32527]), .B(p_input[2527]), .Z(n16607) );
  AND U24913 ( .A(n16609), .B(n16610), .Z(o[2526]) );
  AND U24914 ( .A(p_input[22526]), .B(p_input[12526]), .Z(n16610) );
  AND U24915 ( .A(p_input[32526]), .B(p_input[2526]), .Z(n16609) );
  AND U24916 ( .A(n16611), .B(n16612), .Z(o[2525]) );
  AND U24917 ( .A(p_input[22525]), .B(p_input[12525]), .Z(n16612) );
  AND U24918 ( .A(p_input[32525]), .B(p_input[2525]), .Z(n16611) );
  AND U24919 ( .A(n16613), .B(n16614), .Z(o[2524]) );
  AND U24920 ( .A(p_input[22524]), .B(p_input[12524]), .Z(n16614) );
  AND U24921 ( .A(p_input[32524]), .B(p_input[2524]), .Z(n16613) );
  AND U24922 ( .A(n16615), .B(n16616), .Z(o[2523]) );
  AND U24923 ( .A(p_input[22523]), .B(p_input[12523]), .Z(n16616) );
  AND U24924 ( .A(p_input[32523]), .B(p_input[2523]), .Z(n16615) );
  AND U24925 ( .A(n16617), .B(n16618), .Z(o[2522]) );
  AND U24926 ( .A(p_input[22522]), .B(p_input[12522]), .Z(n16618) );
  AND U24927 ( .A(p_input[32522]), .B(p_input[2522]), .Z(n16617) );
  AND U24928 ( .A(n16619), .B(n16620), .Z(o[2521]) );
  AND U24929 ( .A(p_input[22521]), .B(p_input[12521]), .Z(n16620) );
  AND U24930 ( .A(p_input[32521]), .B(p_input[2521]), .Z(n16619) );
  AND U24931 ( .A(n16621), .B(n16622), .Z(o[2520]) );
  AND U24932 ( .A(p_input[22520]), .B(p_input[12520]), .Z(n16622) );
  AND U24933 ( .A(p_input[32520]), .B(p_input[2520]), .Z(n16621) );
  AND U24934 ( .A(n16623), .B(n16624), .Z(o[251]) );
  AND U24935 ( .A(p_input[20251]), .B(p_input[10251]), .Z(n16624) );
  AND U24936 ( .A(p_input[30251]), .B(p_input[251]), .Z(n16623) );
  AND U24937 ( .A(n16625), .B(n16626), .Z(o[2519]) );
  AND U24938 ( .A(p_input[22519]), .B(p_input[12519]), .Z(n16626) );
  AND U24939 ( .A(p_input[32519]), .B(p_input[2519]), .Z(n16625) );
  AND U24940 ( .A(n16627), .B(n16628), .Z(o[2518]) );
  AND U24941 ( .A(p_input[22518]), .B(p_input[12518]), .Z(n16628) );
  AND U24942 ( .A(p_input[32518]), .B(p_input[2518]), .Z(n16627) );
  AND U24943 ( .A(n16629), .B(n16630), .Z(o[2517]) );
  AND U24944 ( .A(p_input[22517]), .B(p_input[12517]), .Z(n16630) );
  AND U24945 ( .A(p_input[32517]), .B(p_input[2517]), .Z(n16629) );
  AND U24946 ( .A(n16631), .B(n16632), .Z(o[2516]) );
  AND U24947 ( .A(p_input[22516]), .B(p_input[12516]), .Z(n16632) );
  AND U24948 ( .A(p_input[32516]), .B(p_input[2516]), .Z(n16631) );
  AND U24949 ( .A(n16633), .B(n16634), .Z(o[2515]) );
  AND U24950 ( .A(p_input[22515]), .B(p_input[12515]), .Z(n16634) );
  AND U24951 ( .A(p_input[32515]), .B(p_input[2515]), .Z(n16633) );
  AND U24952 ( .A(n16635), .B(n16636), .Z(o[2514]) );
  AND U24953 ( .A(p_input[22514]), .B(p_input[12514]), .Z(n16636) );
  AND U24954 ( .A(p_input[32514]), .B(p_input[2514]), .Z(n16635) );
  AND U24955 ( .A(n16637), .B(n16638), .Z(o[2513]) );
  AND U24956 ( .A(p_input[22513]), .B(p_input[12513]), .Z(n16638) );
  AND U24957 ( .A(p_input[32513]), .B(p_input[2513]), .Z(n16637) );
  AND U24958 ( .A(n16639), .B(n16640), .Z(o[2512]) );
  AND U24959 ( .A(p_input[22512]), .B(p_input[12512]), .Z(n16640) );
  AND U24960 ( .A(p_input[32512]), .B(p_input[2512]), .Z(n16639) );
  AND U24961 ( .A(n16641), .B(n16642), .Z(o[2511]) );
  AND U24962 ( .A(p_input[22511]), .B(p_input[12511]), .Z(n16642) );
  AND U24963 ( .A(p_input[32511]), .B(p_input[2511]), .Z(n16641) );
  AND U24964 ( .A(n16643), .B(n16644), .Z(o[2510]) );
  AND U24965 ( .A(p_input[22510]), .B(p_input[12510]), .Z(n16644) );
  AND U24966 ( .A(p_input[32510]), .B(p_input[2510]), .Z(n16643) );
  AND U24967 ( .A(n16645), .B(n16646), .Z(o[250]) );
  AND U24968 ( .A(p_input[20250]), .B(p_input[10250]), .Z(n16646) );
  AND U24969 ( .A(p_input[30250]), .B(p_input[250]), .Z(n16645) );
  AND U24970 ( .A(n16647), .B(n16648), .Z(o[2509]) );
  AND U24971 ( .A(p_input[22509]), .B(p_input[12509]), .Z(n16648) );
  AND U24972 ( .A(p_input[32509]), .B(p_input[2509]), .Z(n16647) );
  AND U24973 ( .A(n16649), .B(n16650), .Z(o[2508]) );
  AND U24974 ( .A(p_input[22508]), .B(p_input[12508]), .Z(n16650) );
  AND U24975 ( .A(p_input[32508]), .B(p_input[2508]), .Z(n16649) );
  AND U24976 ( .A(n16651), .B(n16652), .Z(o[2507]) );
  AND U24977 ( .A(p_input[22507]), .B(p_input[12507]), .Z(n16652) );
  AND U24978 ( .A(p_input[32507]), .B(p_input[2507]), .Z(n16651) );
  AND U24979 ( .A(n16653), .B(n16654), .Z(o[2506]) );
  AND U24980 ( .A(p_input[22506]), .B(p_input[12506]), .Z(n16654) );
  AND U24981 ( .A(p_input[32506]), .B(p_input[2506]), .Z(n16653) );
  AND U24982 ( .A(n16655), .B(n16656), .Z(o[2505]) );
  AND U24983 ( .A(p_input[22505]), .B(p_input[12505]), .Z(n16656) );
  AND U24984 ( .A(p_input[32505]), .B(p_input[2505]), .Z(n16655) );
  AND U24985 ( .A(n16657), .B(n16658), .Z(o[2504]) );
  AND U24986 ( .A(p_input[22504]), .B(p_input[12504]), .Z(n16658) );
  AND U24987 ( .A(p_input[32504]), .B(p_input[2504]), .Z(n16657) );
  AND U24988 ( .A(n16659), .B(n16660), .Z(o[2503]) );
  AND U24989 ( .A(p_input[22503]), .B(p_input[12503]), .Z(n16660) );
  AND U24990 ( .A(p_input[32503]), .B(p_input[2503]), .Z(n16659) );
  AND U24991 ( .A(n16661), .B(n16662), .Z(o[2502]) );
  AND U24992 ( .A(p_input[22502]), .B(p_input[12502]), .Z(n16662) );
  AND U24993 ( .A(p_input[32502]), .B(p_input[2502]), .Z(n16661) );
  AND U24994 ( .A(n16663), .B(n16664), .Z(o[2501]) );
  AND U24995 ( .A(p_input[22501]), .B(p_input[12501]), .Z(n16664) );
  AND U24996 ( .A(p_input[32501]), .B(p_input[2501]), .Z(n16663) );
  AND U24997 ( .A(n16665), .B(n16666), .Z(o[2500]) );
  AND U24998 ( .A(p_input[22500]), .B(p_input[12500]), .Z(n16666) );
  AND U24999 ( .A(p_input[32500]), .B(p_input[2500]), .Z(n16665) );
  AND U25000 ( .A(n16667), .B(n16668), .Z(o[24]) );
  AND U25001 ( .A(p_input[20024]), .B(p_input[10024]), .Z(n16668) );
  AND U25002 ( .A(p_input[30024]), .B(p_input[24]), .Z(n16667) );
  AND U25003 ( .A(n16669), .B(n16670), .Z(o[249]) );
  AND U25004 ( .A(p_input[20249]), .B(p_input[10249]), .Z(n16670) );
  AND U25005 ( .A(p_input[30249]), .B(p_input[249]), .Z(n16669) );
  AND U25006 ( .A(n16671), .B(n16672), .Z(o[2499]) );
  AND U25007 ( .A(p_input[22499]), .B(p_input[12499]), .Z(n16672) );
  AND U25008 ( .A(p_input[32499]), .B(p_input[2499]), .Z(n16671) );
  AND U25009 ( .A(n16673), .B(n16674), .Z(o[2498]) );
  AND U25010 ( .A(p_input[22498]), .B(p_input[12498]), .Z(n16674) );
  AND U25011 ( .A(p_input[32498]), .B(p_input[2498]), .Z(n16673) );
  AND U25012 ( .A(n16675), .B(n16676), .Z(o[2497]) );
  AND U25013 ( .A(p_input[22497]), .B(p_input[12497]), .Z(n16676) );
  AND U25014 ( .A(p_input[32497]), .B(p_input[2497]), .Z(n16675) );
  AND U25015 ( .A(n16677), .B(n16678), .Z(o[2496]) );
  AND U25016 ( .A(p_input[22496]), .B(p_input[12496]), .Z(n16678) );
  AND U25017 ( .A(p_input[32496]), .B(p_input[2496]), .Z(n16677) );
  AND U25018 ( .A(n16679), .B(n16680), .Z(o[2495]) );
  AND U25019 ( .A(p_input[22495]), .B(p_input[12495]), .Z(n16680) );
  AND U25020 ( .A(p_input[32495]), .B(p_input[2495]), .Z(n16679) );
  AND U25021 ( .A(n16681), .B(n16682), .Z(o[2494]) );
  AND U25022 ( .A(p_input[22494]), .B(p_input[12494]), .Z(n16682) );
  AND U25023 ( .A(p_input[32494]), .B(p_input[2494]), .Z(n16681) );
  AND U25024 ( .A(n16683), .B(n16684), .Z(o[2493]) );
  AND U25025 ( .A(p_input[22493]), .B(p_input[12493]), .Z(n16684) );
  AND U25026 ( .A(p_input[32493]), .B(p_input[2493]), .Z(n16683) );
  AND U25027 ( .A(n16685), .B(n16686), .Z(o[2492]) );
  AND U25028 ( .A(p_input[22492]), .B(p_input[12492]), .Z(n16686) );
  AND U25029 ( .A(p_input[32492]), .B(p_input[2492]), .Z(n16685) );
  AND U25030 ( .A(n16687), .B(n16688), .Z(o[2491]) );
  AND U25031 ( .A(p_input[22491]), .B(p_input[12491]), .Z(n16688) );
  AND U25032 ( .A(p_input[32491]), .B(p_input[2491]), .Z(n16687) );
  AND U25033 ( .A(n16689), .B(n16690), .Z(o[2490]) );
  AND U25034 ( .A(p_input[22490]), .B(p_input[12490]), .Z(n16690) );
  AND U25035 ( .A(p_input[32490]), .B(p_input[2490]), .Z(n16689) );
  AND U25036 ( .A(n16691), .B(n16692), .Z(o[248]) );
  AND U25037 ( .A(p_input[20248]), .B(p_input[10248]), .Z(n16692) );
  AND U25038 ( .A(p_input[30248]), .B(p_input[248]), .Z(n16691) );
  AND U25039 ( .A(n16693), .B(n16694), .Z(o[2489]) );
  AND U25040 ( .A(p_input[22489]), .B(p_input[12489]), .Z(n16694) );
  AND U25041 ( .A(p_input[32489]), .B(p_input[2489]), .Z(n16693) );
  AND U25042 ( .A(n16695), .B(n16696), .Z(o[2488]) );
  AND U25043 ( .A(p_input[22488]), .B(p_input[12488]), .Z(n16696) );
  AND U25044 ( .A(p_input[32488]), .B(p_input[2488]), .Z(n16695) );
  AND U25045 ( .A(n16697), .B(n16698), .Z(o[2487]) );
  AND U25046 ( .A(p_input[22487]), .B(p_input[12487]), .Z(n16698) );
  AND U25047 ( .A(p_input[32487]), .B(p_input[2487]), .Z(n16697) );
  AND U25048 ( .A(n16699), .B(n16700), .Z(o[2486]) );
  AND U25049 ( .A(p_input[22486]), .B(p_input[12486]), .Z(n16700) );
  AND U25050 ( .A(p_input[32486]), .B(p_input[2486]), .Z(n16699) );
  AND U25051 ( .A(n16701), .B(n16702), .Z(o[2485]) );
  AND U25052 ( .A(p_input[22485]), .B(p_input[12485]), .Z(n16702) );
  AND U25053 ( .A(p_input[32485]), .B(p_input[2485]), .Z(n16701) );
  AND U25054 ( .A(n16703), .B(n16704), .Z(o[2484]) );
  AND U25055 ( .A(p_input[22484]), .B(p_input[12484]), .Z(n16704) );
  AND U25056 ( .A(p_input[32484]), .B(p_input[2484]), .Z(n16703) );
  AND U25057 ( .A(n16705), .B(n16706), .Z(o[2483]) );
  AND U25058 ( .A(p_input[22483]), .B(p_input[12483]), .Z(n16706) );
  AND U25059 ( .A(p_input[32483]), .B(p_input[2483]), .Z(n16705) );
  AND U25060 ( .A(n16707), .B(n16708), .Z(o[2482]) );
  AND U25061 ( .A(p_input[22482]), .B(p_input[12482]), .Z(n16708) );
  AND U25062 ( .A(p_input[32482]), .B(p_input[2482]), .Z(n16707) );
  AND U25063 ( .A(n16709), .B(n16710), .Z(o[2481]) );
  AND U25064 ( .A(p_input[22481]), .B(p_input[12481]), .Z(n16710) );
  AND U25065 ( .A(p_input[32481]), .B(p_input[2481]), .Z(n16709) );
  AND U25066 ( .A(n16711), .B(n16712), .Z(o[2480]) );
  AND U25067 ( .A(p_input[22480]), .B(p_input[12480]), .Z(n16712) );
  AND U25068 ( .A(p_input[32480]), .B(p_input[2480]), .Z(n16711) );
  AND U25069 ( .A(n16713), .B(n16714), .Z(o[247]) );
  AND U25070 ( .A(p_input[20247]), .B(p_input[10247]), .Z(n16714) );
  AND U25071 ( .A(p_input[30247]), .B(p_input[247]), .Z(n16713) );
  AND U25072 ( .A(n16715), .B(n16716), .Z(o[2479]) );
  AND U25073 ( .A(p_input[22479]), .B(p_input[12479]), .Z(n16716) );
  AND U25074 ( .A(p_input[32479]), .B(p_input[2479]), .Z(n16715) );
  AND U25075 ( .A(n16717), .B(n16718), .Z(o[2478]) );
  AND U25076 ( .A(p_input[22478]), .B(p_input[12478]), .Z(n16718) );
  AND U25077 ( .A(p_input[32478]), .B(p_input[2478]), .Z(n16717) );
  AND U25078 ( .A(n16719), .B(n16720), .Z(o[2477]) );
  AND U25079 ( .A(p_input[22477]), .B(p_input[12477]), .Z(n16720) );
  AND U25080 ( .A(p_input[32477]), .B(p_input[2477]), .Z(n16719) );
  AND U25081 ( .A(n16721), .B(n16722), .Z(o[2476]) );
  AND U25082 ( .A(p_input[22476]), .B(p_input[12476]), .Z(n16722) );
  AND U25083 ( .A(p_input[32476]), .B(p_input[2476]), .Z(n16721) );
  AND U25084 ( .A(n16723), .B(n16724), .Z(o[2475]) );
  AND U25085 ( .A(p_input[22475]), .B(p_input[12475]), .Z(n16724) );
  AND U25086 ( .A(p_input[32475]), .B(p_input[2475]), .Z(n16723) );
  AND U25087 ( .A(n16725), .B(n16726), .Z(o[2474]) );
  AND U25088 ( .A(p_input[22474]), .B(p_input[12474]), .Z(n16726) );
  AND U25089 ( .A(p_input[32474]), .B(p_input[2474]), .Z(n16725) );
  AND U25090 ( .A(n16727), .B(n16728), .Z(o[2473]) );
  AND U25091 ( .A(p_input[22473]), .B(p_input[12473]), .Z(n16728) );
  AND U25092 ( .A(p_input[32473]), .B(p_input[2473]), .Z(n16727) );
  AND U25093 ( .A(n16729), .B(n16730), .Z(o[2472]) );
  AND U25094 ( .A(p_input[22472]), .B(p_input[12472]), .Z(n16730) );
  AND U25095 ( .A(p_input[32472]), .B(p_input[2472]), .Z(n16729) );
  AND U25096 ( .A(n16731), .B(n16732), .Z(o[2471]) );
  AND U25097 ( .A(p_input[22471]), .B(p_input[12471]), .Z(n16732) );
  AND U25098 ( .A(p_input[32471]), .B(p_input[2471]), .Z(n16731) );
  AND U25099 ( .A(n16733), .B(n16734), .Z(o[2470]) );
  AND U25100 ( .A(p_input[22470]), .B(p_input[12470]), .Z(n16734) );
  AND U25101 ( .A(p_input[32470]), .B(p_input[2470]), .Z(n16733) );
  AND U25102 ( .A(n16735), .B(n16736), .Z(o[246]) );
  AND U25103 ( .A(p_input[20246]), .B(p_input[10246]), .Z(n16736) );
  AND U25104 ( .A(p_input[30246]), .B(p_input[246]), .Z(n16735) );
  AND U25105 ( .A(n16737), .B(n16738), .Z(o[2469]) );
  AND U25106 ( .A(p_input[22469]), .B(p_input[12469]), .Z(n16738) );
  AND U25107 ( .A(p_input[32469]), .B(p_input[2469]), .Z(n16737) );
  AND U25108 ( .A(n16739), .B(n16740), .Z(o[2468]) );
  AND U25109 ( .A(p_input[22468]), .B(p_input[12468]), .Z(n16740) );
  AND U25110 ( .A(p_input[32468]), .B(p_input[2468]), .Z(n16739) );
  AND U25111 ( .A(n16741), .B(n16742), .Z(o[2467]) );
  AND U25112 ( .A(p_input[22467]), .B(p_input[12467]), .Z(n16742) );
  AND U25113 ( .A(p_input[32467]), .B(p_input[2467]), .Z(n16741) );
  AND U25114 ( .A(n16743), .B(n16744), .Z(o[2466]) );
  AND U25115 ( .A(p_input[22466]), .B(p_input[12466]), .Z(n16744) );
  AND U25116 ( .A(p_input[32466]), .B(p_input[2466]), .Z(n16743) );
  AND U25117 ( .A(n16745), .B(n16746), .Z(o[2465]) );
  AND U25118 ( .A(p_input[22465]), .B(p_input[12465]), .Z(n16746) );
  AND U25119 ( .A(p_input[32465]), .B(p_input[2465]), .Z(n16745) );
  AND U25120 ( .A(n16747), .B(n16748), .Z(o[2464]) );
  AND U25121 ( .A(p_input[22464]), .B(p_input[12464]), .Z(n16748) );
  AND U25122 ( .A(p_input[32464]), .B(p_input[2464]), .Z(n16747) );
  AND U25123 ( .A(n16749), .B(n16750), .Z(o[2463]) );
  AND U25124 ( .A(p_input[22463]), .B(p_input[12463]), .Z(n16750) );
  AND U25125 ( .A(p_input[32463]), .B(p_input[2463]), .Z(n16749) );
  AND U25126 ( .A(n16751), .B(n16752), .Z(o[2462]) );
  AND U25127 ( .A(p_input[22462]), .B(p_input[12462]), .Z(n16752) );
  AND U25128 ( .A(p_input[32462]), .B(p_input[2462]), .Z(n16751) );
  AND U25129 ( .A(n16753), .B(n16754), .Z(o[2461]) );
  AND U25130 ( .A(p_input[22461]), .B(p_input[12461]), .Z(n16754) );
  AND U25131 ( .A(p_input[32461]), .B(p_input[2461]), .Z(n16753) );
  AND U25132 ( .A(n16755), .B(n16756), .Z(o[2460]) );
  AND U25133 ( .A(p_input[22460]), .B(p_input[12460]), .Z(n16756) );
  AND U25134 ( .A(p_input[32460]), .B(p_input[2460]), .Z(n16755) );
  AND U25135 ( .A(n16757), .B(n16758), .Z(o[245]) );
  AND U25136 ( .A(p_input[20245]), .B(p_input[10245]), .Z(n16758) );
  AND U25137 ( .A(p_input[30245]), .B(p_input[245]), .Z(n16757) );
  AND U25138 ( .A(n16759), .B(n16760), .Z(o[2459]) );
  AND U25139 ( .A(p_input[22459]), .B(p_input[12459]), .Z(n16760) );
  AND U25140 ( .A(p_input[32459]), .B(p_input[2459]), .Z(n16759) );
  AND U25141 ( .A(n16761), .B(n16762), .Z(o[2458]) );
  AND U25142 ( .A(p_input[22458]), .B(p_input[12458]), .Z(n16762) );
  AND U25143 ( .A(p_input[32458]), .B(p_input[2458]), .Z(n16761) );
  AND U25144 ( .A(n16763), .B(n16764), .Z(o[2457]) );
  AND U25145 ( .A(p_input[22457]), .B(p_input[12457]), .Z(n16764) );
  AND U25146 ( .A(p_input[32457]), .B(p_input[2457]), .Z(n16763) );
  AND U25147 ( .A(n16765), .B(n16766), .Z(o[2456]) );
  AND U25148 ( .A(p_input[22456]), .B(p_input[12456]), .Z(n16766) );
  AND U25149 ( .A(p_input[32456]), .B(p_input[2456]), .Z(n16765) );
  AND U25150 ( .A(n16767), .B(n16768), .Z(o[2455]) );
  AND U25151 ( .A(p_input[22455]), .B(p_input[12455]), .Z(n16768) );
  AND U25152 ( .A(p_input[32455]), .B(p_input[2455]), .Z(n16767) );
  AND U25153 ( .A(n16769), .B(n16770), .Z(o[2454]) );
  AND U25154 ( .A(p_input[22454]), .B(p_input[12454]), .Z(n16770) );
  AND U25155 ( .A(p_input[32454]), .B(p_input[2454]), .Z(n16769) );
  AND U25156 ( .A(n16771), .B(n16772), .Z(o[2453]) );
  AND U25157 ( .A(p_input[22453]), .B(p_input[12453]), .Z(n16772) );
  AND U25158 ( .A(p_input[32453]), .B(p_input[2453]), .Z(n16771) );
  AND U25159 ( .A(n16773), .B(n16774), .Z(o[2452]) );
  AND U25160 ( .A(p_input[22452]), .B(p_input[12452]), .Z(n16774) );
  AND U25161 ( .A(p_input[32452]), .B(p_input[2452]), .Z(n16773) );
  AND U25162 ( .A(n16775), .B(n16776), .Z(o[2451]) );
  AND U25163 ( .A(p_input[22451]), .B(p_input[12451]), .Z(n16776) );
  AND U25164 ( .A(p_input[32451]), .B(p_input[2451]), .Z(n16775) );
  AND U25165 ( .A(n16777), .B(n16778), .Z(o[2450]) );
  AND U25166 ( .A(p_input[22450]), .B(p_input[12450]), .Z(n16778) );
  AND U25167 ( .A(p_input[32450]), .B(p_input[2450]), .Z(n16777) );
  AND U25168 ( .A(n16779), .B(n16780), .Z(o[244]) );
  AND U25169 ( .A(p_input[20244]), .B(p_input[10244]), .Z(n16780) );
  AND U25170 ( .A(p_input[30244]), .B(p_input[244]), .Z(n16779) );
  AND U25171 ( .A(n16781), .B(n16782), .Z(o[2449]) );
  AND U25172 ( .A(p_input[22449]), .B(p_input[12449]), .Z(n16782) );
  AND U25173 ( .A(p_input[32449]), .B(p_input[2449]), .Z(n16781) );
  AND U25174 ( .A(n16783), .B(n16784), .Z(o[2448]) );
  AND U25175 ( .A(p_input[22448]), .B(p_input[12448]), .Z(n16784) );
  AND U25176 ( .A(p_input[32448]), .B(p_input[2448]), .Z(n16783) );
  AND U25177 ( .A(n16785), .B(n16786), .Z(o[2447]) );
  AND U25178 ( .A(p_input[22447]), .B(p_input[12447]), .Z(n16786) );
  AND U25179 ( .A(p_input[32447]), .B(p_input[2447]), .Z(n16785) );
  AND U25180 ( .A(n16787), .B(n16788), .Z(o[2446]) );
  AND U25181 ( .A(p_input[22446]), .B(p_input[12446]), .Z(n16788) );
  AND U25182 ( .A(p_input[32446]), .B(p_input[2446]), .Z(n16787) );
  AND U25183 ( .A(n16789), .B(n16790), .Z(o[2445]) );
  AND U25184 ( .A(p_input[22445]), .B(p_input[12445]), .Z(n16790) );
  AND U25185 ( .A(p_input[32445]), .B(p_input[2445]), .Z(n16789) );
  AND U25186 ( .A(n16791), .B(n16792), .Z(o[2444]) );
  AND U25187 ( .A(p_input[22444]), .B(p_input[12444]), .Z(n16792) );
  AND U25188 ( .A(p_input[32444]), .B(p_input[2444]), .Z(n16791) );
  AND U25189 ( .A(n16793), .B(n16794), .Z(o[2443]) );
  AND U25190 ( .A(p_input[22443]), .B(p_input[12443]), .Z(n16794) );
  AND U25191 ( .A(p_input[32443]), .B(p_input[2443]), .Z(n16793) );
  AND U25192 ( .A(n16795), .B(n16796), .Z(o[2442]) );
  AND U25193 ( .A(p_input[22442]), .B(p_input[12442]), .Z(n16796) );
  AND U25194 ( .A(p_input[32442]), .B(p_input[2442]), .Z(n16795) );
  AND U25195 ( .A(n16797), .B(n16798), .Z(o[2441]) );
  AND U25196 ( .A(p_input[22441]), .B(p_input[12441]), .Z(n16798) );
  AND U25197 ( .A(p_input[32441]), .B(p_input[2441]), .Z(n16797) );
  AND U25198 ( .A(n16799), .B(n16800), .Z(o[2440]) );
  AND U25199 ( .A(p_input[22440]), .B(p_input[12440]), .Z(n16800) );
  AND U25200 ( .A(p_input[32440]), .B(p_input[2440]), .Z(n16799) );
  AND U25201 ( .A(n16801), .B(n16802), .Z(o[243]) );
  AND U25202 ( .A(p_input[20243]), .B(p_input[10243]), .Z(n16802) );
  AND U25203 ( .A(p_input[30243]), .B(p_input[243]), .Z(n16801) );
  AND U25204 ( .A(n16803), .B(n16804), .Z(o[2439]) );
  AND U25205 ( .A(p_input[22439]), .B(p_input[12439]), .Z(n16804) );
  AND U25206 ( .A(p_input[32439]), .B(p_input[2439]), .Z(n16803) );
  AND U25207 ( .A(n16805), .B(n16806), .Z(o[2438]) );
  AND U25208 ( .A(p_input[22438]), .B(p_input[12438]), .Z(n16806) );
  AND U25209 ( .A(p_input[32438]), .B(p_input[2438]), .Z(n16805) );
  AND U25210 ( .A(n16807), .B(n16808), .Z(o[2437]) );
  AND U25211 ( .A(p_input[22437]), .B(p_input[12437]), .Z(n16808) );
  AND U25212 ( .A(p_input[32437]), .B(p_input[2437]), .Z(n16807) );
  AND U25213 ( .A(n16809), .B(n16810), .Z(o[2436]) );
  AND U25214 ( .A(p_input[22436]), .B(p_input[12436]), .Z(n16810) );
  AND U25215 ( .A(p_input[32436]), .B(p_input[2436]), .Z(n16809) );
  AND U25216 ( .A(n16811), .B(n16812), .Z(o[2435]) );
  AND U25217 ( .A(p_input[22435]), .B(p_input[12435]), .Z(n16812) );
  AND U25218 ( .A(p_input[32435]), .B(p_input[2435]), .Z(n16811) );
  AND U25219 ( .A(n16813), .B(n16814), .Z(o[2434]) );
  AND U25220 ( .A(p_input[22434]), .B(p_input[12434]), .Z(n16814) );
  AND U25221 ( .A(p_input[32434]), .B(p_input[2434]), .Z(n16813) );
  AND U25222 ( .A(n16815), .B(n16816), .Z(o[2433]) );
  AND U25223 ( .A(p_input[22433]), .B(p_input[12433]), .Z(n16816) );
  AND U25224 ( .A(p_input[32433]), .B(p_input[2433]), .Z(n16815) );
  AND U25225 ( .A(n16817), .B(n16818), .Z(o[2432]) );
  AND U25226 ( .A(p_input[22432]), .B(p_input[12432]), .Z(n16818) );
  AND U25227 ( .A(p_input[32432]), .B(p_input[2432]), .Z(n16817) );
  AND U25228 ( .A(n16819), .B(n16820), .Z(o[2431]) );
  AND U25229 ( .A(p_input[22431]), .B(p_input[12431]), .Z(n16820) );
  AND U25230 ( .A(p_input[32431]), .B(p_input[2431]), .Z(n16819) );
  AND U25231 ( .A(n16821), .B(n16822), .Z(o[2430]) );
  AND U25232 ( .A(p_input[22430]), .B(p_input[12430]), .Z(n16822) );
  AND U25233 ( .A(p_input[32430]), .B(p_input[2430]), .Z(n16821) );
  AND U25234 ( .A(n16823), .B(n16824), .Z(o[242]) );
  AND U25235 ( .A(p_input[20242]), .B(p_input[10242]), .Z(n16824) );
  AND U25236 ( .A(p_input[30242]), .B(p_input[242]), .Z(n16823) );
  AND U25237 ( .A(n16825), .B(n16826), .Z(o[2429]) );
  AND U25238 ( .A(p_input[22429]), .B(p_input[12429]), .Z(n16826) );
  AND U25239 ( .A(p_input[32429]), .B(p_input[2429]), .Z(n16825) );
  AND U25240 ( .A(n16827), .B(n16828), .Z(o[2428]) );
  AND U25241 ( .A(p_input[22428]), .B(p_input[12428]), .Z(n16828) );
  AND U25242 ( .A(p_input[32428]), .B(p_input[2428]), .Z(n16827) );
  AND U25243 ( .A(n16829), .B(n16830), .Z(o[2427]) );
  AND U25244 ( .A(p_input[22427]), .B(p_input[12427]), .Z(n16830) );
  AND U25245 ( .A(p_input[32427]), .B(p_input[2427]), .Z(n16829) );
  AND U25246 ( .A(n16831), .B(n16832), .Z(o[2426]) );
  AND U25247 ( .A(p_input[22426]), .B(p_input[12426]), .Z(n16832) );
  AND U25248 ( .A(p_input[32426]), .B(p_input[2426]), .Z(n16831) );
  AND U25249 ( .A(n16833), .B(n16834), .Z(o[2425]) );
  AND U25250 ( .A(p_input[22425]), .B(p_input[12425]), .Z(n16834) );
  AND U25251 ( .A(p_input[32425]), .B(p_input[2425]), .Z(n16833) );
  AND U25252 ( .A(n16835), .B(n16836), .Z(o[2424]) );
  AND U25253 ( .A(p_input[22424]), .B(p_input[12424]), .Z(n16836) );
  AND U25254 ( .A(p_input[32424]), .B(p_input[2424]), .Z(n16835) );
  AND U25255 ( .A(n16837), .B(n16838), .Z(o[2423]) );
  AND U25256 ( .A(p_input[22423]), .B(p_input[12423]), .Z(n16838) );
  AND U25257 ( .A(p_input[32423]), .B(p_input[2423]), .Z(n16837) );
  AND U25258 ( .A(n16839), .B(n16840), .Z(o[2422]) );
  AND U25259 ( .A(p_input[22422]), .B(p_input[12422]), .Z(n16840) );
  AND U25260 ( .A(p_input[32422]), .B(p_input[2422]), .Z(n16839) );
  AND U25261 ( .A(n16841), .B(n16842), .Z(o[2421]) );
  AND U25262 ( .A(p_input[22421]), .B(p_input[12421]), .Z(n16842) );
  AND U25263 ( .A(p_input[32421]), .B(p_input[2421]), .Z(n16841) );
  AND U25264 ( .A(n16843), .B(n16844), .Z(o[2420]) );
  AND U25265 ( .A(p_input[22420]), .B(p_input[12420]), .Z(n16844) );
  AND U25266 ( .A(p_input[32420]), .B(p_input[2420]), .Z(n16843) );
  AND U25267 ( .A(n16845), .B(n16846), .Z(o[241]) );
  AND U25268 ( .A(p_input[20241]), .B(p_input[10241]), .Z(n16846) );
  AND U25269 ( .A(p_input[30241]), .B(p_input[241]), .Z(n16845) );
  AND U25270 ( .A(n16847), .B(n16848), .Z(o[2419]) );
  AND U25271 ( .A(p_input[22419]), .B(p_input[12419]), .Z(n16848) );
  AND U25272 ( .A(p_input[32419]), .B(p_input[2419]), .Z(n16847) );
  AND U25273 ( .A(n16849), .B(n16850), .Z(o[2418]) );
  AND U25274 ( .A(p_input[22418]), .B(p_input[12418]), .Z(n16850) );
  AND U25275 ( .A(p_input[32418]), .B(p_input[2418]), .Z(n16849) );
  AND U25276 ( .A(n16851), .B(n16852), .Z(o[2417]) );
  AND U25277 ( .A(p_input[22417]), .B(p_input[12417]), .Z(n16852) );
  AND U25278 ( .A(p_input[32417]), .B(p_input[2417]), .Z(n16851) );
  AND U25279 ( .A(n16853), .B(n16854), .Z(o[2416]) );
  AND U25280 ( .A(p_input[22416]), .B(p_input[12416]), .Z(n16854) );
  AND U25281 ( .A(p_input[32416]), .B(p_input[2416]), .Z(n16853) );
  AND U25282 ( .A(n16855), .B(n16856), .Z(o[2415]) );
  AND U25283 ( .A(p_input[22415]), .B(p_input[12415]), .Z(n16856) );
  AND U25284 ( .A(p_input[32415]), .B(p_input[2415]), .Z(n16855) );
  AND U25285 ( .A(n16857), .B(n16858), .Z(o[2414]) );
  AND U25286 ( .A(p_input[22414]), .B(p_input[12414]), .Z(n16858) );
  AND U25287 ( .A(p_input[32414]), .B(p_input[2414]), .Z(n16857) );
  AND U25288 ( .A(n16859), .B(n16860), .Z(o[2413]) );
  AND U25289 ( .A(p_input[22413]), .B(p_input[12413]), .Z(n16860) );
  AND U25290 ( .A(p_input[32413]), .B(p_input[2413]), .Z(n16859) );
  AND U25291 ( .A(n16861), .B(n16862), .Z(o[2412]) );
  AND U25292 ( .A(p_input[22412]), .B(p_input[12412]), .Z(n16862) );
  AND U25293 ( .A(p_input[32412]), .B(p_input[2412]), .Z(n16861) );
  AND U25294 ( .A(n16863), .B(n16864), .Z(o[2411]) );
  AND U25295 ( .A(p_input[22411]), .B(p_input[12411]), .Z(n16864) );
  AND U25296 ( .A(p_input[32411]), .B(p_input[2411]), .Z(n16863) );
  AND U25297 ( .A(n16865), .B(n16866), .Z(o[2410]) );
  AND U25298 ( .A(p_input[22410]), .B(p_input[12410]), .Z(n16866) );
  AND U25299 ( .A(p_input[32410]), .B(p_input[2410]), .Z(n16865) );
  AND U25300 ( .A(n16867), .B(n16868), .Z(o[240]) );
  AND U25301 ( .A(p_input[20240]), .B(p_input[10240]), .Z(n16868) );
  AND U25302 ( .A(p_input[30240]), .B(p_input[240]), .Z(n16867) );
  AND U25303 ( .A(n16869), .B(n16870), .Z(o[2409]) );
  AND U25304 ( .A(p_input[22409]), .B(p_input[12409]), .Z(n16870) );
  AND U25305 ( .A(p_input[32409]), .B(p_input[2409]), .Z(n16869) );
  AND U25306 ( .A(n16871), .B(n16872), .Z(o[2408]) );
  AND U25307 ( .A(p_input[22408]), .B(p_input[12408]), .Z(n16872) );
  AND U25308 ( .A(p_input[32408]), .B(p_input[2408]), .Z(n16871) );
  AND U25309 ( .A(n16873), .B(n16874), .Z(o[2407]) );
  AND U25310 ( .A(p_input[22407]), .B(p_input[12407]), .Z(n16874) );
  AND U25311 ( .A(p_input[32407]), .B(p_input[2407]), .Z(n16873) );
  AND U25312 ( .A(n16875), .B(n16876), .Z(o[2406]) );
  AND U25313 ( .A(p_input[22406]), .B(p_input[12406]), .Z(n16876) );
  AND U25314 ( .A(p_input[32406]), .B(p_input[2406]), .Z(n16875) );
  AND U25315 ( .A(n16877), .B(n16878), .Z(o[2405]) );
  AND U25316 ( .A(p_input[22405]), .B(p_input[12405]), .Z(n16878) );
  AND U25317 ( .A(p_input[32405]), .B(p_input[2405]), .Z(n16877) );
  AND U25318 ( .A(n16879), .B(n16880), .Z(o[2404]) );
  AND U25319 ( .A(p_input[22404]), .B(p_input[12404]), .Z(n16880) );
  AND U25320 ( .A(p_input[32404]), .B(p_input[2404]), .Z(n16879) );
  AND U25321 ( .A(n16881), .B(n16882), .Z(o[2403]) );
  AND U25322 ( .A(p_input[22403]), .B(p_input[12403]), .Z(n16882) );
  AND U25323 ( .A(p_input[32403]), .B(p_input[2403]), .Z(n16881) );
  AND U25324 ( .A(n16883), .B(n16884), .Z(o[2402]) );
  AND U25325 ( .A(p_input[22402]), .B(p_input[12402]), .Z(n16884) );
  AND U25326 ( .A(p_input[32402]), .B(p_input[2402]), .Z(n16883) );
  AND U25327 ( .A(n16885), .B(n16886), .Z(o[2401]) );
  AND U25328 ( .A(p_input[22401]), .B(p_input[12401]), .Z(n16886) );
  AND U25329 ( .A(p_input[32401]), .B(p_input[2401]), .Z(n16885) );
  AND U25330 ( .A(n16887), .B(n16888), .Z(o[2400]) );
  AND U25331 ( .A(p_input[22400]), .B(p_input[12400]), .Z(n16888) );
  AND U25332 ( .A(p_input[32400]), .B(p_input[2400]), .Z(n16887) );
  AND U25333 ( .A(n16889), .B(n16890), .Z(o[23]) );
  AND U25334 ( .A(p_input[20023]), .B(p_input[10023]), .Z(n16890) );
  AND U25335 ( .A(p_input[30023]), .B(p_input[23]), .Z(n16889) );
  AND U25336 ( .A(n16891), .B(n16892), .Z(o[239]) );
  AND U25337 ( .A(p_input[20239]), .B(p_input[10239]), .Z(n16892) );
  AND U25338 ( .A(p_input[30239]), .B(p_input[239]), .Z(n16891) );
  AND U25339 ( .A(n16893), .B(n16894), .Z(o[2399]) );
  AND U25340 ( .A(p_input[22399]), .B(p_input[12399]), .Z(n16894) );
  AND U25341 ( .A(p_input[32399]), .B(p_input[2399]), .Z(n16893) );
  AND U25342 ( .A(n16895), .B(n16896), .Z(o[2398]) );
  AND U25343 ( .A(p_input[22398]), .B(p_input[12398]), .Z(n16896) );
  AND U25344 ( .A(p_input[32398]), .B(p_input[2398]), .Z(n16895) );
  AND U25345 ( .A(n16897), .B(n16898), .Z(o[2397]) );
  AND U25346 ( .A(p_input[22397]), .B(p_input[12397]), .Z(n16898) );
  AND U25347 ( .A(p_input[32397]), .B(p_input[2397]), .Z(n16897) );
  AND U25348 ( .A(n16899), .B(n16900), .Z(o[2396]) );
  AND U25349 ( .A(p_input[22396]), .B(p_input[12396]), .Z(n16900) );
  AND U25350 ( .A(p_input[32396]), .B(p_input[2396]), .Z(n16899) );
  AND U25351 ( .A(n16901), .B(n16902), .Z(o[2395]) );
  AND U25352 ( .A(p_input[22395]), .B(p_input[12395]), .Z(n16902) );
  AND U25353 ( .A(p_input[32395]), .B(p_input[2395]), .Z(n16901) );
  AND U25354 ( .A(n16903), .B(n16904), .Z(o[2394]) );
  AND U25355 ( .A(p_input[22394]), .B(p_input[12394]), .Z(n16904) );
  AND U25356 ( .A(p_input[32394]), .B(p_input[2394]), .Z(n16903) );
  AND U25357 ( .A(n16905), .B(n16906), .Z(o[2393]) );
  AND U25358 ( .A(p_input[22393]), .B(p_input[12393]), .Z(n16906) );
  AND U25359 ( .A(p_input[32393]), .B(p_input[2393]), .Z(n16905) );
  AND U25360 ( .A(n16907), .B(n16908), .Z(o[2392]) );
  AND U25361 ( .A(p_input[22392]), .B(p_input[12392]), .Z(n16908) );
  AND U25362 ( .A(p_input[32392]), .B(p_input[2392]), .Z(n16907) );
  AND U25363 ( .A(n16909), .B(n16910), .Z(o[2391]) );
  AND U25364 ( .A(p_input[22391]), .B(p_input[12391]), .Z(n16910) );
  AND U25365 ( .A(p_input[32391]), .B(p_input[2391]), .Z(n16909) );
  AND U25366 ( .A(n16911), .B(n16912), .Z(o[2390]) );
  AND U25367 ( .A(p_input[22390]), .B(p_input[12390]), .Z(n16912) );
  AND U25368 ( .A(p_input[32390]), .B(p_input[2390]), .Z(n16911) );
  AND U25369 ( .A(n16913), .B(n16914), .Z(o[238]) );
  AND U25370 ( .A(p_input[20238]), .B(p_input[10238]), .Z(n16914) );
  AND U25371 ( .A(p_input[30238]), .B(p_input[238]), .Z(n16913) );
  AND U25372 ( .A(n16915), .B(n16916), .Z(o[2389]) );
  AND U25373 ( .A(p_input[22389]), .B(p_input[12389]), .Z(n16916) );
  AND U25374 ( .A(p_input[32389]), .B(p_input[2389]), .Z(n16915) );
  AND U25375 ( .A(n16917), .B(n16918), .Z(o[2388]) );
  AND U25376 ( .A(p_input[22388]), .B(p_input[12388]), .Z(n16918) );
  AND U25377 ( .A(p_input[32388]), .B(p_input[2388]), .Z(n16917) );
  AND U25378 ( .A(n16919), .B(n16920), .Z(o[2387]) );
  AND U25379 ( .A(p_input[22387]), .B(p_input[12387]), .Z(n16920) );
  AND U25380 ( .A(p_input[32387]), .B(p_input[2387]), .Z(n16919) );
  AND U25381 ( .A(n16921), .B(n16922), .Z(o[2386]) );
  AND U25382 ( .A(p_input[22386]), .B(p_input[12386]), .Z(n16922) );
  AND U25383 ( .A(p_input[32386]), .B(p_input[2386]), .Z(n16921) );
  AND U25384 ( .A(n16923), .B(n16924), .Z(o[2385]) );
  AND U25385 ( .A(p_input[22385]), .B(p_input[12385]), .Z(n16924) );
  AND U25386 ( .A(p_input[32385]), .B(p_input[2385]), .Z(n16923) );
  AND U25387 ( .A(n16925), .B(n16926), .Z(o[2384]) );
  AND U25388 ( .A(p_input[22384]), .B(p_input[12384]), .Z(n16926) );
  AND U25389 ( .A(p_input[32384]), .B(p_input[2384]), .Z(n16925) );
  AND U25390 ( .A(n16927), .B(n16928), .Z(o[2383]) );
  AND U25391 ( .A(p_input[22383]), .B(p_input[12383]), .Z(n16928) );
  AND U25392 ( .A(p_input[32383]), .B(p_input[2383]), .Z(n16927) );
  AND U25393 ( .A(n16929), .B(n16930), .Z(o[2382]) );
  AND U25394 ( .A(p_input[22382]), .B(p_input[12382]), .Z(n16930) );
  AND U25395 ( .A(p_input[32382]), .B(p_input[2382]), .Z(n16929) );
  AND U25396 ( .A(n16931), .B(n16932), .Z(o[2381]) );
  AND U25397 ( .A(p_input[22381]), .B(p_input[12381]), .Z(n16932) );
  AND U25398 ( .A(p_input[32381]), .B(p_input[2381]), .Z(n16931) );
  AND U25399 ( .A(n16933), .B(n16934), .Z(o[2380]) );
  AND U25400 ( .A(p_input[22380]), .B(p_input[12380]), .Z(n16934) );
  AND U25401 ( .A(p_input[32380]), .B(p_input[2380]), .Z(n16933) );
  AND U25402 ( .A(n16935), .B(n16936), .Z(o[237]) );
  AND U25403 ( .A(p_input[20237]), .B(p_input[10237]), .Z(n16936) );
  AND U25404 ( .A(p_input[30237]), .B(p_input[237]), .Z(n16935) );
  AND U25405 ( .A(n16937), .B(n16938), .Z(o[2379]) );
  AND U25406 ( .A(p_input[22379]), .B(p_input[12379]), .Z(n16938) );
  AND U25407 ( .A(p_input[32379]), .B(p_input[2379]), .Z(n16937) );
  AND U25408 ( .A(n16939), .B(n16940), .Z(o[2378]) );
  AND U25409 ( .A(p_input[22378]), .B(p_input[12378]), .Z(n16940) );
  AND U25410 ( .A(p_input[32378]), .B(p_input[2378]), .Z(n16939) );
  AND U25411 ( .A(n16941), .B(n16942), .Z(o[2377]) );
  AND U25412 ( .A(p_input[22377]), .B(p_input[12377]), .Z(n16942) );
  AND U25413 ( .A(p_input[32377]), .B(p_input[2377]), .Z(n16941) );
  AND U25414 ( .A(n16943), .B(n16944), .Z(o[2376]) );
  AND U25415 ( .A(p_input[22376]), .B(p_input[12376]), .Z(n16944) );
  AND U25416 ( .A(p_input[32376]), .B(p_input[2376]), .Z(n16943) );
  AND U25417 ( .A(n16945), .B(n16946), .Z(o[2375]) );
  AND U25418 ( .A(p_input[22375]), .B(p_input[12375]), .Z(n16946) );
  AND U25419 ( .A(p_input[32375]), .B(p_input[2375]), .Z(n16945) );
  AND U25420 ( .A(n16947), .B(n16948), .Z(o[2374]) );
  AND U25421 ( .A(p_input[22374]), .B(p_input[12374]), .Z(n16948) );
  AND U25422 ( .A(p_input[32374]), .B(p_input[2374]), .Z(n16947) );
  AND U25423 ( .A(n16949), .B(n16950), .Z(o[2373]) );
  AND U25424 ( .A(p_input[22373]), .B(p_input[12373]), .Z(n16950) );
  AND U25425 ( .A(p_input[32373]), .B(p_input[2373]), .Z(n16949) );
  AND U25426 ( .A(n16951), .B(n16952), .Z(o[2372]) );
  AND U25427 ( .A(p_input[22372]), .B(p_input[12372]), .Z(n16952) );
  AND U25428 ( .A(p_input[32372]), .B(p_input[2372]), .Z(n16951) );
  AND U25429 ( .A(n16953), .B(n16954), .Z(o[2371]) );
  AND U25430 ( .A(p_input[22371]), .B(p_input[12371]), .Z(n16954) );
  AND U25431 ( .A(p_input[32371]), .B(p_input[2371]), .Z(n16953) );
  AND U25432 ( .A(n16955), .B(n16956), .Z(o[2370]) );
  AND U25433 ( .A(p_input[22370]), .B(p_input[12370]), .Z(n16956) );
  AND U25434 ( .A(p_input[32370]), .B(p_input[2370]), .Z(n16955) );
  AND U25435 ( .A(n16957), .B(n16958), .Z(o[236]) );
  AND U25436 ( .A(p_input[20236]), .B(p_input[10236]), .Z(n16958) );
  AND U25437 ( .A(p_input[30236]), .B(p_input[236]), .Z(n16957) );
  AND U25438 ( .A(n16959), .B(n16960), .Z(o[2369]) );
  AND U25439 ( .A(p_input[22369]), .B(p_input[12369]), .Z(n16960) );
  AND U25440 ( .A(p_input[32369]), .B(p_input[2369]), .Z(n16959) );
  AND U25441 ( .A(n16961), .B(n16962), .Z(o[2368]) );
  AND U25442 ( .A(p_input[22368]), .B(p_input[12368]), .Z(n16962) );
  AND U25443 ( .A(p_input[32368]), .B(p_input[2368]), .Z(n16961) );
  AND U25444 ( .A(n16963), .B(n16964), .Z(o[2367]) );
  AND U25445 ( .A(p_input[22367]), .B(p_input[12367]), .Z(n16964) );
  AND U25446 ( .A(p_input[32367]), .B(p_input[2367]), .Z(n16963) );
  AND U25447 ( .A(n16965), .B(n16966), .Z(o[2366]) );
  AND U25448 ( .A(p_input[22366]), .B(p_input[12366]), .Z(n16966) );
  AND U25449 ( .A(p_input[32366]), .B(p_input[2366]), .Z(n16965) );
  AND U25450 ( .A(n16967), .B(n16968), .Z(o[2365]) );
  AND U25451 ( .A(p_input[22365]), .B(p_input[12365]), .Z(n16968) );
  AND U25452 ( .A(p_input[32365]), .B(p_input[2365]), .Z(n16967) );
  AND U25453 ( .A(n16969), .B(n16970), .Z(o[2364]) );
  AND U25454 ( .A(p_input[22364]), .B(p_input[12364]), .Z(n16970) );
  AND U25455 ( .A(p_input[32364]), .B(p_input[2364]), .Z(n16969) );
  AND U25456 ( .A(n16971), .B(n16972), .Z(o[2363]) );
  AND U25457 ( .A(p_input[22363]), .B(p_input[12363]), .Z(n16972) );
  AND U25458 ( .A(p_input[32363]), .B(p_input[2363]), .Z(n16971) );
  AND U25459 ( .A(n16973), .B(n16974), .Z(o[2362]) );
  AND U25460 ( .A(p_input[22362]), .B(p_input[12362]), .Z(n16974) );
  AND U25461 ( .A(p_input[32362]), .B(p_input[2362]), .Z(n16973) );
  AND U25462 ( .A(n16975), .B(n16976), .Z(o[2361]) );
  AND U25463 ( .A(p_input[22361]), .B(p_input[12361]), .Z(n16976) );
  AND U25464 ( .A(p_input[32361]), .B(p_input[2361]), .Z(n16975) );
  AND U25465 ( .A(n16977), .B(n16978), .Z(o[2360]) );
  AND U25466 ( .A(p_input[22360]), .B(p_input[12360]), .Z(n16978) );
  AND U25467 ( .A(p_input[32360]), .B(p_input[2360]), .Z(n16977) );
  AND U25468 ( .A(n16979), .B(n16980), .Z(o[235]) );
  AND U25469 ( .A(p_input[20235]), .B(p_input[10235]), .Z(n16980) );
  AND U25470 ( .A(p_input[30235]), .B(p_input[235]), .Z(n16979) );
  AND U25471 ( .A(n16981), .B(n16982), .Z(o[2359]) );
  AND U25472 ( .A(p_input[22359]), .B(p_input[12359]), .Z(n16982) );
  AND U25473 ( .A(p_input[32359]), .B(p_input[2359]), .Z(n16981) );
  AND U25474 ( .A(n16983), .B(n16984), .Z(o[2358]) );
  AND U25475 ( .A(p_input[22358]), .B(p_input[12358]), .Z(n16984) );
  AND U25476 ( .A(p_input[32358]), .B(p_input[2358]), .Z(n16983) );
  AND U25477 ( .A(n16985), .B(n16986), .Z(o[2357]) );
  AND U25478 ( .A(p_input[22357]), .B(p_input[12357]), .Z(n16986) );
  AND U25479 ( .A(p_input[32357]), .B(p_input[2357]), .Z(n16985) );
  AND U25480 ( .A(n16987), .B(n16988), .Z(o[2356]) );
  AND U25481 ( .A(p_input[22356]), .B(p_input[12356]), .Z(n16988) );
  AND U25482 ( .A(p_input[32356]), .B(p_input[2356]), .Z(n16987) );
  AND U25483 ( .A(n16989), .B(n16990), .Z(o[2355]) );
  AND U25484 ( .A(p_input[22355]), .B(p_input[12355]), .Z(n16990) );
  AND U25485 ( .A(p_input[32355]), .B(p_input[2355]), .Z(n16989) );
  AND U25486 ( .A(n16991), .B(n16992), .Z(o[2354]) );
  AND U25487 ( .A(p_input[22354]), .B(p_input[12354]), .Z(n16992) );
  AND U25488 ( .A(p_input[32354]), .B(p_input[2354]), .Z(n16991) );
  AND U25489 ( .A(n16993), .B(n16994), .Z(o[2353]) );
  AND U25490 ( .A(p_input[22353]), .B(p_input[12353]), .Z(n16994) );
  AND U25491 ( .A(p_input[32353]), .B(p_input[2353]), .Z(n16993) );
  AND U25492 ( .A(n16995), .B(n16996), .Z(o[2352]) );
  AND U25493 ( .A(p_input[22352]), .B(p_input[12352]), .Z(n16996) );
  AND U25494 ( .A(p_input[32352]), .B(p_input[2352]), .Z(n16995) );
  AND U25495 ( .A(n16997), .B(n16998), .Z(o[2351]) );
  AND U25496 ( .A(p_input[22351]), .B(p_input[12351]), .Z(n16998) );
  AND U25497 ( .A(p_input[32351]), .B(p_input[2351]), .Z(n16997) );
  AND U25498 ( .A(n16999), .B(n17000), .Z(o[2350]) );
  AND U25499 ( .A(p_input[22350]), .B(p_input[12350]), .Z(n17000) );
  AND U25500 ( .A(p_input[32350]), .B(p_input[2350]), .Z(n16999) );
  AND U25501 ( .A(n17001), .B(n17002), .Z(o[234]) );
  AND U25502 ( .A(p_input[20234]), .B(p_input[10234]), .Z(n17002) );
  AND U25503 ( .A(p_input[30234]), .B(p_input[234]), .Z(n17001) );
  AND U25504 ( .A(n17003), .B(n17004), .Z(o[2349]) );
  AND U25505 ( .A(p_input[22349]), .B(p_input[12349]), .Z(n17004) );
  AND U25506 ( .A(p_input[32349]), .B(p_input[2349]), .Z(n17003) );
  AND U25507 ( .A(n17005), .B(n17006), .Z(o[2348]) );
  AND U25508 ( .A(p_input[22348]), .B(p_input[12348]), .Z(n17006) );
  AND U25509 ( .A(p_input[32348]), .B(p_input[2348]), .Z(n17005) );
  AND U25510 ( .A(n17007), .B(n17008), .Z(o[2347]) );
  AND U25511 ( .A(p_input[22347]), .B(p_input[12347]), .Z(n17008) );
  AND U25512 ( .A(p_input[32347]), .B(p_input[2347]), .Z(n17007) );
  AND U25513 ( .A(n17009), .B(n17010), .Z(o[2346]) );
  AND U25514 ( .A(p_input[22346]), .B(p_input[12346]), .Z(n17010) );
  AND U25515 ( .A(p_input[32346]), .B(p_input[2346]), .Z(n17009) );
  AND U25516 ( .A(n17011), .B(n17012), .Z(o[2345]) );
  AND U25517 ( .A(p_input[22345]), .B(p_input[12345]), .Z(n17012) );
  AND U25518 ( .A(p_input[32345]), .B(p_input[2345]), .Z(n17011) );
  AND U25519 ( .A(n17013), .B(n17014), .Z(o[2344]) );
  AND U25520 ( .A(p_input[22344]), .B(p_input[12344]), .Z(n17014) );
  AND U25521 ( .A(p_input[32344]), .B(p_input[2344]), .Z(n17013) );
  AND U25522 ( .A(n17015), .B(n17016), .Z(o[2343]) );
  AND U25523 ( .A(p_input[22343]), .B(p_input[12343]), .Z(n17016) );
  AND U25524 ( .A(p_input[32343]), .B(p_input[2343]), .Z(n17015) );
  AND U25525 ( .A(n17017), .B(n17018), .Z(o[2342]) );
  AND U25526 ( .A(p_input[22342]), .B(p_input[12342]), .Z(n17018) );
  AND U25527 ( .A(p_input[32342]), .B(p_input[2342]), .Z(n17017) );
  AND U25528 ( .A(n17019), .B(n17020), .Z(o[2341]) );
  AND U25529 ( .A(p_input[22341]), .B(p_input[12341]), .Z(n17020) );
  AND U25530 ( .A(p_input[32341]), .B(p_input[2341]), .Z(n17019) );
  AND U25531 ( .A(n17021), .B(n17022), .Z(o[2340]) );
  AND U25532 ( .A(p_input[22340]), .B(p_input[12340]), .Z(n17022) );
  AND U25533 ( .A(p_input[32340]), .B(p_input[2340]), .Z(n17021) );
  AND U25534 ( .A(n17023), .B(n17024), .Z(o[233]) );
  AND U25535 ( .A(p_input[20233]), .B(p_input[10233]), .Z(n17024) );
  AND U25536 ( .A(p_input[30233]), .B(p_input[233]), .Z(n17023) );
  AND U25537 ( .A(n17025), .B(n17026), .Z(o[2339]) );
  AND U25538 ( .A(p_input[22339]), .B(p_input[12339]), .Z(n17026) );
  AND U25539 ( .A(p_input[32339]), .B(p_input[2339]), .Z(n17025) );
  AND U25540 ( .A(n17027), .B(n17028), .Z(o[2338]) );
  AND U25541 ( .A(p_input[22338]), .B(p_input[12338]), .Z(n17028) );
  AND U25542 ( .A(p_input[32338]), .B(p_input[2338]), .Z(n17027) );
  AND U25543 ( .A(n17029), .B(n17030), .Z(o[2337]) );
  AND U25544 ( .A(p_input[22337]), .B(p_input[12337]), .Z(n17030) );
  AND U25545 ( .A(p_input[32337]), .B(p_input[2337]), .Z(n17029) );
  AND U25546 ( .A(n17031), .B(n17032), .Z(o[2336]) );
  AND U25547 ( .A(p_input[22336]), .B(p_input[12336]), .Z(n17032) );
  AND U25548 ( .A(p_input[32336]), .B(p_input[2336]), .Z(n17031) );
  AND U25549 ( .A(n17033), .B(n17034), .Z(o[2335]) );
  AND U25550 ( .A(p_input[22335]), .B(p_input[12335]), .Z(n17034) );
  AND U25551 ( .A(p_input[32335]), .B(p_input[2335]), .Z(n17033) );
  AND U25552 ( .A(n17035), .B(n17036), .Z(o[2334]) );
  AND U25553 ( .A(p_input[22334]), .B(p_input[12334]), .Z(n17036) );
  AND U25554 ( .A(p_input[32334]), .B(p_input[2334]), .Z(n17035) );
  AND U25555 ( .A(n17037), .B(n17038), .Z(o[2333]) );
  AND U25556 ( .A(p_input[22333]), .B(p_input[12333]), .Z(n17038) );
  AND U25557 ( .A(p_input[32333]), .B(p_input[2333]), .Z(n17037) );
  AND U25558 ( .A(n17039), .B(n17040), .Z(o[2332]) );
  AND U25559 ( .A(p_input[22332]), .B(p_input[12332]), .Z(n17040) );
  AND U25560 ( .A(p_input[32332]), .B(p_input[2332]), .Z(n17039) );
  AND U25561 ( .A(n17041), .B(n17042), .Z(o[2331]) );
  AND U25562 ( .A(p_input[22331]), .B(p_input[12331]), .Z(n17042) );
  AND U25563 ( .A(p_input[32331]), .B(p_input[2331]), .Z(n17041) );
  AND U25564 ( .A(n17043), .B(n17044), .Z(o[2330]) );
  AND U25565 ( .A(p_input[22330]), .B(p_input[12330]), .Z(n17044) );
  AND U25566 ( .A(p_input[32330]), .B(p_input[2330]), .Z(n17043) );
  AND U25567 ( .A(n17045), .B(n17046), .Z(o[232]) );
  AND U25568 ( .A(p_input[20232]), .B(p_input[10232]), .Z(n17046) );
  AND U25569 ( .A(p_input[30232]), .B(p_input[232]), .Z(n17045) );
  AND U25570 ( .A(n17047), .B(n17048), .Z(o[2329]) );
  AND U25571 ( .A(p_input[22329]), .B(p_input[12329]), .Z(n17048) );
  AND U25572 ( .A(p_input[32329]), .B(p_input[2329]), .Z(n17047) );
  AND U25573 ( .A(n17049), .B(n17050), .Z(o[2328]) );
  AND U25574 ( .A(p_input[22328]), .B(p_input[12328]), .Z(n17050) );
  AND U25575 ( .A(p_input[32328]), .B(p_input[2328]), .Z(n17049) );
  AND U25576 ( .A(n17051), .B(n17052), .Z(o[2327]) );
  AND U25577 ( .A(p_input[22327]), .B(p_input[12327]), .Z(n17052) );
  AND U25578 ( .A(p_input[32327]), .B(p_input[2327]), .Z(n17051) );
  AND U25579 ( .A(n17053), .B(n17054), .Z(o[2326]) );
  AND U25580 ( .A(p_input[22326]), .B(p_input[12326]), .Z(n17054) );
  AND U25581 ( .A(p_input[32326]), .B(p_input[2326]), .Z(n17053) );
  AND U25582 ( .A(n17055), .B(n17056), .Z(o[2325]) );
  AND U25583 ( .A(p_input[22325]), .B(p_input[12325]), .Z(n17056) );
  AND U25584 ( .A(p_input[32325]), .B(p_input[2325]), .Z(n17055) );
  AND U25585 ( .A(n17057), .B(n17058), .Z(o[2324]) );
  AND U25586 ( .A(p_input[22324]), .B(p_input[12324]), .Z(n17058) );
  AND U25587 ( .A(p_input[32324]), .B(p_input[2324]), .Z(n17057) );
  AND U25588 ( .A(n17059), .B(n17060), .Z(o[2323]) );
  AND U25589 ( .A(p_input[22323]), .B(p_input[12323]), .Z(n17060) );
  AND U25590 ( .A(p_input[32323]), .B(p_input[2323]), .Z(n17059) );
  AND U25591 ( .A(n17061), .B(n17062), .Z(o[2322]) );
  AND U25592 ( .A(p_input[22322]), .B(p_input[12322]), .Z(n17062) );
  AND U25593 ( .A(p_input[32322]), .B(p_input[2322]), .Z(n17061) );
  AND U25594 ( .A(n17063), .B(n17064), .Z(o[2321]) );
  AND U25595 ( .A(p_input[22321]), .B(p_input[12321]), .Z(n17064) );
  AND U25596 ( .A(p_input[32321]), .B(p_input[2321]), .Z(n17063) );
  AND U25597 ( .A(n17065), .B(n17066), .Z(o[2320]) );
  AND U25598 ( .A(p_input[22320]), .B(p_input[12320]), .Z(n17066) );
  AND U25599 ( .A(p_input[32320]), .B(p_input[2320]), .Z(n17065) );
  AND U25600 ( .A(n17067), .B(n17068), .Z(o[231]) );
  AND U25601 ( .A(p_input[20231]), .B(p_input[10231]), .Z(n17068) );
  AND U25602 ( .A(p_input[30231]), .B(p_input[231]), .Z(n17067) );
  AND U25603 ( .A(n17069), .B(n17070), .Z(o[2319]) );
  AND U25604 ( .A(p_input[22319]), .B(p_input[12319]), .Z(n17070) );
  AND U25605 ( .A(p_input[32319]), .B(p_input[2319]), .Z(n17069) );
  AND U25606 ( .A(n17071), .B(n17072), .Z(o[2318]) );
  AND U25607 ( .A(p_input[22318]), .B(p_input[12318]), .Z(n17072) );
  AND U25608 ( .A(p_input[32318]), .B(p_input[2318]), .Z(n17071) );
  AND U25609 ( .A(n17073), .B(n17074), .Z(o[2317]) );
  AND U25610 ( .A(p_input[22317]), .B(p_input[12317]), .Z(n17074) );
  AND U25611 ( .A(p_input[32317]), .B(p_input[2317]), .Z(n17073) );
  AND U25612 ( .A(n17075), .B(n17076), .Z(o[2316]) );
  AND U25613 ( .A(p_input[22316]), .B(p_input[12316]), .Z(n17076) );
  AND U25614 ( .A(p_input[32316]), .B(p_input[2316]), .Z(n17075) );
  AND U25615 ( .A(n17077), .B(n17078), .Z(o[2315]) );
  AND U25616 ( .A(p_input[22315]), .B(p_input[12315]), .Z(n17078) );
  AND U25617 ( .A(p_input[32315]), .B(p_input[2315]), .Z(n17077) );
  AND U25618 ( .A(n17079), .B(n17080), .Z(o[2314]) );
  AND U25619 ( .A(p_input[22314]), .B(p_input[12314]), .Z(n17080) );
  AND U25620 ( .A(p_input[32314]), .B(p_input[2314]), .Z(n17079) );
  AND U25621 ( .A(n17081), .B(n17082), .Z(o[2313]) );
  AND U25622 ( .A(p_input[22313]), .B(p_input[12313]), .Z(n17082) );
  AND U25623 ( .A(p_input[32313]), .B(p_input[2313]), .Z(n17081) );
  AND U25624 ( .A(n17083), .B(n17084), .Z(o[2312]) );
  AND U25625 ( .A(p_input[22312]), .B(p_input[12312]), .Z(n17084) );
  AND U25626 ( .A(p_input[32312]), .B(p_input[2312]), .Z(n17083) );
  AND U25627 ( .A(n17085), .B(n17086), .Z(o[2311]) );
  AND U25628 ( .A(p_input[22311]), .B(p_input[12311]), .Z(n17086) );
  AND U25629 ( .A(p_input[32311]), .B(p_input[2311]), .Z(n17085) );
  AND U25630 ( .A(n17087), .B(n17088), .Z(o[2310]) );
  AND U25631 ( .A(p_input[22310]), .B(p_input[12310]), .Z(n17088) );
  AND U25632 ( .A(p_input[32310]), .B(p_input[2310]), .Z(n17087) );
  AND U25633 ( .A(n17089), .B(n17090), .Z(o[230]) );
  AND U25634 ( .A(p_input[20230]), .B(p_input[10230]), .Z(n17090) );
  AND U25635 ( .A(p_input[30230]), .B(p_input[230]), .Z(n17089) );
  AND U25636 ( .A(n17091), .B(n17092), .Z(o[2309]) );
  AND U25637 ( .A(p_input[22309]), .B(p_input[12309]), .Z(n17092) );
  AND U25638 ( .A(p_input[32309]), .B(p_input[2309]), .Z(n17091) );
  AND U25639 ( .A(n17093), .B(n17094), .Z(o[2308]) );
  AND U25640 ( .A(p_input[22308]), .B(p_input[12308]), .Z(n17094) );
  AND U25641 ( .A(p_input[32308]), .B(p_input[2308]), .Z(n17093) );
  AND U25642 ( .A(n17095), .B(n17096), .Z(o[2307]) );
  AND U25643 ( .A(p_input[22307]), .B(p_input[12307]), .Z(n17096) );
  AND U25644 ( .A(p_input[32307]), .B(p_input[2307]), .Z(n17095) );
  AND U25645 ( .A(n17097), .B(n17098), .Z(o[2306]) );
  AND U25646 ( .A(p_input[22306]), .B(p_input[12306]), .Z(n17098) );
  AND U25647 ( .A(p_input[32306]), .B(p_input[2306]), .Z(n17097) );
  AND U25648 ( .A(n17099), .B(n17100), .Z(o[2305]) );
  AND U25649 ( .A(p_input[22305]), .B(p_input[12305]), .Z(n17100) );
  AND U25650 ( .A(p_input[32305]), .B(p_input[2305]), .Z(n17099) );
  AND U25651 ( .A(n17101), .B(n17102), .Z(o[2304]) );
  AND U25652 ( .A(p_input[22304]), .B(p_input[12304]), .Z(n17102) );
  AND U25653 ( .A(p_input[32304]), .B(p_input[2304]), .Z(n17101) );
  AND U25654 ( .A(n17103), .B(n17104), .Z(o[2303]) );
  AND U25655 ( .A(p_input[22303]), .B(p_input[12303]), .Z(n17104) );
  AND U25656 ( .A(p_input[32303]), .B(p_input[2303]), .Z(n17103) );
  AND U25657 ( .A(n17105), .B(n17106), .Z(o[2302]) );
  AND U25658 ( .A(p_input[22302]), .B(p_input[12302]), .Z(n17106) );
  AND U25659 ( .A(p_input[32302]), .B(p_input[2302]), .Z(n17105) );
  AND U25660 ( .A(n17107), .B(n17108), .Z(o[2301]) );
  AND U25661 ( .A(p_input[22301]), .B(p_input[12301]), .Z(n17108) );
  AND U25662 ( .A(p_input[32301]), .B(p_input[2301]), .Z(n17107) );
  AND U25663 ( .A(n17109), .B(n17110), .Z(o[2300]) );
  AND U25664 ( .A(p_input[22300]), .B(p_input[12300]), .Z(n17110) );
  AND U25665 ( .A(p_input[32300]), .B(p_input[2300]), .Z(n17109) );
  AND U25666 ( .A(n17111), .B(n17112), .Z(o[22]) );
  AND U25667 ( .A(p_input[20022]), .B(p_input[10022]), .Z(n17112) );
  AND U25668 ( .A(p_input[30022]), .B(p_input[22]), .Z(n17111) );
  AND U25669 ( .A(n17113), .B(n17114), .Z(o[229]) );
  AND U25670 ( .A(p_input[20229]), .B(p_input[10229]), .Z(n17114) );
  AND U25671 ( .A(p_input[30229]), .B(p_input[229]), .Z(n17113) );
  AND U25672 ( .A(n17115), .B(n17116), .Z(o[2299]) );
  AND U25673 ( .A(p_input[22299]), .B(p_input[12299]), .Z(n17116) );
  AND U25674 ( .A(p_input[32299]), .B(p_input[2299]), .Z(n17115) );
  AND U25675 ( .A(n17117), .B(n17118), .Z(o[2298]) );
  AND U25676 ( .A(p_input[22298]), .B(p_input[12298]), .Z(n17118) );
  AND U25677 ( .A(p_input[32298]), .B(p_input[2298]), .Z(n17117) );
  AND U25678 ( .A(n17119), .B(n17120), .Z(o[2297]) );
  AND U25679 ( .A(p_input[22297]), .B(p_input[12297]), .Z(n17120) );
  AND U25680 ( .A(p_input[32297]), .B(p_input[2297]), .Z(n17119) );
  AND U25681 ( .A(n17121), .B(n17122), .Z(o[2296]) );
  AND U25682 ( .A(p_input[22296]), .B(p_input[12296]), .Z(n17122) );
  AND U25683 ( .A(p_input[32296]), .B(p_input[2296]), .Z(n17121) );
  AND U25684 ( .A(n17123), .B(n17124), .Z(o[2295]) );
  AND U25685 ( .A(p_input[22295]), .B(p_input[12295]), .Z(n17124) );
  AND U25686 ( .A(p_input[32295]), .B(p_input[2295]), .Z(n17123) );
  AND U25687 ( .A(n17125), .B(n17126), .Z(o[2294]) );
  AND U25688 ( .A(p_input[22294]), .B(p_input[12294]), .Z(n17126) );
  AND U25689 ( .A(p_input[32294]), .B(p_input[2294]), .Z(n17125) );
  AND U25690 ( .A(n17127), .B(n17128), .Z(o[2293]) );
  AND U25691 ( .A(p_input[22293]), .B(p_input[12293]), .Z(n17128) );
  AND U25692 ( .A(p_input[32293]), .B(p_input[2293]), .Z(n17127) );
  AND U25693 ( .A(n17129), .B(n17130), .Z(o[2292]) );
  AND U25694 ( .A(p_input[22292]), .B(p_input[12292]), .Z(n17130) );
  AND U25695 ( .A(p_input[32292]), .B(p_input[2292]), .Z(n17129) );
  AND U25696 ( .A(n17131), .B(n17132), .Z(o[2291]) );
  AND U25697 ( .A(p_input[22291]), .B(p_input[12291]), .Z(n17132) );
  AND U25698 ( .A(p_input[32291]), .B(p_input[2291]), .Z(n17131) );
  AND U25699 ( .A(n17133), .B(n17134), .Z(o[2290]) );
  AND U25700 ( .A(p_input[22290]), .B(p_input[12290]), .Z(n17134) );
  AND U25701 ( .A(p_input[32290]), .B(p_input[2290]), .Z(n17133) );
  AND U25702 ( .A(n17135), .B(n17136), .Z(o[228]) );
  AND U25703 ( .A(p_input[20228]), .B(p_input[10228]), .Z(n17136) );
  AND U25704 ( .A(p_input[30228]), .B(p_input[228]), .Z(n17135) );
  AND U25705 ( .A(n17137), .B(n17138), .Z(o[2289]) );
  AND U25706 ( .A(p_input[22289]), .B(p_input[12289]), .Z(n17138) );
  AND U25707 ( .A(p_input[32289]), .B(p_input[2289]), .Z(n17137) );
  AND U25708 ( .A(n17139), .B(n17140), .Z(o[2288]) );
  AND U25709 ( .A(p_input[22288]), .B(p_input[12288]), .Z(n17140) );
  AND U25710 ( .A(p_input[32288]), .B(p_input[2288]), .Z(n17139) );
  AND U25711 ( .A(n17141), .B(n17142), .Z(o[2287]) );
  AND U25712 ( .A(p_input[22287]), .B(p_input[12287]), .Z(n17142) );
  AND U25713 ( .A(p_input[32287]), .B(p_input[2287]), .Z(n17141) );
  AND U25714 ( .A(n17143), .B(n17144), .Z(o[2286]) );
  AND U25715 ( .A(p_input[22286]), .B(p_input[12286]), .Z(n17144) );
  AND U25716 ( .A(p_input[32286]), .B(p_input[2286]), .Z(n17143) );
  AND U25717 ( .A(n17145), .B(n17146), .Z(o[2285]) );
  AND U25718 ( .A(p_input[22285]), .B(p_input[12285]), .Z(n17146) );
  AND U25719 ( .A(p_input[32285]), .B(p_input[2285]), .Z(n17145) );
  AND U25720 ( .A(n17147), .B(n17148), .Z(o[2284]) );
  AND U25721 ( .A(p_input[22284]), .B(p_input[12284]), .Z(n17148) );
  AND U25722 ( .A(p_input[32284]), .B(p_input[2284]), .Z(n17147) );
  AND U25723 ( .A(n17149), .B(n17150), .Z(o[2283]) );
  AND U25724 ( .A(p_input[22283]), .B(p_input[12283]), .Z(n17150) );
  AND U25725 ( .A(p_input[32283]), .B(p_input[2283]), .Z(n17149) );
  AND U25726 ( .A(n17151), .B(n17152), .Z(o[2282]) );
  AND U25727 ( .A(p_input[22282]), .B(p_input[12282]), .Z(n17152) );
  AND U25728 ( .A(p_input[32282]), .B(p_input[2282]), .Z(n17151) );
  AND U25729 ( .A(n17153), .B(n17154), .Z(o[2281]) );
  AND U25730 ( .A(p_input[22281]), .B(p_input[12281]), .Z(n17154) );
  AND U25731 ( .A(p_input[32281]), .B(p_input[2281]), .Z(n17153) );
  AND U25732 ( .A(n17155), .B(n17156), .Z(o[2280]) );
  AND U25733 ( .A(p_input[22280]), .B(p_input[12280]), .Z(n17156) );
  AND U25734 ( .A(p_input[32280]), .B(p_input[2280]), .Z(n17155) );
  AND U25735 ( .A(n17157), .B(n17158), .Z(o[227]) );
  AND U25736 ( .A(p_input[20227]), .B(p_input[10227]), .Z(n17158) );
  AND U25737 ( .A(p_input[30227]), .B(p_input[227]), .Z(n17157) );
  AND U25738 ( .A(n17159), .B(n17160), .Z(o[2279]) );
  AND U25739 ( .A(p_input[22279]), .B(p_input[12279]), .Z(n17160) );
  AND U25740 ( .A(p_input[32279]), .B(p_input[2279]), .Z(n17159) );
  AND U25741 ( .A(n17161), .B(n17162), .Z(o[2278]) );
  AND U25742 ( .A(p_input[22278]), .B(p_input[12278]), .Z(n17162) );
  AND U25743 ( .A(p_input[32278]), .B(p_input[2278]), .Z(n17161) );
  AND U25744 ( .A(n17163), .B(n17164), .Z(o[2277]) );
  AND U25745 ( .A(p_input[22277]), .B(p_input[12277]), .Z(n17164) );
  AND U25746 ( .A(p_input[32277]), .B(p_input[2277]), .Z(n17163) );
  AND U25747 ( .A(n17165), .B(n17166), .Z(o[2276]) );
  AND U25748 ( .A(p_input[22276]), .B(p_input[12276]), .Z(n17166) );
  AND U25749 ( .A(p_input[32276]), .B(p_input[2276]), .Z(n17165) );
  AND U25750 ( .A(n17167), .B(n17168), .Z(o[2275]) );
  AND U25751 ( .A(p_input[22275]), .B(p_input[12275]), .Z(n17168) );
  AND U25752 ( .A(p_input[32275]), .B(p_input[2275]), .Z(n17167) );
  AND U25753 ( .A(n17169), .B(n17170), .Z(o[2274]) );
  AND U25754 ( .A(p_input[22274]), .B(p_input[12274]), .Z(n17170) );
  AND U25755 ( .A(p_input[32274]), .B(p_input[2274]), .Z(n17169) );
  AND U25756 ( .A(n17171), .B(n17172), .Z(o[2273]) );
  AND U25757 ( .A(p_input[22273]), .B(p_input[12273]), .Z(n17172) );
  AND U25758 ( .A(p_input[32273]), .B(p_input[2273]), .Z(n17171) );
  AND U25759 ( .A(n17173), .B(n17174), .Z(o[2272]) );
  AND U25760 ( .A(p_input[22272]), .B(p_input[12272]), .Z(n17174) );
  AND U25761 ( .A(p_input[32272]), .B(p_input[2272]), .Z(n17173) );
  AND U25762 ( .A(n17175), .B(n17176), .Z(o[2271]) );
  AND U25763 ( .A(p_input[22271]), .B(p_input[12271]), .Z(n17176) );
  AND U25764 ( .A(p_input[32271]), .B(p_input[2271]), .Z(n17175) );
  AND U25765 ( .A(n17177), .B(n17178), .Z(o[2270]) );
  AND U25766 ( .A(p_input[22270]), .B(p_input[12270]), .Z(n17178) );
  AND U25767 ( .A(p_input[32270]), .B(p_input[2270]), .Z(n17177) );
  AND U25768 ( .A(n17179), .B(n17180), .Z(o[226]) );
  AND U25769 ( .A(p_input[20226]), .B(p_input[10226]), .Z(n17180) );
  AND U25770 ( .A(p_input[30226]), .B(p_input[226]), .Z(n17179) );
  AND U25771 ( .A(n17181), .B(n17182), .Z(o[2269]) );
  AND U25772 ( .A(p_input[22269]), .B(p_input[12269]), .Z(n17182) );
  AND U25773 ( .A(p_input[32269]), .B(p_input[2269]), .Z(n17181) );
  AND U25774 ( .A(n17183), .B(n17184), .Z(o[2268]) );
  AND U25775 ( .A(p_input[22268]), .B(p_input[12268]), .Z(n17184) );
  AND U25776 ( .A(p_input[32268]), .B(p_input[2268]), .Z(n17183) );
  AND U25777 ( .A(n17185), .B(n17186), .Z(o[2267]) );
  AND U25778 ( .A(p_input[22267]), .B(p_input[12267]), .Z(n17186) );
  AND U25779 ( .A(p_input[32267]), .B(p_input[2267]), .Z(n17185) );
  AND U25780 ( .A(n17187), .B(n17188), .Z(o[2266]) );
  AND U25781 ( .A(p_input[22266]), .B(p_input[12266]), .Z(n17188) );
  AND U25782 ( .A(p_input[32266]), .B(p_input[2266]), .Z(n17187) );
  AND U25783 ( .A(n17189), .B(n17190), .Z(o[2265]) );
  AND U25784 ( .A(p_input[22265]), .B(p_input[12265]), .Z(n17190) );
  AND U25785 ( .A(p_input[32265]), .B(p_input[2265]), .Z(n17189) );
  AND U25786 ( .A(n17191), .B(n17192), .Z(o[2264]) );
  AND U25787 ( .A(p_input[22264]), .B(p_input[12264]), .Z(n17192) );
  AND U25788 ( .A(p_input[32264]), .B(p_input[2264]), .Z(n17191) );
  AND U25789 ( .A(n17193), .B(n17194), .Z(o[2263]) );
  AND U25790 ( .A(p_input[22263]), .B(p_input[12263]), .Z(n17194) );
  AND U25791 ( .A(p_input[32263]), .B(p_input[2263]), .Z(n17193) );
  AND U25792 ( .A(n17195), .B(n17196), .Z(o[2262]) );
  AND U25793 ( .A(p_input[22262]), .B(p_input[12262]), .Z(n17196) );
  AND U25794 ( .A(p_input[32262]), .B(p_input[2262]), .Z(n17195) );
  AND U25795 ( .A(n17197), .B(n17198), .Z(o[2261]) );
  AND U25796 ( .A(p_input[22261]), .B(p_input[12261]), .Z(n17198) );
  AND U25797 ( .A(p_input[32261]), .B(p_input[2261]), .Z(n17197) );
  AND U25798 ( .A(n17199), .B(n17200), .Z(o[2260]) );
  AND U25799 ( .A(p_input[22260]), .B(p_input[12260]), .Z(n17200) );
  AND U25800 ( .A(p_input[32260]), .B(p_input[2260]), .Z(n17199) );
  AND U25801 ( .A(n17201), .B(n17202), .Z(o[225]) );
  AND U25802 ( .A(p_input[20225]), .B(p_input[10225]), .Z(n17202) );
  AND U25803 ( .A(p_input[30225]), .B(p_input[225]), .Z(n17201) );
  AND U25804 ( .A(n17203), .B(n17204), .Z(o[2259]) );
  AND U25805 ( .A(p_input[22259]), .B(p_input[12259]), .Z(n17204) );
  AND U25806 ( .A(p_input[32259]), .B(p_input[2259]), .Z(n17203) );
  AND U25807 ( .A(n17205), .B(n17206), .Z(o[2258]) );
  AND U25808 ( .A(p_input[22258]), .B(p_input[12258]), .Z(n17206) );
  AND U25809 ( .A(p_input[32258]), .B(p_input[2258]), .Z(n17205) );
  AND U25810 ( .A(n17207), .B(n17208), .Z(o[2257]) );
  AND U25811 ( .A(p_input[22257]), .B(p_input[12257]), .Z(n17208) );
  AND U25812 ( .A(p_input[32257]), .B(p_input[2257]), .Z(n17207) );
  AND U25813 ( .A(n17209), .B(n17210), .Z(o[2256]) );
  AND U25814 ( .A(p_input[22256]), .B(p_input[12256]), .Z(n17210) );
  AND U25815 ( .A(p_input[32256]), .B(p_input[2256]), .Z(n17209) );
  AND U25816 ( .A(n17211), .B(n17212), .Z(o[2255]) );
  AND U25817 ( .A(p_input[22255]), .B(p_input[12255]), .Z(n17212) );
  AND U25818 ( .A(p_input[32255]), .B(p_input[2255]), .Z(n17211) );
  AND U25819 ( .A(n17213), .B(n17214), .Z(o[2254]) );
  AND U25820 ( .A(p_input[22254]), .B(p_input[12254]), .Z(n17214) );
  AND U25821 ( .A(p_input[32254]), .B(p_input[2254]), .Z(n17213) );
  AND U25822 ( .A(n17215), .B(n17216), .Z(o[2253]) );
  AND U25823 ( .A(p_input[22253]), .B(p_input[12253]), .Z(n17216) );
  AND U25824 ( .A(p_input[32253]), .B(p_input[2253]), .Z(n17215) );
  AND U25825 ( .A(n17217), .B(n17218), .Z(o[2252]) );
  AND U25826 ( .A(p_input[22252]), .B(p_input[12252]), .Z(n17218) );
  AND U25827 ( .A(p_input[32252]), .B(p_input[2252]), .Z(n17217) );
  AND U25828 ( .A(n17219), .B(n17220), .Z(o[2251]) );
  AND U25829 ( .A(p_input[22251]), .B(p_input[12251]), .Z(n17220) );
  AND U25830 ( .A(p_input[32251]), .B(p_input[2251]), .Z(n17219) );
  AND U25831 ( .A(n17221), .B(n17222), .Z(o[2250]) );
  AND U25832 ( .A(p_input[22250]), .B(p_input[12250]), .Z(n17222) );
  AND U25833 ( .A(p_input[32250]), .B(p_input[2250]), .Z(n17221) );
  AND U25834 ( .A(n17223), .B(n17224), .Z(o[224]) );
  AND U25835 ( .A(p_input[20224]), .B(p_input[10224]), .Z(n17224) );
  AND U25836 ( .A(p_input[30224]), .B(p_input[224]), .Z(n17223) );
  AND U25837 ( .A(n17225), .B(n17226), .Z(o[2249]) );
  AND U25838 ( .A(p_input[22249]), .B(p_input[12249]), .Z(n17226) );
  AND U25839 ( .A(p_input[32249]), .B(p_input[2249]), .Z(n17225) );
  AND U25840 ( .A(n17227), .B(n17228), .Z(o[2248]) );
  AND U25841 ( .A(p_input[22248]), .B(p_input[12248]), .Z(n17228) );
  AND U25842 ( .A(p_input[32248]), .B(p_input[2248]), .Z(n17227) );
  AND U25843 ( .A(n17229), .B(n17230), .Z(o[2247]) );
  AND U25844 ( .A(p_input[22247]), .B(p_input[12247]), .Z(n17230) );
  AND U25845 ( .A(p_input[32247]), .B(p_input[2247]), .Z(n17229) );
  AND U25846 ( .A(n17231), .B(n17232), .Z(o[2246]) );
  AND U25847 ( .A(p_input[22246]), .B(p_input[12246]), .Z(n17232) );
  AND U25848 ( .A(p_input[32246]), .B(p_input[2246]), .Z(n17231) );
  AND U25849 ( .A(n17233), .B(n17234), .Z(o[2245]) );
  AND U25850 ( .A(p_input[22245]), .B(p_input[12245]), .Z(n17234) );
  AND U25851 ( .A(p_input[32245]), .B(p_input[2245]), .Z(n17233) );
  AND U25852 ( .A(n17235), .B(n17236), .Z(o[2244]) );
  AND U25853 ( .A(p_input[22244]), .B(p_input[12244]), .Z(n17236) );
  AND U25854 ( .A(p_input[32244]), .B(p_input[2244]), .Z(n17235) );
  AND U25855 ( .A(n17237), .B(n17238), .Z(o[2243]) );
  AND U25856 ( .A(p_input[22243]), .B(p_input[12243]), .Z(n17238) );
  AND U25857 ( .A(p_input[32243]), .B(p_input[2243]), .Z(n17237) );
  AND U25858 ( .A(n17239), .B(n17240), .Z(o[2242]) );
  AND U25859 ( .A(p_input[22242]), .B(p_input[12242]), .Z(n17240) );
  AND U25860 ( .A(p_input[32242]), .B(p_input[2242]), .Z(n17239) );
  AND U25861 ( .A(n17241), .B(n17242), .Z(o[2241]) );
  AND U25862 ( .A(p_input[22241]), .B(p_input[12241]), .Z(n17242) );
  AND U25863 ( .A(p_input[32241]), .B(p_input[2241]), .Z(n17241) );
  AND U25864 ( .A(n17243), .B(n17244), .Z(o[2240]) );
  AND U25865 ( .A(p_input[22240]), .B(p_input[12240]), .Z(n17244) );
  AND U25866 ( .A(p_input[32240]), .B(p_input[2240]), .Z(n17243) );
  AND U25867 ( .A(n17245), .B(n17246), .Z(o[223]) );
  AND U25868 ( .A(p_input[20223]), .B(p_input[10223]), .Z(n17246) );
  AND U25869 ( .A(p_input[30223]), .B(p_input[223]), .Z(n17245) );
  AND U25870 ( .A(n17247), .B(n17248), .Z(o[2239]) );
  AND U25871 ( .A(p_input[22239]), .B(p_input[12239]), .Z(n17248) );
  AND U25872 ( .A(p_input[32239]), .B(p_input[2239]), .Z(n17247) );
  AND U25873 ( .A(n17249), .B(n17250), .Z(o[2238]) );
  AND U25874 ( .A(p_input[22238]), .B(p_input[12238]), .Z(n17250) );
  AND U25875 ( .A(p_input[32238]), .B(p_input[2238]), .Z(n17249) );
  AND U25876 ( .A(n17251), .B(n17252), .Z(o[2237]) );
  AND U25877 ( .A(p_input[22237]), .B(p_input[12237]), .Z(n17252) );
  AND U25878 ( .A(p_input[32237]), .B(p_input[2237]), .Z(n17251) );
  AND U25879 ( .A(n17253), .B(n17254), .Z(o[2236]) );
  AND U25880 ( .A(p_input[22236]), .B(p_input[12236]), .Z(n17254) );
  AND U25881 ( .A(p_input[32236]), .B(p_input[2236]), .Z(n17253) );
  AND U25882 ( .A(n17255), .B(n17256), .Z(o[2235]) );
  AND U25883 ( .A(p_input[22235]), .B(p_input[12235]), .Z(n17256) );
  AND U25884 ( .A(p_input[32235]), .B(p_input[2235]), .Z(n17255) );
  AND U25885 ( .A(n17257), .B(n17258), .Z(o[2234]) );
  AND U25886 ( .A(p_input[22234]), .B(p_input[12234]), .Z(n17258) );
  AND U25887 ( .A(p_input[32234]), .B(p_input[2234]), .Z(n17257) );
  AND U25888 ( .A(n17259), .B(n17260), .Z(o[2233]) );
  AND U25889 ( .A(p_input[22233]), .B(p_input[12233]), .Z(n17260) );
  AND U25890 ( .A(p_input[32233]), .B(p_input[2233]), .Z(n17259) );
  AND U25891 ( .A(n17261), .B(n17262), .Z(o[2232]) );
  AND U25892 ( .A(p_input[22232]), .B(p_input[12232]), .Z(n17262) );
  AND U25893 ( .A(p_input[32232]), .B(p_input[2232]), .Z(n17261) );
  AND U25894 ( .A(n17263), .B(n17264), .Z(o[2231]) );
  AND U25895 ( .A(p_input[22231]), .B(p_input[12231]), .Z(n17264) );
  AND U25896 ( .A(p_input[32231]), .B(p_input[2231]), .Z(n17263) );
  AND U25897 ( .A(n17265), .B(n17266), .Z(o[2230]) );
  AND U25898 ( .A(p_input[22230]), .B(p_input[12230]), .Z(n17266) );
  AND U25899 ( .A(p_input[32230]), .B(p_input[2230]), .Z(n17265) );
  AND U25900 ( .A(n17267), .B(n17268), .Z(o[222]) );
  AND U25901 ( .A(p_input[20222]), .B(p_input[10222]), .Z(n17268) );
  AND U25902 ( .A(p_input[30222]), .B(p_input[222]), .Z(n17267) );
  AND U25903 ( .A(n17269), .B(n17270), .Z(o[2229]) );
  AND U25904 ( .A(p_input[22229]), .B(p_input[12229]), .Z(n17270) );
  AND U25905 ( .A(p_input[32229]), .B(p_input[2229]), .Z(n17269) );
  AND U25906 ( .A(n17271), .B(n17272), .Z(o[2228]) );
  AND U25907 ( .A(p_input[22228]), .B(p_input[12228]), .Z(n17272) );
  AND U25908 ( .A(p_input[32228]), .B(p_input[2228]), .Z(n17271) );
  AND U25909 ( .A(n17273), .B(n17274), .Z(o[2227]) );
  AND U25910 ( .A(p_input[22227]), .B(p_input[12227]), .Z(n17274) );
  AND U25911 ( .A(p_input[32227]), .B(p_input[2227]), .Z(n17273) );
  AND U25912 ( .A(n17275), .B(n17276), .Z(o[2226]) );
  AND U25913 ( .A(p_input[22226]), .B(p_input[12226]), .Z(n17276) );
  AND U25914 ( .A(p_input[32226]), .B(p_input[2226]), .Z(n17275) );
  AND U25915 ( .A(n17277), .B(n17278), .Z(o[2225]) );
  AND U25916 ( .A(p_input[22225]), .B(p_input[12225]), .Z(n17278) );
  AND U25917 ( .A(p_input[32225]), .B(p_input[2225]), .Z(n17277) );
  AND U25918 ( .A(n17279), .B(n17280), .Z(o[2224]) );
  AND U25919 ( .A(p_input[22224]), .B(p_input[12224]), .Z(n17280) );
  AND U25920 ( .A(p_input[32224]), .B(p_input[2224]), .Z(n17279) );
  AND U25921 ( .A(n17281), .B(n17282), .Z(o[2223]) );
  AND U25922 ( .A(p_input[22223]), .B(p_input[12223]), .Z(n17282) );
  AND U25923 ( .A(p_input[32223]), .B(p_input[2223]), .Z(n17281) );
  AND U25924 ( .A(n17283), .B(n17284), .Z(o[2222]) );
  AND U25925 ( .A(p_input[22222]), .B(p_input[12222]), .Z(n17284) );
  AND U25926 ( .A(p_input[32222]), .B(p_input[2222]), .Z(n17283) );
  AND U25927 ( .A(n17285), .B(n17286), .Z(o[2221]) );
  AND U25928 ( .A(p_input[2221]), .B(p_input[12221]), .Z(n17286) );
  AND U25929 ( .A(p_input[32221]), .B(p_input[22221]), .Z(n17285) );
  AND U25930 ( .A(n17287), .B(n17288), .Z(o[2220]) );
  AND U25931 ( .A(p_input[2220]), .B(p_input[12220]), .Z(n17288) );
  AND U25932 ( .A(p_input[32220]), .B(p_input[22220]), .Z(n17287) );
  AND U25933 ( .A(n17289), .B(n17290), .Z(o[221]) );
  AND U25934 ( .A(p_input[20221]), .B(p_input[10221]), .Z(n17290) );
  AND U25935 ( .A(p_input[30221]), .B(p_input[221]), .Z(n17289) );
  AND U25936 ( .A(n17291), .B(n17292), .Z(o[2219]) );
  AND U25937 ( .A(p_input[2219]), .B(p_input[12219]), .Z(n17292) );
  AND U25938 ( .A(p_input[32219]), .B(p_input[22219]), .Z(n17291) );
  AND U25939 ( .A(n17293), .B(n17294), .Z(o[2218]) );
  AND U25940 ( .A(p_input[2218]), .B(p_input[12218]), .Z(n17294) );
  AND U25941 ( .A(p_input[32218]), .B(p_input[22218]), .Z(n17293) );
  AND U25942 ( .A(n17295), .B(n17296), .Z(o[2217]) );
  AND U25943 ( .A(p_input[2217]), .B(p_input[12217]), .Z(n17296) );
  AND U25944 ( .A(p_input[32217]), .B(p_input[22217]), .Z(n17295) );
  AND U25945 ( .A(n17297), .B(n17298), .Z(o[2216]) );
  AND U25946 ( .A(p_input[2216]), .B(p_input[12216]), .Z(n17298) );
  AND U25947 ( .A(p_input[32216]), .B(p_input[22216]), .Z(n17297) );
  AND U25948 ( .A(n17299), .B(n17300), .Z(o[2215]) );
  AND U25949 ( .A(p_input[2215]), .B(p_input[12215]), .Z(n17300) );
  AND U25950 ( .A(p_input[32215]), .B(p_input[22215]), .Z(n17299) );
  AND U25951 ( .A(n17301), .B(n17302), .Z(o[2214]) );
  AND U25952 ( .A(p_input[2214]), .B(p_input[12214]), .Z(n17302) );
  AND U25953 ( .A(p_input[32214]), .B(p_input[22214]), .Z(n17301) );
  AND U25954 ( .A(n17303), .B(n17304), .Z(o[2213]) );
  AND U25955 ( .A(p_input[2213]), .B(p_input[12213]), .Z(n17304) );
  AND U25956 ( .A(p_input[32213]), .B(p_input[22213]), .Z(n17303) );
  AND U25957 ( .A(n17305), .B(n17306), .Z(o[2212]) );
  AND U25958 ( .A(p_input[2212]), .B(p_input[12212]), .Z(n17306) );
  AND U25959 ( .A(p_input[32212]), .B(p_input[22212]), .Z(n17305) );
  AND U25960 ( .A(n17307), .B(n17308), .Z(o[2211]) );
  AND U25961 ( .A(p_input[2211]), .B(p_input[12211]), .Z(n17308) );
  AND U25962 ( .A(p_input[32211]), .B(p_input[22211]), .Z(n17307) );
  AND U25963 ( .A(n17309), .B(n17310), .Z(o[2210]) );
  AND U25964 ( .A(p_input[2210]), .B(p_input[12210]), .Z(n17310) );
  AND U25965 ( .A(p_input[32210]), .B(p_input[22210]), .Z(n17309) );
  AND U25966 ( .A(n17311), .B(n17312), .Z(o[220]) );
  AND U25967 ( .A(p_input[20220]), .B(p_input[10220]), .Z(n17312) );
  AND U25968 ( .A(p_input[30220]), .B(p_input[220]), .Z(n17311) );
  AND U25969 ( .A(n17313), .B(n17314), .Z(o[2209]) );
  AND U25970 ( .A(p_input[2209]), .B(p_input[12209]), .Z(n17314) );
  AND U25971 ( .A(p_input[32209]), .B(p_input[22209]), .Z(n17313) );
  AND U25972 ( .A(n17315), .B(n17316), .Z(o[2208]) );
  AND U25973 ( .A(p_input[2208]), .B(p_input[12208]), .Z(n17316) );
  AND U25974 ( .A(p_input[32208]), .B(p_input[22208]), .Z(n17315) );
  AND U25975 ( .A(n17317), .B(n17318), .Z(o[2207]) );
  AND U25976 ( .A(p_input[2207]), .B(p_input[12207]), .Z(n17318) );
  AND U25977 ( .A(p_input[32207]), .B(p_input[22207]), .Z(n17317) );
  AND U25978 ( .A(n17319), .B(n17320), .Z(o[2206]) );
  AND U25979 ( .A(p_input[2206]), .B(p_input[12206]), .Z(n17320) );
  AND U25980 ( .A(p_input[32206]), .B(p_input[22206]), .Z(n17319) );
  AND U25981 ( .A(n17321), .B(n17322), .Z(o[2205]) );
  AND U25982 ( .A(p_input[2205]), .B(p_input[12205]), .Z(n17322) );
  AND U25983 ( .A(p_input[32205]), .B(p_input[22205]), .Z(n17321) );
  AND U25984 ( .A(n17323), .B(n17324), .Z(o[2204]) );
  AND U25985 ( .A(p_input[2204]), .B(p_input[12204]), .Z(n17324) );
  AND U25986 ( .A(p_input[32204]), .B(p_input[22204]), .Z(n17323) );
  AND U25987 ( .A(n17325), .B(n17326), .Z(o[2203]) );
  AND U25988 ( .A(p_input[2203]), .B(p_input[12203]), .Z(n17326) );
  AND U25989 ( .A(p_input[32203]), .B(p_input[22203]), .Z(n17325) );
  AND U25990 ( .A(n17327), .B(n17328), .Z(o[2202]) );
  AND U25991 ( .A(p_input[2202]), .B(p_input[12202]), .Z(n17328) );
  AND U25992 ( .A(p_input[32202]), .B(p_input[22202]), .Z(n17327) );
  AND U25993 ( .A(n17329), .B(n17330), .Z(o[2201]) );
  AND U25994 ( .A(p_input[2201]), .B(p_input[12201]), .Z(n17330) );
  AND U25995 ( .A(p_input[32201]), .B(p_input[22201]), .Z(n17329) );
  AND U25996 ( .A(n17331), .B(n17332), .Z(o[2200]) );
  AND U25997 ( .A(p_input[2200]), .B(p_input[12200]), .Z(n17332) );
  AND U25998 ( .A(p_input[32200]), .B(p_input[22200]), .Z(n17331) );
  AND U25999 ( .A(n17333), .B(n17334), .Z(o[21]) );
  AND U26000 ( .A(p_input[20021]), .B(p_input[10021]), .Z(n17334) );
  AND U26001 ( .A(p_input[30021]), .B(p_input[21]), .Z(n17333) );
  AND U26002 ( .A(n17335), .B(n17336), .Z(o[219]) );
  AND U26003 ( .A(p_input[20219]), .B(p_input[10219]), .Z(n17336) );
  AND U26004 ( .A(p_input[30219]), .B(p_input[219]), .Z(n17335) );
  AND U26005 ( .A(n17337), .B(n17338), .Z(o[2199]) );
  AND U26006 ( .A(p_input[2199]), .B(p_input[12199]), .Z(n17338) );
  AND U26007 ( .A(p_input[32199]), .B(p_input[22199]), .Z(n17337) );
  AND U26008 ( .A(n17339), .B(n17340), .Z(o[2198]) );
  AND U26009 ( .A(p_input[2198]), .B(p_input[12198]), .Z(n17340) );
  AND U26010 ( .A(p_input[32198]), .B(p_input[22198]), .Z(n17339) );
  AND U26011 ( .A(n17341), .B(n17342), .Z(o[2197]) );
  AND U26012 ( .A(p_input[2197]), .B(p_input[12197]), .Z(n17342) );
  AND U26013 ( .A(p_input[32197]), .B(p_input[22197]), .Z(n17341) );
  AND U26014 ( .A(n17343), .B(n17344), .Z(o[2196]) );
  AND U26015 ( .A(p_input[2196]), .B(p_input[12196]), .Z(n17344) );
  AND U26016 ( .A(p_input[32196]), .B(p_input[22196]), .Z(n17343) );
  AND U26017 ( .A(n17345), .B(n17346), .Z(o[2195]) );
  AND U26018 ( .A(p_input[2195]), .B(p_input[12195]), .Z(n17346) );
  AND U26019 ( .A(p_input[32195]), .B(p_input[22195]), .Z(n17345) );
  AND U26020 ( .A(n17347), .B(n17348), .Z(o[2194]) );
  AND U26021 ( .A(p_input[2194]), .B(p_input[12194]), .Z(n17348) );
  AND U26022 ( .A(p_input[32194]), .B(p_input[22194]), .Z(n17347) );
  AND U26023 ( .A(n17349), .B(n17350), .Z(o[2193]) );
  AND U26024 ( .A(p_input[2193]), .B(p_input[12193]), .Z(n17350) );
  AND U26025 ( .A(p_input[32193]), .B(p_input[22193]), .Z(n17349) );
  AND U26026 ( .A(n17351), .B(n17352), .Z(o[2192]) );
  AND U26027 ( .A(p_input[2192]), .B(p_input[12192]), .Z(n17352) );
  AND U26028 ( .A(p_input[32192]), .B(p_input[22192]), .Z(n17351) );
  AND U26029 ( .A(n17353), .B(n17354), .Z(o[2191]) );
  AND U26030 ( .A(p_input[2191]), .B(p_input[12191]), .Z(n17354) );
  AND U26031 ( .A(p_input[32191]), .B(p_input[22191]), .Z(n17353) );
  AND U26032 ( .A(n17355), .B(n17356), .Z(o[2190]) );
  AND U26033 ( .A(p_input[2190]), .B(p_input[12190]), .Z(n17356) );
  AND U26034 ( .A(p_input[32190]), .B(p_input[22190]), .Z(n17355) );
  AND U26035 ( .A(n17357), .B(n17358), .Z(o[218]) );
  AND U26036 ( .A(p_input[20218]), .B(p_input[10218]), .Z(n17358) );
  AND U26037 ( .A(p_input[30218]), .B(p_input[218]), .Z(n17357) );
  AND U26038 ( .A(n17359), .B(n17360), .Z(o[2189]) );
  AND U26039 ( .A(p_input[2189]), .B(p_input[12189]), .Z(n17360) );
  AND U26040 ( .A(p_input[32189]), .B(p_input[22189]), .Z(n17359) );
  AND U26041 ( .A(n17361), .B(n17362), .Z(o[2188]) );
  AND U26042 ( .A(p_input[2188]), .B(p_input[12188]), .Z(n17362) );
  AND U26043 ( .A(p_input[32188]), .B(p_input[22188]), .Z(n17361) );
  AND U26044 ( .A(n17363), .B(n17364), .Z(o[2187]) );
  AND U26045 ( .A(p_input[2187]), .B(p_input[12187]), .Z(n17364) );
  AND U26046 ( .A(p_input[32187]), .B(p_input[22187]), .Z(n17363) );
  AND U26047 ( .A(n17365), .B(n17366), .Z(o[2186]) );
  AND U26048 ( .A(p_input[2186]), .B(p_input[12186]), .Z(n17366) );
  AND U26049 ( .A(p_input[32186]), .B(p_input[22186]), .Z(n17365) );
  AND U26050 ( .A(n17367), .B(n17368), .Z(o[2185]) );
  AND U26051 ( .A(p_input[2185]), .B(p_input[12185]), .Z(n17368) );
  AND U26052 ( .A(p_input[32185]), .B(p_input[22185]), .Z(n17367) );
  AND U26053 ( .A(n17369), .B(n17370), .Z(o[2184]) );
  AND U26054 ( .A(p_input[2184]), .B(p_input[12184]), .Z(n17370) );
  AND U26055 ( .A(p_input[32184]), .B(p_input[22184]), .Z(n17369) );
  AND U26056 ( .A(n17371), .B(n17372), .Z(o[2183]) );
  AND U26057 ( .A(p_input[2183]), .B(p_input[12183]), .Z(n17372) );
  AND U26058 ( .A(p_input[32183]), .B(p_input[22183]), .Z(n17371) );
  AND U26059 ( .A(n17373), .B(n17374), .Z(o[2182]) );
  AND U26060 ( .A(p_input[2182]), .B(p_input[12182]), .Z(n17374) );
  AND U26061 ( .A(p_input[32182]), .B(p_input[22182]), .Z(n17373) );
  AND U26062 ( .A(n17375), .B(n17376), .Z(o[2181]) );
  AND U26063 ( .A(p_input[2181]), .B(p_input[12181]), .Z(n17376) );
  AND U26064 ( .A(p_input[32181]), .B(p_input[22181]), .Z(n17375) );
  AND U26065 ( .A(n17377), .B(n17378), .Z(o[2180]) );
  AND U26066 ( .A(p_input[2180]), .B(p_input[12180]), .Z(n17378) );
  AND U26067 ( .A(p_input[32180]), .B(p_input[22180]), .Z(n17377) );
  AND U26068 ( .A(n17379), .B(n17380), .Z(o[217]) );
  AND U26069 ( .A(p_input[20217]), .B(p_input[10217]), .Z(n17380) );
  AND U26070 ( .A(p_input[30217]), .B(p_input[217]), .Z(n17379) );
  AND U26071 ( .A(n17381), .B(n17382), .Z(o[2179]) );
  AND U26072 ( .A(p_input[2179]), .B(p_input[12179]), .Z(n17382) );
  AND U26073 ( .A(p_input[32179]), .B(p_input[22179]), .Z(n17381) );
  AND U26074 ( .A(n17383), .B(n17384), .Z(o[2178]) );
  AND U26075 ( .A(p_input[2178]), .B(p_input[12178]), .Z(n17384) );
  AND U26076 ( .A(p_input[32178]), .B(p_input[22178]), .Z(n17383) );
  AND U26077 ( .A(n17385), .B(n17386), .Z(o[2177]) );
  AND U26078 ( .A(p_input[2177]), .B(p_input[12177]), .Z(n17386) );
  AND U26079 ( .A(p_input[32177]), .B(p_input[22177]), .Z(n17385) );
  AND U26080 ( .A(n17387), .B(n17388), .Z(o[2176]) );
  AND U26081 ( .A(p_input[2176]), .B(p_input[12176]), .Z(n17388) );
  AND U26082 ( .A(p_input[32176]), .B(p_input[22176]), .Z(n17387) );
  AND U26083 ( .A(n17389), .B(n17390), .Z(o[2175]) );
  AND U26084 ( .A(p_input[2175]), .B(p_input[12175]), .Z(n17390) );
  AND U26085 ( .A(p_input[32175]), .B(p_input[22175]), .Z(n17389) );
  AND U26086 ( .A(n17391), .B(n17392), .Z(o[2174]) );
  AND U26087 ( .A(p_input[2174]), .B(p_input[12174]), .Z(n17392) );
  AND U26088 ( .A(p_input[32174]), .B(p_input[22174]), .Z(n17391) );
  AND U26089 ( .A(n17393), .B(n17394), .Z(o[2173]) );
  AND U26090 ( .A(p_input[2173]), .B(p_input[12173]), .Z(n17394) );
  AND U26091 ( .A(p_input[32173]), .B(p_input[22173]), .Z(n17393) );
  AND U26092 ( .A(n17395), .B(n17396), .Z(o[2172]) );
  AND U26093 ( .A(p_input[2172]), .B(p_input[12172]), .Z(n17396) );
  AND U26094 ( .A(p_input[32172]), .B(p_input[22172]), .Z(n17395) );
  AND U26095 ( .A(n17397), .B(n17398), .Z(o[2171]) );
  AND U26096 ( .A(p_input[2171]), .B(p_input[12171]), .Z(n17398) );
  AND U26097 ( .A(p_input[32171]), .B(p_input[22171]), .Z(n17397) );
  AND U26098 ( .A(n17399), .B(n17400), .Z(o[2170]) );
  AND U26099 ( .A(p_input[2170]), .B(p_input[12170]), .Z(n17400) );
  AND U26100 ( .A(p_input[32170]), .B(p_input[22170]), .Z(n17399) );
  AND U26101 ( .A(n17401), .B(n17402), .Z(o[216]) );
  AND U26102 ( .A(p_input[20216]), .B(p_input[10216]), .Z(n17402) );
  AND U26103 ( .A(p_input[30216]), .B(p_input[216]), .Z(n17401) );
  AND U26104 ( .A(n17403), .B(n17404), .Z(o[2169]) );
  AND U26105 ( .A(p_input[2169]), .B(p_input[12169]), .Z(n17404) );
  AND U26106 ( .A(p_input[32169]), .B(p_input[22169]), .Z(n17403) );
  AND U26107 ( .A(n17405), .B(n17406), .Z(o[2168]) );
  AND U26108 ( .A(p_input[2168]), .B(p_input[12168]), .Z(n17406) );
  AND U26109 ( .A(p_input[32168]), .B(p_input[22168]), .Z(n17405) );
  AND U26110 ( .A(n17407), .B(n17408), .Z(o[2167]) );
  AND U26111 ( .A(p_input[2167]), .B(p_input[12167]), .Z(n17408) );
  AND U26112 ( .A(p_input[32167]), .B(p_input[22167]), .Z(n17407) );
  AND U26113 ( .A(n17409), .B(n17410), .Z(o[2166]) );
  AND U26114 ( .A(p_input[2166]), .B(p_input[12166]), .Z(n17410) );
  AND U26115 ( .A(p_input[32166]), .B(p_input[22166]), .Z(n17409) );
  AND U26116 ( .A(n17411), .B(n17412), .Z(o[2165]) );
  AND U26117 ( .A(p_input[2165]), .B(p_input[12165]), .Z(n17412) );
  AND U26118 ( .A(p_input[32165]), .B(p_input[22165]), .Z(n17411) );
  AND U26119 ( .A(n17413), .B(n17414), .Z(o[2164]) );
  AND U26120 ( .A(p_input[2164]), .B(p_input[12164]), .Z(n17414) );
  AND U26121 ( .A(p_input[32164]), .B(p_input[22164]), .Z(n17413) );
  AND U26122 ( .A(n17415), .B(n17416), .Z(o[2163]) );
  AND U26123 ( .A(p_input[2163]), .B(p_input[12163]), .Z(n17416) );
  AND U26124 ( .A(p_input[32163]), .B(p_input[22163]), .Z(n17415) );
  AND U26125 ( .A(n17417), .B(n17418), .Z(o[2162]) );
  AND U26126 ( .A(p_input[2162]), .B(p_input[12162]), .Z(n17418) );
  AND U26127 ( .A(p_input[32162]), .B(p_input[22162]), .Z(n17417) );
  AND U26128 ( .A(n17419), .B(n17420), .Z(o[2161]) );
  AND U26129 ( .A(p_input[2161]), .B(p_input[12161]), .Z(n17420) );
  AND U26130 ( .A(p_input[32161]), .B(p_input[22161]), .Z(n17419) );
  AND U26131 ( .A(n17421), .B(n17422), .Z(o[2160]) );
  AND U26132 ( .A(p_input[2160]), .B(p_input[12160]), .Z(n17422) );
  AND U26133 ( .A(p_input[32160]), .B(p_input[22160]), .Z(n17421) );
  AND U26134 ( .A(n17423), .B(n17424), .Z(o[215]) );
  AND U26135 ( .A(p_input[20215]), .B(p_input[10215]), .Z(n17424) );
  AND U26136 ( .A(p_input[30215]), .B(p_input[215]), .Z(n17423) );
  AND U26137 ( .A(n17425), .B(n17426), .Z(o[2159]) );
  AND U26138 ( .A(p_input[2159]), .B(p_input[12159]), .Z(n17426) );
  AND U26139 ( .A(p_input[32159]), .B(p_input[22159]), .Z(n17425) );
  AND U26140 ( .A(n17427), .B(n17428), .Z(o[2158]) );
  AND U26141 ( .A(p_input[2158]), .B(p_input[12158]), .Z(n17428) );
  AND U26142 ( .A(p_input[32158]), .B(p_input[22158]), .Z(n17427) );
  AND U26143 ( .A(n17429), .B(n17430), .Z(o[2157]) );
  AND U26144 ( .A(p_input[2157]), .B(p_input[12157]), .Z(n17430) );
  AND U26145 ( .A(p_input[32157]), .B(p_input[22157]), .Z(n17429) );
  AND U26146 ( .A(n17431), .B(n17432), .Z(o[2156]) );
  AND U26147 ( .A(p_input[2156]), .B(p_input[12156]), .Z(n17432) );
  AND U26148 ( .A(p_input[32156]), .B(p_input[22156]), .Z(n17431) );
  AND U26149 ( .A(n17433), .B(n17434), .Z(o[2155]) );
  AND U26150 ( .A(p_input[2155]), .B(p_input[12155]), .Z(n17434) );
  AND U26151 ( .A(p_input[32155]), .B(p_input[22155]), .Z(n17433) );
  AND U26152 ( .A(n17435), .B(n17436), .Z(o[2154]) );
  AND U26153 ( .A(p_input[2154]), .B(p_input[12154]), .Z(n17436) );
  AND U26154 ( .A(p_input[32154]), .B(p_input[22154]), .Z(n17435) );
  AND U26155 ( .A(n17437), .B(n17438), .Z(o[2153]) );
  AND U26156 ( .A(p_input[2153]), .B(p_input[12153]), .Z(n17438) );
  AND U26157 ( .A(p_input[32153]), .B(p_input[22153]), .Z(n17437) );
  AND U26158 ( .A(n17439), .B(n17440), .Z(o[2152]) );
  AND U26159 ( .A(p_input[2152]), .B(p_input[12152]), .Z(n17440) );
  AND U26160 ( .A(p_input[32152]), .B(p_input[22152]), .Z(n17439) );
  AND U26161 ( .A(n17441), .B(n17442), .Z(o[2151]) );
  AND U26162 ( .A(p_input[2151]), .B(p_input[12151]), .Z(n17442) );
  AND U26163 ( .A(p_input[32151]), .B(p_input[22151]), .Z(n17441) );
  AND U26164 ( .A(n17443), .B(n17444), .Z(o[2150]) );
  AND U26165 ( .A(p_input[2150]), .B(p_input[12150]), .Z(n17444) );
  AND U26166 ( .A(p_input[32150]), .B(p_input[22150]), .Z(n17443) );
  AND U26167 ( .A(n17445), .B(n17446), .Z(o[214]) );
  AND U26168 ( .A(p_input[20214]), .B(p_input[10214]), .Z(n17446) );
  AND U26169 ( .A(p_input[30214]), .B(p_input[214]), .Z(n17445) );
  AND U26170 ( .A(n17447), .B(n17448), .Z(o[2149]) );
  AND U26171 ( .A(p_input[2149]), .B(p_input[12149]), .Z(n17448) );
  AND U26172 ( .A(p_input[32149]), .B(p_input[22149]), .Z(n17447) );
  AND U26173 ( .A(n17449), .B(n17450), .Z(o[2148]) );
  AND U26174 ( .A(p_input[2148]), .B(p_input[12148]), .Z(n17450) );
  AND U26175 ( .A(p_input[32148]), .B(p_input[22148]), .Z(n17449) );
  AND U26176 ( .A(n17451), .B(n17452), .Z(o[2147]) );
  AND U26177 ( .A(p_input[2147]), .B(p_input[12147]), .Z(n17452) );
  AND U26178 ( .A(p_input[32147]), .B(p_input[22147]), .Z(n17451) );
  AND U26179 ( .A(n17453), .B(n17454), .Z(o[2146]) );
  AND U26180 ( .A(p_input[2146]), .B(p_input[12146]), .Z(n17454) );
  AND U26181 ( .A(p_input[32146]), .B(p_input[22146]), .Z(n17453) );
  AND U26182 ( .A(n17455), .B(n17456), .Z(o[2145]) );
  AND U26183 ( .A(p_input[2145]), .B(p_input[12145]), .Z(n17456) );
  AND U26184 ( .A(p_input[32145]), .B(p_input[22145]), .Z(n17455) );
  AND U26185 ( .A(n17457), .B(n17458), .Z(o[2144]) );
  AND U26186 ( .A(p_input[2144]), .B(p_input[12144]), .Z(n17458) );
  AND U26187 ( .A(p_input[32144]), .B(p_input[22144]), .Z(n17457) );
  AND U26188 ( .A(n17459), .B(n17460), .Z(o[2143]) );
  AND U26189 ( .A(p_input[2143]), .B(p_input[12143]), .Z(n17460) );
  AND U26190 ( .A(p_input[32143]), .B(p_input[22143]), .Z(n17459) );
  AND U26191 ( .A(n17461), .B(n17462), .Z(o[2142]) );
  AND U26192 ( .A(p_input[2142]), .B(p_input[12142]), .Z(n17462) );
  AND U26193 ( .A(p_input[32142]), .B(p_input[22142]), .Z(n17461) );
  AND U26194 ( .A(n17463), .B(n17464), .Z(o[2141]) );
  AND U26195 ( .A(p_input[2141]), .B(p_input[12141]), .Z(n17464) );
  AND U26196 ( .A(p_input[32141]), .B(p_input[22141]), .Z(n17463) );
  AND U26197 ( .A(n17465), .B(n17466), .Z(o[2140]) );
  AND U26198 ( .A(p_input[2140]), .B(p_input[12140]), .Z(n17466) );
  AND U26199 ( .A(p_input[32140]), .B(p_input[22140]), .Z(n17465) );
  AND U26200 ( .A(n17467), .B(n17468), .Z(o[213]) );
  AND U26201 ( .A(p_input[20213]), .B(p_input[10213]), .Z(n17468) );
  AND U26202 ( .A(p_input[30213]), .B(p_input[213]), .Z(n17467) );
  AND U26203 ( .A(n17469), .B(n17470), .Z(o[2139]) );
  AND U26204 ( .A(p_input[2139]), .B(p_input[12139]), .Z(n17470) );
  AND U26205 ( .A(p_input[32139]), .B(p_input[22139]), .Z(n17469) );
  AND U26206 ( .A(n17471), .B(n17472), .Z(o[2138]) );
  AND U26207 ( .A(p_input[2138]), .B(p_input[12138]), .Z(n17472) );
  AND U26208 ( .A(p_input[32138]), .B(p_input[22138]), .Z(n17471) );
  AND U26209 ( .A(n17473), .B(n17474), .Z(o[2137]) );
  AND U26210 ( .A(p_input[2137]), .B(p_input[12137]), .Z(n17474) );
  AND U26211 ( .A(p_input[32137]), .B(p_input[22137]), .Z(n17473) );
  AND U26212 ( .A(n17475), .B(n17476), .Z(o[2136]) );
  AND U26213 ( .A(p_input[2136]), .B(p_input[12136]), .Z(n17476) );
  AND U26214 ( .A(p_input[32136]), .B(p_input[22136]), .Z(n17475) );
  AND U26215 ( .A(n17477), .B(n17478), .Z(o[2135]) );
  AND U26216 ( .A(p_input[2135]), .B(p_input[12135]), .Z(n17478) );
  AND U26217 ( .A(p_input[32135]), .B(p_input[22135]), .Z(n17477) );
  AND U26218 ( .A(n17479), .B(n17480), .Z(o[2134]) );
  AND U26219 ( .A(p_input[2134]), .B(p_input[12134]), .Z(n17480) );
  AND U26220 ( .A(p_input[32134]), .B(p_input[22134]), .Z(n17479) );
  AND U26221 ( .A(n17481), .B(n17482), .Z(o[2133]) );
  AND U26222 ( .A(p_input[2133]), .B(p_input[12133]), .Z(n17482) );
  AND U26223 ( .A(p_input[32133]), .B(p_input[22133]), .Z(n17481) );
  AND U26224 ( .A(n17483), .B(n17484), .Z(o[2132]) );
  AND U26225 ( .A(p_input[2132]), .B(p_input[12132]), .Z(n17484) );
  AND U26226 ( .A(p_input[32132]), .B(p_input[22132]), .Z(n17483) );
  AND U26227 ( .A(n17485), .B(n17486), .Z(o[2131]) );
  AND U26228 ( .A(p_input[2131]), .B(p_input[12131]), .Z(n17486) );
  AND U26229 ( .A(p_input[32131]), .B(p_input[22131]), .Z(n17485) );
  AND U26230 ( .A(n17487), .B(n17488), .Z(o[2130]) );
  AND U26231 ( .A(p_input[2130]), .B(p_input[12130]), .Z(n17488) );
  AND U26232 ( .A(p_input[32130]), .B(p_input[22130]), .Z(n17487) );
  AND U26233 ( .A(n17489), .B(n17490), .Z(o[212]) );
  AND U26234 ( .A(p_input[20212]), .B(p_input[10212]), .Z(n17490) );
  AND U26235 ( .A(p_input[30212]), .B(p_input[212]), .Z(n17489) );
  AND U26236 ( .A(n17491), .B(n17492), .Z(o[2129]) );
  AND U26237 ( .A(p_input[2129]), .B(p_input[12129]), .Z(n17492) );
  AND U26238 ( .A(p_input[32129]), .B(p_input[22129]), .Z(n17491) );
  AND U26239 ( .A(n17493), .B(n17494), .Z(o[2128]) );
  AND U26240 ( .A(p_input[2128]), .B(p_input[12128]), .Z(n17494) );
  AND U26241 ( .A(p_input[32128]), .B(p_input[22128]), .Z(n17493) );
  AND U26242 ( .A(n17495), .B(n17496), .Z(o[2127]) );
  AND U26243 ( .A(p_input[2127]), .B(p_input[12127]), .Z(n17496) );
  AND U26244 ( .A(p_input[32127]), .B(p_input[22127]), .Z(n17495) );
  AND U26245 ( .A(n17497), .B(n17498), .Z(o[2126]) );
  AND U26246 ( .A(p_input[2126]), .B(p_input[12126]), .Z(n17498) );
  AND U26247 ( .A(p_input[32126]), .B(p_input[22126]), .Z(n17497) );
  AND U26248 ( .A(n17499), .B(n17500), .Z(o[2125]) );
  AND U26249 ( .A(p_input[2125]), .B(p_input[12125]), .Z(n17500) );
  AND U26250 ( .A(p_input[32125]), .B(p_input[22125]), .Z(n17499) );
  AND U26251 ( .A(n17501), .B(n17502), .Z(o[2124]) );
  AND U26252 ( .A(p_input[2124]), .B(p_input[12124]), .Z(n17502) );
  AND U26253 ( .A(p_input[32124]), .B(p_input[22124]), .Z(n17501) );
  AND U26254 ( .A(n17503), .B(n17504), .Z(o[2123]) );
  AND U26255 ( .A(p_input[2123]), .B(p_input[12123]), .Z(n17504) );
  AND U26256 ( .A(p_input[32123]), .B(p_input[22123]), .Z(n17503) );
  AND U26257 ( .A(n17505), .B(n17506), .Z(o[2122]) );
  AND U26258 ( .A(p_input[2122]), .B(p_input[12122]), .Z(n17506) );
  AND U26259 ( .A(p_input[32122]), .B(p_input[22122]), .Z(n17505) );
  AND U26260 ( .A(n17507), .B(n17508), .Z(o[2121]) );
  AND U26261 ( .A(p_input[2121]), .B(p_input[12121]), .Z(n17508) );
  AND U26262 ( .A(p_input[32121]), .B(p_input[22121]), .Z(n17507) );
  AND U26263 ( .A(n17509), .B(n17510), .Z(o[2120]) );
  AND U26264 ( .A(p_input[2120]), .B(p_input[12120]), .Z(n17510) );
  AND U26265 ( .A(p_input[32120]), .B(p_input[22120]), .Z(n17509) );
  AND U26266 ( .A(n17511), .B(n17512), .Z(o[211]) );
  AND U26267 ( .A(p_input[20211]), .B(p_input[10211]), .Z(n17512) );
  AND U26268 ( .A(p_input[30211]), .B(p_input[211]), .Z(n17511) );
  AND U26269 ( .A(n17513), .B(n17514), .Z(o[2119]) );
  AND U26270 ( .A(p_input[2119]), .B(p_input[12119]), .Z(n17514) );
  AND U26271 ( .A(p_input[32119]), .B(p_input[22119]), .Z(n17513) );
  AND U26272 ( .A(n17515), .B(n17516), .Z(o[2118]) );
  AND U26273 ( .A(p_input[2118]), .B(p_input[12118]), .Z(n17516) );
  AND U26274 ( .A(p_input[32118]), .B(p_input[22118]), .Z(n17515) );
  AND U26275 ( .A(n17517), .B(n17518), .Z(o[2117]) );
  AND U26276 ( .A(p_input[2117]), .B(p_input[12117]), .Z(n17518) );
  AND U26277 ( .A(p_input[32117]), .B(p_input[22117]), .Z(n17517) );
  AND U26278 ( .A(n17519), .B(n17520), .Z(o[2116]) );
  AND U26279 ( .A(p_input[2116]), .B(p_input[12116]), .Z(n17520) );
  AND U26280 ( .A(p_input[32116]), .B(p_input[22116]), .Z(n17519) );
  AND U26281 ( .A(n17521), .B(n17522), .Z(o[2115]) );
  AND U26282 ( .A(p_input[2115]), .B(p_input[12115]), .Z(n17522) );
  AND U26283 ( .A(p_input[32115]), .B(p_input[22115]), .Z(n17521) );
  AND U26284 ( .A(n17523), .B(n17524), .Z(o[2114]) );
  AND U26285 ( .A(p_input[2114]), .B(p_input[12114]), .Z(n17524) );
  AND U26286 ( .A(p_input[32114]), .B(p_input[22114]), .Z(n17523) );
  AND U26287 ( .A(n17525), .B(n17526), .Z(o[2113]) );
  AND U26288 ( .A(p_input[2113]), .B(p_input[12113]), .Z(n17526) );
  AND U26289 ( .A(p_input[32113]), .B(p_input[22113]), .Z(n17525) );
  AND U26290 ( .A(n17527), .B(n17528), .Z(o[2112]) );
  AND U26291 ( .A(p_input[2112]), .B(p_input[12112]), .Z(n17528) );
  AND U26292 ( .A(p_input[32112]), .B(p_input[22112]), .Z(n17527) );
  AND U26293 ( .A(n17529), .B(n17530), .Z(o[2111]) );
  AND U26294 ( .A(p_input[2111]), .B(p_input[12111]), .Z(n17530) );
  AND U26295 ( .A(p_input[32111]), .B(p_input[22111]), .Z(n17529) );
  AND U26296 ( .A(n17531), .B(n17532), .Z(o[2110]) );
  AND U26297 ( .A(p_input[2110]), .B(p_input[12110]), .Z(n17532) );
  AND U26298 ( .A(p_input[32110]), .B(p_input[22110]), .Z(n17531) );
  AND U26299 ( .A(n17533), .B(n17534), .Z(o[210]) );
  AND U26300 ( .A(p_input[20210]), .B(p_input[10210]), .Z(n17534) );
  AND U26301 ( .A(p_input[30210]), .B(p_input[210]), .Z(n17533) );
  AND U26302 ( .A(n17535), .B(n17536), .Z(o[2109]) );
  AND U26303 ( .A(p_input[2109]), .B(p_input[12109]), .Z(n17536) );
  AND U26304 ( .A(p_input[32109]), .B(p_input[22109]), .Z(n17535) );
  AND U26305 ( .A(n17537), .B(n17538), .Z(o[2108]) );
  AND U26306 ( .A(p_input[2108]), .B(p_input[12108]), .Z(n17538) );
  AND U26307 ( .A(p_input[32108]), .B(p_input[22108]), .Z(n17537) );
  AND U26308 ( .A(n17539), .B(n17540), .Z(o[2107]) );
  AND U26309 ( .A(p_input[2107]), .B(p_input[12107]), .Z(n17540) );
  AND U26310 ( .A(p_input[32107]), .B(p_input[22107]), .Z(n17539) );
  AND U26311 ( .A(n17541), .B(n17542), .Z(o[2106]) );
  AND U26312 ( .A(p_input[2106]), .B(p_input[12106]), .Z(n17542) );
  AND U26313 ( .A(p_input[32106]), .B(p_input[22106]), .Z(n17541) );
  AND U26314 ( .A(n17543), .B(n17544), .Z(o[2105]) );
  AND U26315 ( .A(p_input[2105]), .B(p_input[12105]), .Z(n17544) );
  AND U26316 ( .A(p_input[32105]), .B(p_input[22105]), .Z(n17543) );
  AND U26317 ( .A(n17545), .B(n17546), .Z(o[2104]) );
  AND U26318 ( .A(p_input[2104]), .B(p_input[12104]), .Z(n17546) );
  AND U26319 ( .A(p_input[32104]), .B(p_input[22104]), .Z(n17545) );
  AND U26320 ( .A(n17547), .B(n17548), .Z(o[2103]) );
  AND U26321 ( .A(p_input[2103]), .B(p_input[12103]), .Z(n17548) );
  AND U26322 ( .A(p_input[32103]), .B(p_input[22103]), .Z(n17547) );
  AND U26323 ( .A(n17549), .B(n17550), .Z(o[2102]) );
  AND U26324 ( .A(p_input[2102]), .B(p_input[12102]), .Z(n17550) );
  AND U26325 ( .A(p_input[32102]), .B(p_input[22102]), .Z(n17549) );
  AND U26326 ( .A(n17551), .B(n17552), .Z(o[2101]) );
  AND U26327 ( .A(p_input[2101]), .B(p_input[12101]), .Z(n17552) );
  AND U26328 ( .A(p_input[32101]), .B(p_input[22101]), .Z(n17551) );
  AND U26329 ( .A(n17553), .B(n17554), .Z(o[2100]) );
  AND U26330 ( .A(p_input[2100]), .B(p_input[12100]), .Z(n17554) );
  AND U26331 ( .A(p_input[32100]), .B(p_input[22100]), .Z(n17553) );
  AND U26332 ( .A(n17555), .B(n17556), .Z(o[20]) );
  AND U26333 ( .A(p_input[20020]), .B(p_input[10020]), .Z(n17556) );
  AND U26334 ( .A(p_input[30020]), .B(p_input[20]), .Z(n17555) );
  AND U26335 ( .A(n17557), .B(n17558), .Z(o[209]) );
  AND U26336 ( .A(p_input[20209]), .B(p_input[10209]), .Z(n17558) );
  AND U26337 ( .A(p_input[30209]), .B(p_input[209]), .Z(n17557) );
  AND U26338 ( .A(n17559), .B(n17560), .Z(o[2099]) );
  AND U26339 ( .A(p_input[2099]), .B(p_input[12099]), .Z(n17560) );
  AND U26340 ( .A(p_input[32099]), .B(p_input[22099]), .Z(n17559) );
  AND U26341 ( .A(n17561), .B(n17562), .Z(o[2098]) );
  AND U26342 ( .A(p_input[2098]), .B(p_input[12098]), .Z(n17562) );
  AND U26343 ( .A(p_input[32098]), .B(p_input[22098]), .Z(n17561) );
  AND U26344 ( .A(n17563), .B(n17564), .Z(o[2097]) );
  AND U26345 ( .A(p_input[2097]), .B(p_input[12097]), .Z(n17564) );
  AND U26346 ( .A(p_input[32097]), .B(p_input[22097]), .Z(n17563) );
  AND U26347 ( .A(n17565), .B(n17566), .Z(o[2096]) );
  AND U26348 ( .A(p_input[2096]), .B(p_input[12096]), .Z(n17566) );
  AND U26349 ( .A(p_input[32096]), .B(p_input[22096]), .Z(n17565) );
  AND U26350 ( .A(n17567), .B(n17568), .Z(o[2095]) );
  AND U26351 ( .A(p_input[2095]), .B(p_input[12095]), .Z(n17568) );
  AND U26352 ( .A(p_input[32095]), .B(p_input[22095]), .Z(n17567) );
  AND U26353 ( .A(n17569), .B(n17570), .Z(o[2094]) );
  AND U26354 ( .A(p_input[2094]), .B(p_input[12094]), .Z(n17570) );
  AND U26355 ( .A(p_input[32094]), .B(p_input[22094]), .Z(n17569) );
  AND U26356 ( .A(n17571), .B(n17572), .Z(o[2093]) );
  AND U26357 ( .A(p_input[2093]), .B(p_input[12093]), .Z(n17572) );
  AND U26358 ( .A(p_input[32093]), .B(p_input[22093]), .Z(n17571) );
  AND U26359 ( .A(n17573), .B(n17574), .Z(o[2092]) );
  AND U26360 ( .A(p_input[2092]), .B(p_input[12092]), .Z(n17574) );
  AND U26361 ( .A(p_input[32092]), .B(p_input[22092]), .Z(n17573) );
  AND U26362 ( .A(n17575), .B(n17576), .Z(o[2091]) );
  AND U26363 ( .A(p_input[2091]), .B(p_input[12091]), .Z(n17576) );
  AND U26364 ( .A(p_input[32091]), .B(p_input[22091]), .Z(n17575) );
  AND U26365 ( .A(n17577), .B(n17578), .Z(o[2090]) );
  AND U26366 ( .A(p_input[2090]), .B(p_input[12090]), .Z(n17578) );
  AND U26367 ( .A(p_input[32090]), .B(p_input[22090]), .Z(n17577) );
  AND U26368 ( .A(n17579), .B(n17580), .Z(o[208]) );
  AND U26369 ( .A(p_input[20208]), .B(p_input[10208]), .Z(n17580) );
  AND U26370 ( .A(p_input[30208]), .B(p_input[208]), .Z(n17579) );
  AND U26371 ( .A(n17581), .B(n17582), .Z(o[2089]) );
  AND U26372 ( .A(p_input[2089]), .B(p_input[12089]), .Z(n17582) );
  AND U26373 ( .A(p_input[32089]), .B(p_input[22089]), .Z(n17581) );
  AND U26374 ( .A(n17583), .B(n17584), .Z(o[2088]) );
  AND U26375 ( .A(p_input[2088]), .B(p_input[12088]), .Z(n17584) );
  AND U26376 ( .A(p_input[32088]), .B(p_input[22088]), .Z(n17583) );
  AND U26377 ( .A(n17585), .B(n17586), .Z(o[2087]) );
  AND U26378 ( .A(p_input[2087]), .B(p_input[12087]), .Z(n17586) );
  AND U26379 ( .A(p_input[32087]), .B(p_input[22087]), .Z(n17585) );
  AND U26380 ( .A(n17587), .B(n17588), .Z(o[2086]) );
  AND U26381 ( .A(p_input[2086]), .B(p_input[12086]), .Z(n17588) );
  AND U26382 ( .A(p_input[32086]), .B(p_input[22086]), .Z(n17587) );
  AND U26383 ( .A(n17589), .B(n17590), .Z(o[2085]) );
  AND U26384 ( .A(p_input[2085]), .B(p_input[12085]), .Z(n17590) );
  AND U26385 ( .A(p_input[32085]), .B(p_input[22085]), .Z(n17589) );
  AND U26386 ( .A(n17591), .B(n17592), .Z(o[2084]) );
  AND U26387 ( .A(p_input[2084]), .B(p_input[12084]), .Z(n17592) );
  AND U26388 ( .A(p_input[32084]), .B(p_input[22084]), .Z(n17591) );
  AND U26389 ( .A(n17593), .B(n17594), .Z(o[2083]) );
  AND U26390 ( .A(p_input[2083]), .B(p_input[12083]), .Z(n17594) );
  AND U26391 ( .A(p_input[32083]), .B(p_input[22083]), .Z(n17593) );
  AND U26392 ( .A(n17595), .B(n17596), .Z(o[2082]) );
  AND U26393 ( .A(p_input[2082]), .B(p_input[12082]), .Z(n17596) );
  AND U26394 ( .A(p_input[32082]), .B(p_input[22082]), .Z(n17595) );
  AND U26395 ( .A(n17597), .B(n17598), .Z(o[2081]) );
  AND U26396 ( .A(p_input[2081]), .B(p_input[12081]), .Z(n17598) );
  AND U26397 ( .A(p_input[32081]), .B(p_input[22081]), .Z(n17597) );
  AND U26398 ( .A(n17599), .B(n17600), .Z(o[2080]) );
  AND U26399 ( .A(p_input[2080]), .B(p_input[12080]), .Z(n17600) );
  AND U26400 ( .A(p_input[32080]), .B(p_input[22080]), .Z(n17599) );
  AND U26401 ( .A(n17601), .B(n17602), .Z(o[207]) );
  AND U26402 ( .A(p_input[20207]), .B(p_input[10207]), .Z(n17602) );
  AND U26403 ( .A(p_input[30207]), .B(p_input[207]), .Z(n17601) );
  AND U26404 ( .A(n17603), .B(n17604), .Z(o[2079]) );
  AND U26405 ( .A(p_input[2079]), .B(p_input[12079]), .Z(n17604) );
  AND U26406 ( .A(p_input[32079]), .B(p_input[22079]), .Z(n17603) );
  AND U26407 ( .A(n17605), .B(n17606), .Z(o[2078]) );
  AND U26408 ( .A(p_input[2078]), .B(p_input[12078]), .Z(n17606) );
  AND U26409 ( .A(p_input[32078]), .B(p_input[22078]), .Z(n17605) );
  AND U26410 ( .A(n17607), .B(n17608), .Z(o[2077]) );
  AND U26411 ( .A(p_input[2077]), .B(p_input[12077]), .Z(n17608) );
  AND U26412 ( .A(p_input[32077]), .B(p_input[22077]), .Z(n17607) );
  AND U26413 ( .A(n17609), .B(n17610), .Z(o[2076]) );
  AND U26414 ( .A(p_input[2076]), .B(p_input[12076]), .Z(n17610) );
  AND U26415 ( .A(p_input[32076]), .B(p_input[22076]), .Z(n17609) );
  AND U26416 ( .A(n17611), .B(n17612), .Z(o[2075]) );
  AND U26417 ( .A(p_input[2075]), .B(p_input[12075]), .Z(n17612) );
  AND U26418 ( .A(p_input[32075]), .B(p_input[22075]), .Z(n17611) );
  AND U26419 ( .A(n17613), .B(n17614), .Z(o[2074]) );
  AND U26420 ( .A(p_input[2074]), .B(p_input[12074]), .Z(n17614) );
  AND U26421 ( .A(p_input[32074]), .B(p_input[22074]), .Z(n17613) );
  AND U26422 ( .A(n17615), .B(n17616), .Z(o[2073]) );
  AND U26423 ( .A(p_input[2073]), .B(p_input[12073]), .Z(n17616) );
  AND U26424 ( .A(p_input[32073]), .B(p_input[22073]), .Z(n17615) );
  AND U26425 ( .A(n17617), .B(n17618), .Z(o[2072]) );
  AND U26426 ( .A(p_input[2072]), .B(p_input[12072]), .Z(n17618) );
  AND U26427 ( .A(p_input[32072]), .B(p_input[22072]), .Z(n17617) );
  AND U26428 ( .A(n17619), .B(n17620), .Z(o[2071]) );
  AND U26429 ( .A(p_input[2071]), .B(p_input[12071]), .Z(n17620) );
  AND U26430 ( .A(p_input[32071]), .B(p_input[22071]), .Z(n17619) );
  AND U26431 ( .A(n17621), .B(n17622), .Z(o[2070]) );
  AND U26432 ( .A(p_input[2070]), .B(p_input[12070]), .Z(n17622) );
  AND U26433 ( .A(p_input[32070]), .B(p_input[22070]), .Z(n17621) );
  AND U26434 ( .A(n17623), .B(n17624), .Z(o[206]) );
  AND U26435 ( .A(p_input[20206]), .B(p_input[10206]), .Z(n17624) );
  AND U26436 ( .A(p_input[30206]), .B(p_input[206]), .Z(n17623) );
  AND U26437 ( .A(n17625), .B(n17626), .Z(o[2069]) );
  AND U26438 ( .A(p_input[2069]), .B(p_input[12069]), .Z(n17626) );
  AND U26439 ( .A(p_input[32069]), .B(p_input[22069]), .Z(n17625) );
  AND U26440 ( .A(n17627), .B(n17628), .Z(o[2068]) );
  AND U26441 ( .A(p_input[2068]), .B(p_input[12068]), .Z(n17628) );
  AND U26442 ( .A(p_input[32068]), .B(p_input[22068]), .Z(n17627) );
  AND U26443 ( .A(n17629), .B(n17630), .Z(o[2067]) );
  AND U26444 ( .A(p_input[2067]), .B(p_input[12067]), .Z(n17630) );
  AND U26445 ( .A(p_input[32067]), .B(p_input[22067]), .Z(n17629) );
  AND U26446 ( .A(n17631), .B(n17632), .Z(o[2066]) );
  AND U26447 ( .A(p_input[2066]), .B(p_input[12066]), .Z(n17632) );
  AND U26448 ( .A(p_input[32066]), .B(p_input[22066]), .Z(n17631) );
  AND U26449 ( .A(n17633), .B(n17634), .Z(o[2065]) );
  AND U26450 ( .A(p_input[2065]), .B(p_input[12065]), .Z(n17634) );
  AND U26451 ( .A(p_input[32065]), .B(p_input[22065]), .Z(n17633) );
  AND U26452 ( .A(n17635), .B(n17636), .Z(o[2064]) );
  AND U26453 ( .A(p_input[2064]), .B(p_input[12064]), .Z(n17636) );
  AND U26454 ( .A(p_input[32064]), .B(p_input[22064]), .Z(n17635) );
  AND U26455 ( .A(n17637), .B(n17638), .Z(o[2063]) );
  AND U26456 ( .A(p_input[2063]), .B(p_input[12063]), .Z(n17638) );
  AND U26457 ( .A(p_input[32063]), .B(p_input[22063]), .Z(n17637) );
  AND U26458 ( .A(n17639), .B(n17640), .Z(o[2062]) );
  AND U26459 ( .A(p_input[2062]), .B(p_input[12062]), .Z(n17640) );
  AND U26460 ( .A(p_input[32062]), .B(p_input[22062]), .Z(n17639) );
  AND U26461 ( .A(n17641), .B(n17642), .Z(o[2061]) );
  AND U26462 ( .A(p_input[2061]), .B(p_input[12061]), .Z(n17642) );
  AND U26463 ( .A(p_input[32061]), .B(p_input[22061]), .Z(n17641) );
  AND U26464 ( .A(n17643), .B(n17644), .Z(o[2060]) );
  AND U26465 ( .A(p_input[2060]), .B(p_input[12060]), .Z(n17644) );
  AND U26466 ( .A(p_input[32060]), .B(p_input[22060]), .Z(n17643) );
  AND U26467 ( .A(n17645), .B(n17646), .Z(o[205]) );
  AND U26468 ( .A(p_input[20205]), .B(p_input[10205]), .Z(n17646) );
  AND U26469 ( .A(p_input[30205]), .B(p_input[205]), .Z(n17645) );
  AND U26470 ( .A(n17647), .B(n17648), .Z(o[2059]) );
  AND U26471 ( .A(p_input[2059]), .B(p_input[12059]), .Z(n17648) );
  AND U26472 ( .A(p_input[32059]), .B(p_input[22059]), .Z(n17647) );
  AND U26473 ( .A(n17649), .B(n17650), .Z(o[2058]) );
  AND U26474 ( .A(p_input[2058]), .B(p_input[12058]), .Z(n17650) );
  AND U26475 ( .A(p_input[32058]), .B(p_input[22058]), .Z(n17649) );
  AND U26476 ( .A(n17651), .B(n17652), .Z(o[2057]) );
  AND U26477 ( .A(p_input[2057]), .B(p_input[12057]), .Z(n17652) );
  AND U26478 ( .A(p_input[32057]), .B(p_input[22057]), .Z(n17651) );
  AND U26479 ( .A(n17653), .B(n17654), .Z(o[2056]) );
  AND U26480 ( .A(p_input[2056]), .B(p_input[12056]), .Z(n17654) );
  AND U26481 ( .A(p_input[32056]), .B(p_input[22056]), .Z(n17653) );
  AND U26482 ( .A(n17655), .B(n17656), .Z(o[2055]) );
  AND U26483 ( .A(p_input[2055]), .B(p_input[12055]), .Z(n17656) );
  AND U26484 ( .A(p_input[32055]), .B(p_input[22055]), .Z(n17655) );
  AND U26485 ( .A(n17657), .B(n17658), .Z(o[2054]) );
  AND U26486 ( .A(p_input[2054]), .B(p_input[12054]), .Z(n17658) );
  AND U26487 ( .A(p_input[32054]), .B(p_input[22054]), .Z(n17657) );
  AND U26488 ( .A(n17659), .B(n17660), .Z(o[2053]) );
  AND U26489 ( .A(p_input[2053]), .B(p_input[12053]), .Z(n17660) );
  AND U26490 ( .A(p_input[32053]), .B(p_input[22053]), .Z(n17659) );
  AND U26491 ( .A(n17661), .B(n17662), .Z(o[2052]) );
  AND U26492 ( .A(p_input[2052]), .B(p_input[12052]), .Z(n17662) );
  AND U26493 ( .A(p_input[32052]), .B(p_input[22052]), .Z(n17661) );
  AND U26494 ( .A(n17663), .B(n17664), .Z(o[2051]) );
  AND U26495 ( .A(p_input[2051]), .B(p_input[12051]), .Z(n17664) );
  AND U26496 ( .A(p_input[32051]), .B(p_input[22051]), .Z(n17663) );
  AND U26497 ( .A(n17665), .B(n17666), .Z(o[2050]) );
  AND U26498 ( .A(p_input[2050]), .B(p_input[12050]), .Z(n17666) );
  AND U26499 ( .A(p_input[32050]), .B(p_input[22050]), .Z(n17665) );
  AND U26500 ( .A(n17667), .B(n17668), .Z(o[204]) );
  AND U26501 ( .A(p_input[20204]), .B(p_input[10204]), .Z(n17668) );
  AND U26502 ( .A(p_input[30204]), .B(p_input[204]), .Z(n17667) );
  AND U26503 ( .A(n17669), .B(n17670), .Z(o[2049]) );
  AND U26504 ( .A(p_input[2049]), .B(p_input[12049]), .Z(n17670) );
  AND U26505 ( .A(p_input[32049]), .B(p_input[22049]), .Z(n17669) );
  AND U26506 ( .A(n17671), .B(n17672), .Z(o[2048]) );
  AND U26507 ( .A(p_input[2048]), .B(p_input[12048]), .Z(n17672) );
  AND U26508 ( .A(p_input[32048]), .B(p_input[22048]), .Z(n17671) );
  AND U26509 ( .A(n17673), .B(n17674), .Z(o[2047]) );
  AND U26510 ( .A(p_input[2047]), .B(p_input[12047]), .Z(n17674) );
  AND U26511 ( .A(p_input[32047]), .B(p_input[22047]), .Z(n17673) );
  AND U26512 ( .A(n17675), .B(n17676), .Z(o[2046]) );
  AND U26513 ( .A(p_input[2046]), .B(p_input[12046]), .Z(n17676) );
  AND U26514 ( .A(p_input[32046]), .B(p_input[22046]), .Z(n17675) );
  AND U26515 ( .A(n17677), .B(n17678), .Z(o[2045]) );
  AND U26516 ( .A(p_input[2045]), .B(p_input[12045]), .Z(n17678) );
  AND U26517 ( .A(p_input[32045]), .B(p_input[22045]), .Z(n17677) );
  AND U26518 ( .A(n17679), .B(n17680), .Z(o[2044]) );
  AND U26519 ( .A(p_input[2044]), .B(p_input[12044]), .Z(n17680) );
  AND U26520 ( .A(p_input[32044]), .B(p_input[22044]), .Z(n17679) );
  AND U26521 ( .A(n17681), .B(n17682), .Z(o[2043]) );
  AND U26522 ( .A(p_input[2043]), .B(p_input[12043]), .Z(n17682) );
  AND U26523 ( .A(p_input[32043]), .B(p_input[22043]), .Z(n17681) );
  AND U26524 ( .A(n17683), .B(n17684), .Z(o[2042]) );
  AND U26525 ( .A(p_input[2042]), .B(p_input[12042]), .Z(n17684) );
  AND U26526 ( .A(p_input[32042]), .B(p_input[22042]), .Z(n17683) );
  AND U26527 ( .A(n17685), .B(n17686), .Z(o[2041]) );
  AND U26528 ( .A(p_input[2041]), .B(p_input[12041]), .Z(n17686) );
  AND U26529 ( .A(p_input[32041]), .B(p_input[22041]), .Z(n17685) );
  AND U26530 ( .A(n17687), .B(n17688), .Z(o[2040]) );
  AND U26531 ( .A(p_input[2040]), .B(p_input[12040]), .Z(n17688) );
  AND U26532 ( .A(p_input[32040]), .B(p_input[22040]), .Z(n17687) );
  AND U26533 ( .A(n17689), .B(n17690), .Z(o[203]) );
  AND U26534 ( .A(p_input[20203]), .B(p_input[10203]), .Z(n17690) );
  AND U26535 ( .A(p_input[30203]), .B(p_input[203]), .Z(n17689) );
  AND U26536 ( .A(n17691), .B(n17692), .Z(o[2039]) );
  AND U26537 ( .A(p_input[2039]), .B(p_input[12039]), .Z(n17692) );
  AND U26538 ( .A(p_input[32039]), .B(p_input[22039]), .Z(n17691) );
  AND U26539 ( .A(n17693), .B(n17694), .Z(o[2038]) );
  AND U26540 ( .A(p_input[2038]), .B(p_input[12038]), .Z(n17694) );
  AND U26541 ( .A(p_input[32038]), .B(p_input[22038]), .Z(n17693) );
  AND U26542 ( .A(n17695), .B(n17696), .Z(o[2037]) );
  AND U26543 ( .A(p_input[2037]), .B(p_input[12037]), .Z(n17696) );
  AND U26544 ( .A(p_input[32037]), .B(p_input[22037]), .Z(n17695) );
  AND U26545 ( .A(n17697), .B(n17698), .Z(o[2036]) );
  AND U26546 ( .A(p_input[2036]), .B(p_input[12036]), .Z(n17698) );
  AND U26547 ( .A(p_input[32036]), .B(p_input[22036]), .Z(n17697) );
  AND U26548 ( .A(n17699), .B(n17700), .Z(o[2035]) );
  AND U26549 ( .A(p_input[2035]), .B(p_input[12035]), .Z(n17700) );
  AND U26550 ( .A(p_input[32035]), .B(p_input[22035]), .Z(n17699) );
  AND U26551 ( .A(n17701), .B(n17702), .Z(o[2034]) );
  AND U26552 ( .A(p_input[2034]), .B(p_input[12034]), .Z(n17702) );
  AND U26553 ( .A(p_input[32034]), .B(p_input[22034]), .Z(n17701) );
  AND U26554 ( .A(n17703), .B(n17704), .Z(o[2033]) );
  AND U26555 ( .A(p_input[2033]), .B(p_input[12033]), .Z(n17704) );
  AND U26556 ( .A(p_input[32033]), .B(p_input[22033]), .Z(n17703) );
  AND U26557 ( .A(n17705), .B(n17706), .Z(o[2032]) );
  AND U26558 ( .A(p_input[2032]), .B(p_input[12032]), .Z(n17706) );
  AND U26559 ( .A(p_input[32032]), .B(p_input[22032]), .Z(n17705) );
  AND U26560 ( .A(n17707), .B(n17708), .Z(o[2031]) );
  AND U26561 ( .A(p_input[2031]), .B(p_input[12031]), .Z(n17708) );
  AND U26562 ( .A(p_input[32031]), .B(p_input[22031]), .Z(n17707) );
  AND U26563 ( .A(n17709), .B(n17710), .Z(o[2030]) );
  AND U26564 ( .A(p_input[2030]), .B(p_input[12030]), .Z(n17710) );
  AND U26565 ( .A(p_input[32030]), .B(p_input[22030]), .Z(n17709) );
  AND U26566 ( .A(n17711), .B(n17712), .Z(o[202]) );
  AND U26567 ( .A(p_input[20202]), .B(p_input[10202]), .Z(n17712) );
  AND U26568 ( .A(p_input[30202]), .B(p_input[202]), .Z(n17711) );
  AND U26569 ( .A(n17713), .B(n17714), .Z(o[2029]) );
  AND U26570 ( .A(p_input[2029]), .B(p_input[12029]), .Z(n17714) );
  AND U26571 ( .A(p_input[32029]), .B(p_input[22029]), .Z(n17713) );
  AND U26572 ( .A(n17715), .B(n17716), .Z(o[2028]) );
  AND U26573 ( .A(p_input[2028]), .B(p_input[12028]), .Z(n17716) );
  AND U26574 ( .A(p_input[32028]), .B(p_input[22028]), .Z(n17715) );
  AND U26575 ( .A(n17717), .B(n17718), .Z(o[2027]) );
  AND U26576 ( .A(p_input[2027]), .B(p_input[12027]), .Z(n17718) );
  AND U26577 ( .A(p_input[32027]), .B(p_input[22027]), .Z(n17717) );
  AND U26578 ( .A(n17719), .B(n17720), .Z(o[2026]) );
  AND U26579 ( .A(p_input[2026]), .B(p_input[12026]), .Z(n17720) );
  AND U26580 ( .A(p_input[32026]), .B(p_input[22026]), .Z(n17719) );
  AND U26581 ( .A(n17721), .B(n17722), .Z(o[2025]) );
  AND U26582 ( .A(p_input[2025]), .B(p_input[12025]), .Z(n17722) );
  AND U26583 ( .A(p_input[32025]), .B(p_input[22025]), .Z(n17721) );
  AND U26584 ( .A(n17723), .B(n17724), .Z(o[2024]) );
  AND U26585 ( .A(p_input[2024]), .B(p_input[12024]), .Z(n17724) );
  AND U26586 ( .A(p_input[32024]), .B(p_input[22024]), .Z(n17723) );
  AND U26587 ( .A(n17725), .B(n17726), .Z(o[2023]) );
  AND U26588 ( .A(p_input[2023]), .B(p_input[12023]), .Z(n17726) );
  AND U26589 ( .A(p_input[32023]), .B(p_input[22023]), .Z(n17725) );
  AND U26590 ( .A(n17727), .B(n17728), .Z(o[2022]) );
  AND U26591 ( .A(p_input[2022]), .B(p_input[12022]), .Z(n17728) );
  AND U26592 ( .A(p_input[32022]), .B(p_input[22022]), .Z(n17727) );
  AND U26593 ( .A(n17729), .B(n17730), .Z(o[2021]) );
  AND U26594 ( .A(p_input[2021]), .B(p_input[12021]), .Z(n17730) );
  AND U26595 ( .A(p_input[32021]), .B(p_input[22021]), .Z(n17729) );
  AND U26596 ( .A(n17731), .B(n17732), .Z(o[2020]) );
  AND U26597 ( .A(p_input[2020]), .B(p_input[12020]), .Z(n17732) );
  AND U26598 ( .A(p_input[32020]), .B(p_input[22020]), .Z(n17731) );
  AND U26599 ( .A(n17733), .B(n17734), .Z(o[201]) );
  AND U26600 ( .A(p_input[201]), .B(p_input[10201]), .Z(n17734) );
  AND U26601 ( .A(p_input[30201]), .B(p_input[20201]), .Z(n17733) );
  AND U26602 ( .A(n17735), .B(n17736), .Z(o[2019]) );
  AND U26603 ( .A(p_input[2019]), .B(p_input[12019]), .Z(n17736) );
  AND U26604 ( .A(p_input[32019]), .B(p_input[22019]), .Z(n17735) );
  AND U26605 ( .A(n17737), .B(n17738), .Z(o[2018]) );
  AND U26606 ( .A(p_input[2018]), .B(p_input[12018]), .Z(n17738) );
  AND U26607 ( .A(p_input[32018]), .B(p_input[22018]), .Z(n17737) );
  AND U26608 ( .A(n17739), .B(n17740), .Z(o[2017]) );
  AND U26609 ( .A(p_input[2017]), .B(p_input[12017]), .Z(n17740) );
  AND U26610 ( .A(p_input[32017]), .B(p_input[22017]), .Z(n17739) );
  AND U26611 ( .A(n17741), .B(n17742), .Z(o[2016]) );
  AND U26612 ( .A(p_input[2016]), .B(p_input[12016]), .Z(n17742) );
  AND U26613 ( .A(p_input[32016]), .B(p_input[22016]), .Z(n17741) );
  AND U26614 ( .A(n17743), .B(n17744), .Z(o[2015]) );
  AND U26615 ( .A(p_input[2015]), .B(p_input[12015]), .Z(n17744) );
  AND U26616 ( .A(p_input[32015]), .B(p_input[22015]), .Z(n17743) );
  AND U26617 ( .A(n17745), .B(n17746), .Z(o[2014]) );
  AND U26618 ( .A(p_input[2014]), .B(p_input[12014]), .Z(n17746) );
  AND U26619 ( .A(p_input[32014]), .B(p_input[22014]), .Z(n17745) );
  AND U26620 ( .A(n17747), .B(n17748), .Z(o[2013]) );
  AND U26621 ( .A(p_input[2013]), .B(p_input[12013]), .Z(n17748) );
  AND U26622 ( .A(p_input[32013]), .B(p_input[22013]), .Z(n17747) );
  AND U26623 ( .A(n17749), .B(n17750), .Z(o[2012]) );
  AND U26624 ( .A(p_input[2012]), .B(p_input[12012]), .Z(n17750) );
  AND U26625 ( .A(p_input[32012]), .B(p_input[22012]), .Z(n17749) );
  AND U26626 ( .A(n17751), .B(n17752), .Z(o[2011]) );
  AND U26627 ( .A(p_input[2011]), .B(p_input[12011]), .Z(n17752) );
  AND U26628 ( .A(p_input[32011]), .B(p_input[22011]), .Z(n17751) );
  AND U26629 ( .A(n17753), .B(n17754), .Z(o[2010]) );
  AND U26630 ( .A(p_input[2010]), .B(p_input[12010]), .Z(n17754) );
  AND U26631 ( .A(p_input[32010]), .B(p_input[22010]), .Z(n17753) );
  AND U26632 ( .A(n17755), .B(n17756), .Z(o[200]) );
  AND U26633 ( .A(p_input[200]), .B(p_input[10200]), .Z(n17756) );
  AND U26634 ( .A(p_input[30200]), .B(p_input[20200]), .Z(n17755) );
  AND U26635 ( .A(n17757), .B(n17758), .Z(o[2009]) );
  AND U26636 ( .A(p_input[2009]), .B(p_input[12009]), .Z(n17758) );
  AND U26637 ( .A(p_input[32009]), .B(p_input[22009]), .Z(n17757) );
  AND U26638 ( .A(n17759), .B(n17760), .Z(o[2008]) );
  AND U26639 ( .A(p_input[2008]), .B(p_input[12008]), .Z(n17760) );
  AND U26640 ( .A(p_input[32008]), .B(p_input[22008]), .Z(n17759) );
  AND U26641 ( .A(n17761), .B(n17762), .Z(o[2007]) );
  AND U26642 ( .A(p_input[2007]), .B(p_input[12007]), .Z(n17762) );
  AND U26643 ( .A(p_input[32007]), .B(p_input[22007]), .Z(n17761) );
  AND U26644 ( .A(n17763), .B(n17764), .Z(o[2006]) );
  AND U26645 ( .A(p_input[2006]), .B(p_input[12006]), .Z(n17764) );
  AND U26646 ( .A(p_input[32006]), .B(p_input[22006]), .Z(n17763) );
  AND U26647 ( .A(n17765), .B(n17766), .Z(o[2005]) );
  AND U26648 ( .A(p_input[2005]), .B(p_input[12005]), .Z(n17766) );
  AND U26649 ( .A(p_input[32005]), .B(p_input[22005]), .Z(n17765) );
  AND U26650 ( .A(n17767), .B(n17768), .Z(o[2004]) );
  AND U26651 ( .A(p_input[2004]), .B(p_input[12004]), .Z(n17768) );
  AND U26652 ( .A(p_input[32004]), .B(p_input[22004]), .Z(n17767) );
  AND U26653 ( .A(n17769), .B(n17770), .Z(o[2003]) );
  AND U26654 ( .A(p_input[2003]), .B(p_input[12003]), .Z(n17770) );
  AND U26655 ( .A(p_input[32003]), .B(p_input[22003]), .Z(n17769) );
  AND U26656 ( .A(n17771), .B(n17772), .Z(o[2002]) );
  AND U26657 ( .A(p_input[2002]), .B(p_input[12002]), .Z(n17772) );
  AND U26658 ( .A(p_input[32002]), .B(p_input[22002]), .Z(n17771) );
  AND U26659 ( .A(n17773), .B(n17774), .Z(o[2001]) );
  AND U26660 ( .A(p_input[2001]), .B(p_input[12001]), .Z(n17774) );
  AND U26661 ( .A(p_input[32001]), .B(p_input[22001]), .Z(n17773) );
  AND U26662 ( .A(n17775), .B(n17776), .Z(o[2000]) );
  AND U26663 ( .A(p_input[2000]), .B(p_input[12000]), .Z(n17776) );
  AND U26664 ( .A(p_input[32000]), .B(p_input[22000]), .Z(n17775) );
  AND U26665 ( .A(n17777), .B(n17778), .Z(o[1]) );
  AND U26666 ( .A(p_input[1]), .B(p_input[10001]), .Z(n17778) );
  AND U26667 ( .A(p_input[30001]), .B(p_input[20001]), .Z(n17777) );
  AND U26668 ( .A(n17779), .B(n17780), .Z(o[19]) );
  AND U26669 ( .A(p_input[19]), .B(p_input[10019]), .Z(n17780) );
  AND U26670 ( .A(p_input[30019]), .B(p_input[20019]), .Z(n17779) );
  AND U26671 ( .A(n17781), .B(n17782), .Z(o[199]) );
  AND U26672 ( .A(p_input[199]), .B(p_input[10199]), .Z(n17782) );
  AND U26673 ( .A(p_input[30199]), .B(p_input[20199]), .Z(n17781) );
  AND U26674 ( .A(n17783), .B(n17784), .Z(o[1999]) );
  AND U26675 ( .A(p_input[1999]), .B(p_input[11999]), .Z(n17784) );
  AND U26676 ( .A(p_input[31999]), .B(p_input[21999]), .Z(n17783) );
  AND U26677 ( .A(n17785), .B(n17786), .Z(o[1998]) );
  AND U26678 ( .A(p_input[1998]), .B(p_input[11998]), .Z(n17786) );
  AND U26679 ( .A(p_input[31998]), .B(p_input[21998]), .Z(n17785) );
  AND U26680 ( .A(n17787), .B(n17788), .Z(o[1997]) );
  AND U26681 ( .A(p_input[1997]), .B(p_input[11997]), .Z(n17788) );
  AND U26682 ( .A(p_input[31997]), .B(p_input[21997]), .Z(n17787) );
  AND U26683 ( .A(n17789), .B(n17790), .Z(o[1996]) );
  AND U26684 ( .A(p_input[1996]), .B(p_input[11996]), .Z(n17790) );
  AND U26685 ( .A(p_input[31996]), .B(p_input[21996]), .Z(n17789) );
  AND U26686 ( .A(n17791), .B(n17792), .Z(o[1995]) );
  AND U26687 ( .A(p_input[1995]), .B(p_input[11995]), .Z(n17792) );
  AND U26688 ( .A(p_input[31995]), .B(p_input[21995]), .Z(n17791) );
  AND U26689 ( .A(n17793), .B(n17794), .Z(o[1994]) );
  AND U26690 ( .A(p_input[1994]), .B(p_input[11994]), .Z(n17794) );
  AND U26691 ( .A(p_input[31994]), .B(p_input[21994]), .Z(n17793) );
  AND U26692 ( .A(n17795), .B(n17796), .Z(o[1993]) );
  AND U26693 ( .A(p_input[1993]), .B(p_input[11993]), .Z(n17796) );
  AND U26694 ( .A(p_input[31993]), .B(p_input[21993]), .Z(n17795) );
  AND U26695 ( .A(n17797), .B(n17798), .Z(o[1992]) );
  AND U26696 ( .A(p_input[1992]), .B(p_input[11992]), .Z(n17798) );
  AND U26697 ( .A(p_input[31992]), .B(p_input[21992]), .Z(n17797) );
  AND U26698 ( .A(n17799), .B(n17800), .Z(o[1991]) );
  AND U26699 ( .A(p_input[1991]), .B(p_input[11991]), .Z(n17800) );
  AND U26700 ( .A(p_input[31991]), .B(p_input[21991]), .Z(n17799) );
  AND U26701 ( .A(n17801), .B(n17802), .Z(o[1990]) );
  AND U26702 ( .A(p_input[1990]), .B(p_input[11990]), .Z(n17802) );
  AND U26703 ( .A(p_input[31990]), .B(p_input[21990]), .Z(n17801) );
  AND U26704 ( .A(n17803), .B(n17804), .Z(o[198]) );
  AND U26705 ( .A(p_input[198]), .B(p_input[10198]), .Z(n17804) );
  AND U26706 ( .A(p_input[30198]), .B(p_input[20198]), .Z(n17803) );
  AND U26707 ( .A(n17805), .B(n17806), .Z(o[1989]) );
  AND U26708 ( .A(p_input[1989]), .B(p_input[11989]), .Z(n17806) );
  AND U26709 ( .A(p_input[31989]), .B(p_input[21989]), .Z(n17805) );
  AND U26710 ( .A(n17807), .B(n17808), .Z(o[1988]) );
  AND U26711 ( .A(p_input[1988]), .B(p_input[11988]), .Z(n17808) );
  AND U26712 ( .A(p_input[31988]), .B(p_input[21988]), .Z(n17807) );
  AND U26713 ( .A(n17809), .B(n17810), .Z(o[1987]) );
  AND U26714 ( .A(p_input[1987]), .B(p_input[11987]), .Z(n17810) );
  AND U26715 ( .A(p_input[31987]), .B(p_input[21987]), .Z(n17809) );
  AND U26716 ( .A(n17811), .B(n17812), .Z(o[1986]) );
  AND U26717 ( .A(p_input[1986]), .B(p_input[11986]), .Z(n17812) );
  AND U26718 ( .A(p_input[31986]), .B(p_input[21986]), .Z(n17811) );
  AND U26719 ( .A(n17813), .B(n17814), .Z(o[1985]) );
  AND U26720 ( .A(p_input[1985]), .B(p_input[11985]), .Z(n17814) );
  AND U26721 ( .A(p_input[31985]), .B(p_input[21985]), .Z(n17813) );
  AND U26722 ( .A(n17815), .B(n17816), .Z(o[1984]) );
  AND U26723 ( .A(p_input[1984]), .B(p_input[11984]), .Z(n17816) );
  AND U26724 ( .A(p_input[31984]), .B(p_input[21984]), .Z(n17815) );
  AND U26725 ( .A(n17817), .B(n17818), .Z(o[1983]) );
  AND U26726 ( .A(p_input[1983]), .B(p_input[11983]), .Z(n17818) );
  AND U26727 ( .A(p_input[31983]), .B(p_input[21983]), .Z(n17817) );
  AND U26728 ( .A(n17819), .B(n17820), .Z(o[1982]) );
  AND U26729 ( .A(p_input[1982]), .B(p_input[11982]), .Z(n17820) );
  AND U26730 ( .A(p_input[31982]), .B(p_input[21982]), .Z(n17819) );
  AND U26731 ( .A(n17821), .B(n17822), .Z(o[1981]) );
  AND U26732 ( .A(p_input[1981]), .B(p_input[11981]), .Z(n17822) );
  AND U26733 ( .A(p_input[31981]), .B(p_input[21981]), .Z(n17821) );
  AND U26734 ( .A(n17823), .B(n17824), .Z(o[1980]) );
  AND U26735 ( .A(p_input[1980]), .B(p_input[11980]), .Z(n17824) );
  AND U26736 ( .A(p_input[31980]), .B(p_input[21980]), .Z(n17823) );
  AND U26737 ( .A(n17825), .B(n17826), .Z(o[197]) );
  AND U26738 ( .A(p_input[197]), .B(p_input[10197]), .Z(n17826) );
  AND U26739 ( .A(p_input[30197]), .B(p_input[20197]), .Z(n17825) );
  AND U26740 ( .A(n17827), .B(n17828), .Z(o[1979]) );
  AND U26741 ( .A(p_input[1979]), .B(p_input[11979]), .Z(n17828) );
  AND U26742 ( .A(p_input[31979]), .B(p_input[21979]), .Z(n17827) );
  AND U26743 ( .A(n17829), .B(n17830), .Z(o[1978]) );
  AND U26744 ( .A(p_input[1978]), .B(p_input[11978]), .Z(n17830) );
  AND U26745 ( .A(p_input[31978]), .B(p_input[21978]), .Z(n17829) );
  AND U26746 ( .A(n17831), .B(n17832), .Z(o[1977]) );
  AND U26747 ( .A(p_input[1977]), .B(p_input[11977]), .Z(n17832) );
  AND U26748 ( .A(p_input[31977]), .B(p_input[21977]), .Z(n17831) );
  AND U26749 ( .A(n17833), .B(n17834), .Z(o[1976]) );
  AND U26750 ( .A(p_input[1976]), .B(p_input[11976]), .Z(n17834) );
  AND U26751 ( .A(p_input[31976]), .B(p_input[21976]), .Z(n17833) );
  AND U26752 ( .A(n17835), .B(n17836), .Z(o[1975]) );
  AND U26753 ( .A(p_input[1975]), .B(p_input[11975]), .Z(n17836) );
  AND U26754 ( .A(p_input[31975]), .B(p_input[21975]), .Z(n17835) );
  AND U26755 ( .A(n17837), .B(n17838), .Z(o[1974]) );
  AND U26756 ( .A(p_input[1974]), .B(p_input[11974]), .Z(n17838) );
  AND U26757 ( .A(p_input[31974]), .B(p_input[21974]), .Z(n17837) );
  AND U26758 ( .A(n17839), .B(n17840), .Z(o[1973]) );
  AND U26759 ( .A(p_input[1973]), .B(p_input[11973]), .Z(n17840) );
  AND U26760 ( .A(p_input[31973]), .B(p_input[21973]), .Z(n17839) );
  AND U26761 ( .A(n17841), .B(n17842), .Z(o[1972]) );
  AND U26762 ( .A(p_input[1972]), .B(p_input[11972]), .Z(n17842) );
  AND U26763 ( .A(p_input[31972]), .B(p_input[21972]), .Z(n17841) );
  AND U26764 ( .A(n17843), .B(n17844), .Z(o[1971]) );
  AND U26765 ( .A(p_input[1971]), .B(p_input[11971]), .Z(n17844) );
  AND U26766 ( .A(p_input[31971]), .B(p_input[21971]), .Z(n17843) );
  AND U26767 ( .A(n17845), .B(n17846), .Z(o[1970]) );
  AND U26768 ( .A(p_input[1970]), .B(p_input[11970]), .Z(n17846) );
  AND U26769 ( .A(p_input[31970]), .B(p_input[21970]), .Z(n17845) );
  AND U26770 ( .A(n17847), .B(n17848), .Z(o[196]) );
  AND U26771 ( .A(p_input[196]), .B(p_input[10196]), .Z(n17848) );
  AND U26772 ( .A(p_input[30196]), .B(p_input[20196]), .Z(n17847) );
  AND U26773 ( .A(n17849), .B(n17850), .Z(o[1969]) );
  AND U26774 ( .A(p_input[1969]), .B(p_input[11969]), .Z(n17850) );
  AND U26775 ( .A(p_input[31969]), .B(p_input[21969]), .Z(n17849) );
  AND U26776 ( .A(n17851), .B(n17852), .Z(o[1968]) );
  AND U26777 ( .A(p_input[1968]), .B(p_input[11968]), .Z(n17852) );
  AND U26778 ( .A(p_input[31968]), .B(p_input[21968]), .Z(n17851) );
  AND U26779 ( .A(n17853), .B(n17854), .Z(o[1967]) );
  AND U26780 ( .A(p_input[1967]), .B(p_input[11967]), .Z(n17854) );
  AND U26781 ( .A(p_input[31967]), .B(p_input[21967]), .Z(n17853) );
  AND U26782 ( .A(n17855), .B(n17856), .Z(o[1966]) );
  AND U26783 ( .A(p_input[1966]), .B(p_input[11966]), .Z(n17856) );
  AND U26784 ( .A(p_input[31966]), .B(p_input[21966]), .Z(n17855) );
  AND U26785 ( .A(n17857), .B(n17858), .Z(o[1965]) );
  AND U26786 ( .A(p_input[1965]), .B(p_input[11965]), .Z(n17858) );
  AND U26787 ( .A(p_input[31965]), .B(p_input[21965]), .Z(n17857) );
  AND U26788 ( .A(n17859), .B(n17860), .Z(o[1964]) );
  AND U26789 ( .A(p_input[1964]), .B(p_input[11964]), .Z(n17860) );
  AND U26790 ( .A(p_input[31964]), .B(p_input[21964]), .Z(n17859) );
  AND U26791 ( .A(n17861), .B(n17862), .Z(o[1963]) );
  AND U26792 ( .A(p_input[1963]), .B(p_input[11963]), .Z(n17862) );
  AND U26793 ( .A(p_input[31963]), .B(p_input[21963]), .Z(n17861) );
  AND U26794 ( .A(n17863), .B(n17864), .Z(o[1962]) );
  AND U26795 ( .A(p_input[1962]), .B(p_input[11962]), .Z(n17864) );
  AND U26796 ( .A(p_input[31962]), .B(p_input[21962]), .Z(n17863) );
  AND U26797 ( .A(n17865), .B(n17866), .Z(o[1961]) );
  AND U26798 ( .A(p_input[1961]), .B(p_input[11961]), .Z(n17866) );
  AND U26799 ( .A(p_input[31961]), .B(p_input[21961]), .Z(n17865) );
  AND U26800 ( .A(n17867), .B(n17868), .Z(o[1960]) );
  AND U26801 ( .A(p_input[1960]), .B(p_input[11960]), .Z(n17868) );
  AND U26802 ( .A(p_input[31960]), .B(p_input[21960]), .Z(n17867) );
  AND U26803 ( .A(n17869), .B(n17870), .Z(o[195]) );
  AND U26804 ( .A(p_input[195]), .B(p_input[10195]), .Z(n17870) );
  AND U26805 ( .A(p_input[30195]), .B(p_input[20195]), .Z(n17869) );
  AND U26806 ( .A(n17871), .B(n17872), .Z(o[1959]) );
  AND U26807 ( .A(p_input[1959]), .B(p_input[11959]), .Z(n17872) );
  AND U26808 ( .A(p_input[31959]), .B(p_input[21959]), .Z(n17871) );
  AND U26809 ( .A(n17873), .B(n17874), .Z(o[1958]) );
  AND U26810 ( .A(p_input[1958]), .B(p_input[11958]), .Z(n17874) );
  AND U26811 ( .A(p_input[31958]), .B(p_input[21958]), .Z(n17873) );
  AND U26812 ( .A(n17875), .B(n17876), .Z(o[1957]) );
  AND U26813 ( .A(p_input[1957]), .B(p_input[11957]), .Z(n17876) );
  AND U26814 ( .A(p_input[31957]), .B(p_input[21957]), .Z(n17875) );
  AND U26815 ( .A(n17877), .B(n17878), .Z(o[1956]) );
  AND U26816 ( .A(p_input[1956]), .B(p_input[11956]), .Z(n17878) );
  AND U26817 ( .A(p_input[31956]), .B(p_input[21956]), .Z(n17877) );
  AND U26818 ( .A(n17879), .B(n17880), .Z(o[1955]) );
  AND U26819 ( .A(p_input[1955]), .B(p_input[11955]), .Z(n17880) );
  AND U26820 ( .A(p_input[31955]), .B(p_input[21955]), .Z(n17879) );
  AND U26821 ( .A(n17881), .B(n17882), .Z(o[1954]) );
  AND U26822 ( .A(p_input[1954]), .B(p_input[11954]), .Z(n17882) );
  AND U26823 ( .A(p_input[31954]), .B(p_input[21954]), .Z(n17881) );
  AND U26824 ( .A(n17883), .B(n17884), .Z(o[1953]) );
  AND U26825 ( .A(p_input[1953]), .B(p_input[11953]), .Z(n17884) );
  AND U26826 ( .A(p_input[31953]), .B(p_input[21953]), .Z(n17883) );
  AND U26827 ( .A(n17885), .B(n17886), .Z(o[1952]) );
  AND U26828 ( .A(p_input[1952]), .B(p_input[11952]), .Z(n17886) );
  AND U26829 ( .A(p_input[31952]), .B(p_input[21952]), .Z(n17885) );
  AND U26830 ( .A(n17887), .B(n17888), .Z(o[1951]) );
  AND U26831 ( .A(p_input[1951]), .B(p_input[11951]), .Z(n17888) );
  AND U26832 ( .A(p_input[31951]), .B(p_input[21951]), .Z(n17887) );
  AND U26833 ( .A(n17889), .B(n17890), .Z(o[1950]) );
  AND U26834 ( .A(p_input[1950]), .B(p_input[11950]), .Z(n17890) );
  AND U26835 ( .A(p_input[31950]), .B(p_input[21950]), .Z(n17889) );
  AND U26836 ( .A(n17891), .B(n17892), .Z(o[194]) );
  AND U26837 ( .A(p_input[194]), .B(p_input[10194]), .Z(n17892) );
  AND U26838 ( .A(p_input[30194]), .B(p_input[20194]), .Z(n17891) );
  AND U26839 ( .A(n17893), .B(n17894), .Z(o[1949]) );
  AND U26840 ( .A(p_input[1949]), .B(p_input[11949]), .Z(n17894) );
  AND U26841 ( .A(p_input[31949]), .B(p_input[21949]), .Z(n17893) );
  AND U26842 ( .A(n17895), .B(n17896), .Z(o[1948]) );
  AND U26843 ( .A(p_input[1948]), .B(p_input[11948]), .Z(n17896) );
  AND U26844 ( .A(p_input[31948]), .B(p_input[21948]), .Z(n17895) );
  AND U26845 ( .A(n17897), .B(n17898), .Z(o[1947]) );
  AND U26846 ( .A(p_input[1947]), .B(p_input[11947]), .Z(n17898) );
  AND U26847 ( .A(p_input[31947]), .B(p_input[21947]), .Z(n17897) );
  AND U26848 ( .A(n17899), .B(n17900), .Z(o[1946]) );
  AND U26849 ( .A(p_input[1946]), .B(p_input[11946]), .Z(n17900) );
  AND U26850 ( .A(p_input[31946]), .B(p_input[21946]), .Z(n17899) );
  AND U26851 ( .A(n17901), .B(n17902), .Z(o[1945]) );
  AND U26852 ( .A(p_input[1945]), .B(p_input[11945]), .Z(n17902) );
  AND U26853 ( .A(p_input[31945]), .B(p_input[21945]), .Z(n17901) );
  AND U26854 ( .A(n17903), .B(n17904), .Z(o[1944]) );
  AND U26855 ( .A(p_input[1944]), .B(p_input[11944]), .Z(n17904) );
  AND U26856 ( .A(p_input[31944]), .B(p_input[21944]), .Z(n17903) );
  AND U26857 ( .A(n17905), .B(n17906), .Z(o[1943]) );
  AND U26858 ( .A(p_input[1943]), .B(p_input[11943]), .Z(n17906) );
  AND U26859 ( .A(p_input[31943]), .B(p_input[21943]), .Z(n17905) );
  AND U26860 ( .A(n17907), .B(n17908), .Z(o[1942]) );
  AND U26861 ( .A(p_input[1942]), .B(p_input[11942]), .Z(n17908) );
  AND U26862 ( .A(p_input[31942]), .B(p_input[21942]), .Z(n17907) );
  AND U26863 ( .A(n17909), .B(n17910), .Z(o[1941]) );
  AND U26864 ( .A(p_input[1941]), .B(p_input[11941]), .Z(n17910) );
  AND U26865 ( .A(p_input[31941]), .B(p_input[21941]), .Z(n17909) );
  AND U26866 ( .A(n17911), .B(n17912), .Z(o[1940]) );
  AND U26867 ( .A(p_input[1940]), .B(p_input[11940]), .Z(n17912) );
  AND U26868 ( .A(p_input[31940]), .B(p_input[21940]), .Z(n17911) );
  AND U26869 ( .A(n17913), .B(n17914), .Z(o[193]) );
  AND U26870 ( .A(p_input[193]), .B(p_input[10193]), .Z(n17914) );
  AND U26871 ( .A(p_input[30193]), .B(p_input[20193]), .Z(n17913) );
  AND U26872 ( .A(n17915), .B(n17916), .Z(o[1939]) );
  AND U26873 ( .A(p_input[1939]), .B(p_input[11939]), .Z(n17916) );
  AND U26874 ( .A(p_input[31939]), .B(p_input[21939]), .Z(n17915) );
  AND U26875 ( .A(n17917), .B(n17918), .Z(o[1938]) );
  AND U26876 ( .A(p_input[1938]), .B(p_input[11938]), .Z(n17918) );
  AND U26877 ( .A(p_input[31938]), .B(p_input[21938]), .Z(n17917) );
  AND U26878 ( .A(n17919), .B(n17920), .Z(o[1937]) );
  AND U26879 ( .A(p_input[1937]), .B(p_input[11937]), .Z(n17920) );
  AND U26880 ( .A(p_input[31937]), .B(p_input[21937]), .Z(n17919) );
  AND U26881 ( .A(n17921), .B(n17922), .Z(o[1936]) );
  AND U26882 ( .A(p_input[1936]), .B(p_input[11936]), .Z(n17922) );
  AND U26883 ( .A(p_input[31936]), .B(p_input[21936]), .Z(n17921) );
  AND U26884 ( .A(n17923), .B(n17924), .Z(o[1935]) );
  AND U26885 ( .A(p_input[1935]), .B(p_input[11935]), .Z(n17924) );
  AND U26886 ( .A(p_input[31935]), .B(p_input[21935]), .Z(n17923) );
  AND U26887 ( .A(n17925), .B(n17926), .Z(o[1934]) );
  AND U26888 ( .A(p_input[1934]), .B(p_input[11934]), .Z(n17926) );
  AND U26889 ( .A(p_input[31934]), .B(p_input[21934]), .Z(n17925) );
  AND U26890 ( .A(n17927), .B(n17928), .Z(o[1933]) );
  AND U26891 ( .A(p_input[1933]), .B(p_input[11933]), .Z(n17928) );
  AND U26892 ( .A(p_input[31933]), .B(p_input[21933]), .Z(n17927) );
  AND U26893 ( .A(n17929), .B(n17930), .Z(o[1932]) );
  AND U26894 ( .A(p_input[1932]), .B(p_input[11932]), .Z(n17930) );
  AND U26895 ( .A(p_input[31932]), .B(p_input[21932]), .Z(n17929) );
  AND U26896 ( .A(n17931), .B(n17932), .Z(o[1931]) );
  AND U26897 ( .A(p_input[1931]), .B(p_input[11931]), .Z(n17932) );
  AND U26898 ( .A(p_input[31931]), .B(p_input[21931]), .Z(n17931) );
  AND U26899 ( .A(n17933), .B(n17934), .Z(o[1930]) );
  AND U26900 ( .A(p_input[1930]), .B(p_input[11930]), .Z(n17934) );
  AND U26901 ( .A(p_input[31930]), .B(p_input[21930]), .Z(n17933) );
  AND U26902 ( .A(n17935), .B(n17936), .Z(o[192]) );
  AND U26903 ( .A(p_input[192]), .B(p_input[10192]), .Z(n17936) );
  AND U26904 ( .A(p_input[30192]), .B(p_input[20192]), .Z(n17935) );
  AND U26905 ( .A(n17937), .B(n17938), .Z(o[1929]) );
  AND U26906 ( .A(p_input[1929]), .B(p_input[11929]), .Z(n17938) );
  AND U26907 ( .A(p_input[31929]), .B(p_input[21929]), .Z(n17937) );
  AND U26908 ( .A(n17939), .B(n17940), .Z(o[1928]) );
  AND U26909 ( .A(p_input[1928]), .B(p_input[11928]), .Z(n17940) );
  AND U26910 ( .A(p_input[31928]), .B(p_input[21928]), .Z(n17939) );
  AND U26911 ( .A(n17941), .B(n17942), .Z(o[1927]) );
  AND U26912 ( .A(p_input[1927]), .B(p_input[11927]), .Z(n17942) );
  AND U26913 ( .A(p_input[31927]), .B(p_input[21927]), .Z(n17941) );
  AND U26914 ( .A(n17943), .B(n17944), .Z(o[1926]) );
  AND U26915 ( .A(p_input[1926]), .B(p_input[11926]), .Z(n17944) );
  AND U26916 ( .A(p_input[31926]), .B(p_input[21926]), .Z(n17943) );
  AND U26917 ( .A(n17945), .B(n17946), .Z(o[1925]) );
  AND U26918 ( .A(p_input[1925]), .B(p_input[11925]), .Z(n17946) );
  AND U26919 ( .A(p_input[31925]), .B(p_input[21925]), .Z(n17945) );
  AND U26920 ( .A(n17947), .B(n17948), .Z(o[1924]) );
  AND U26921 ( .A(p_input[1924]), .B(p_input[11924]), .Z(n17948) );
  AND U26922 ( .A(p_input[31924]), .B(p_input[21924]), .Z(n17947) );
  AND U26923 ( .A(n17949), .B(n17950), .Z(o[1923]) );
  AND U26924 ( .A(p_input[1923]), .B(p_input[11923]), .Z(n17950) );
  AND U26925 ( .A(p_input[31923]), .B(p_input[21923]), .Z(n17949) );
  AND U26926 ( .A(n17951), .B(n17952), .Z(o[1922]) );
  AND U26927 ( .A(p_input[1922]), .B(p_input[11922]), .Z(n17952) );
  AND U26928 ( .A(p_input[31922]), .B(p_input[21922]), .Z(n17951) );
  AND U26929 ( .A(n17953), .B(n17954), .Z(o[1921]) );
  AND U26930 ( .A(p_input[1921]), .B(p_input[11921]), .Z(n17954) );
  AND U26931 ( .A(p_input[31921]), .B(p_input[21921]), .Z(n17953) );
  AND U26932 ( .A(n17955), .B(n17956), .Z(o[1920]) );
  AND U26933 ( .A(p_input[1920]), .B(p_input[11920]), .Z(n17956) );
  AND U26934 ( .A(p_input[31920]), .B(p_input[21920]), .Z(n17955) );
  AND U26935 ( .A(n17957), .B(n17958), .Z(o[191]) );
  AND U26936 ( .A(p_input[191]), .B(p_input[10191]), .Z(n17958) );
  AND U26937 ( .A(p_input[30191]), .B(p_input[20191]), .Z(n17957) );
  AND U26938 ( .A(n17959), .B(n17960), .Z(o[1919]) );
  AND U26939 ( .A(p_input[1919]), .B(p_input[11919]), .Z(n17960) );
  AND U26940 ( .A(p_input[31919]), .B(p_input[21919]), .Z(n17959) );
  AND U26941 ( .A(n17961), .B(n17962), .Z(o[1918]) );
  AND U26942 ( .A(p_input[1918]), .B(p_input[11918]), .Z(n17962) );
  AND U26943 ( .A(p_input[31918]), .B(p_input[21918]), .Z(n17961) );
  AND U26944 ( .A(n17963), .B(n17964), .Z(o[1917]) );
  AND U26945 ( .A(p_input[1917]), .B(p_input[11917]), .Z(n17964) );
  AND U26946 ( .A(p_input[31917]), .B(p_input[21917]), .Z(n17963) );
  AND U26947 ( .A(n17965), .B(n17966), .Z(o[1916]) );
  AND U26948 ( .A(p_input[1916]), .B(p_input[11916]), .Z(n17966) );
  AND U26949 ( .A(p_input[31916]), .B(p_input[21916]), .Z(n17965) );
  AND U26950 ( .A(n17967), .B(n17968), .Z(o[1915]) );
  AND U26951 ( .A(p_input[1915]), .B(p_input[11915]), .Z(n17968) );
  AND U26952 ( .A(p_input[31915]), .B(p_input[21915]), .Z(n17967) );
  AND U26953 ( .A(n17969), .B(n17970), .Z(o[1914]) );
  AND U26954 ( .A(p_input[1914]), .B(p_input[11914]), .Z(n17970) );
  AND U26955 ( .A(p_input[31914]), .B(p_input[21914]), .Z(n17969) );
  AND U26956 ( .A(n17971), .B(n17972), .Z(o[1913]) );
  AND U26957 ( .A(p_input[1913]), .B(p_input[11913]), .Z(n17972) );
  AND U26958 ( .A(p_input[31913]), .B(p_input[21913]), .Z(n17971) );
  AND U26959 ( .A(n17973), .B(n17974), .Z(o[1912]) );
  AND U26960 ( .A(p_input[1912]), .B(p_input[11912]), .Z(n17974) );
  AND U26961 ( .A(p_input[31912]), .B(p_input[21912]), .Z(n17973) );
  AND U26962 ( .A(n17975), .B(n17976), .Z(o[1911]) );
  AND U26963 ( .A(p_input[1911]), .B(p_input[11911]), .Z(n17976) );
  AND U26964 ( .A(p_input[31911]), .B(p_input[21911]), .Z(n17975) );
  AND U26965 ( .A(n17977), .B(n17978), .Z(o[1910]) );
  AND U26966 ( .A(p_input[1910]), .B(p_input[11910]), .Z(n17978) );
  AND U26967 ( .A(p_input[31910]), .B(p_input[21910]), .Z(n17977) );
  AND U26968 ( .A(n17979), .B(n17980), .Z(o[190]) );
  AND U26969 ( .A(p_input[190]), .B(p_input[10190]), .Z(n17980) );
  AND U26970 ( .A(p_input[30190]), .B(p_input[20190]), .Z(n17979) );
  AND U26971 ( .A(n17981), .B(n17982), .Z(o[1909]) );
  AND U26972 ( .A(p_input[1909]), .B(p_input[11909]), .Z(n17982) );
  AND U26973 ( .A(p_input[31909]), .B(p_input[21909]), .Z(n17981) );
  AND U26974 ( .A(n17983), .B(n17984), .Z(o[1908]) );
  AND U26975 ( .A(p_input[1908]), .B(p_input[11908]), .Z(n17984) );
  AND U26976 ( .A(p_input[31908]), .B(p_input[21908]), .Z(n17983) );
  AND U26977 ( .A(n17985), .B(n17986), .Z(o[1907]) );
  AND U26978 ( .A(p_input[1907]), .B(p_input[11907]), .Z(n17986) );
  AND U26979 ( .A(p_input[31907]), .B(p_input[21907]), .Z(n17985) );
  AND U26980 ( .A(n17987), .B(n17988), .Z(o[1906]) );
  AND U26981 ( .A(p_input[1906]), .B(p_input[11906]), .Z(n17988) );
  AND U26982 ( .A(p_input[31906]), .B(p_input[21906]), .Z(n17987) );
  AND U26983 ( .A(n17989), .B(n17990), .Z(o[1905]) );
  AND U26984 ( .A(p_input[1905]), .B(p_input[11905]), .Z(n17990) );
  AND U26985 ( .A(p_input[31905]), .B(p_input[21905]), .Z(n17989) );
  AND U26986 ( .A(n17991), .B(n17992), .Z(o[1904]) );
  AND U26987 ( .A(p_input[1904]), .B(p_input[11904]), .Z(n17992) );
  AND U26988 ( .A(p_input[31904]), .B(p_input[21904]), .Z(n17991) );
  AND U26989 ( .A(n17993), .B(n17994), .Z(o[1903]) );
  AND U26990 ( .A(p_input[1903]), .B(p_input[11903]), .Z(n17994) );
  AND U26991 ( .A(p_input[31903]), .B(p_input[21903]), .Z(n17993) );
  AND U26992 ( .A(n17995), .B(n17996), .Z(o[1902]) );
  AND U26993 ( .A(p_input[1902]), .B(p_input[11902]), .Z(n17996) );
  AND U26994 ( .A(p_input[31902]), .B(p_input[21902]), .Z(n17995) );
  AND U26995 ( .A(n17997), .B(n17998), .Z(o[1901]) );
  AND U26996 ( .A(p_input[1901]), .B(p_input[11901]), .Z(n17998) );
  AND U26997 ( .A(p_input[31901]), .B(p_input[21901]), .Z(n17997) );
  AND U26998 ( .A(n17999), .B(n18000), .Z(o[1900]) );
  AND U26999 ( .A(p_input[1900]), .B(p_input[11900]), .Z(n18000) );
  AND U27000 ( .A(p_input[31900]), .B(p_input[21900]), .Z(n17999) );
  AND U27001 ( .A(n18001), .B(n18002), .Z(o[18]) );
  AND U27002 ( .A(p_input[18]), .B(p_input[10018]), .Z(n18002) );
  AND U27003 ( .A(p_input[30018]), .B(p_input[20018]), .Z(n18001) );
  AND U27004 ( .A(n18003), .B(n18004), .Z(o[189]) );
  AND U27005 ( .A(p_input[189]), .B(p_input[10189]), .Z(n18004) );
  AND U27006 ( .A(p_input[30189]), .B(p_input[20189]), .Z(n18003) );
  AND U27007 ( .A(n18005), .B(n18006), .Z(o[1899]) );
  AND U27008 ( .A(p_input[1899]), .B(p_input[11899]), .Z(n18006) );
  AND U27009 ( .A(p_input[31899]), .B(p_input[21899]), .Z(n18005) );
  AND U27010 ( .A(n18007), .B(n18008), .Z(o[1898]) );
  AND U27011 ( .A(p_input[1898]), .B(p_input[11898]), .Z(n18008) );
  AND U27012 ( .A(p_input[31898]), .B(p_input[21898]), .Z(n18007) );
  AND U27013 ( .A(n18009), .B(n18010), .Z(o[1897]) );
  AND U27014 ( .A(p_input[1897]), .B(p_input[11897]), .Z(n18010) );
  AND U27015 ( .A(p_input[31897]), .B(p_input[21897]), .Z(n18009) );
  AND U27016 ( .A(n18011), .B(n18012), .Z(o[1896]) );
  AND U27017 ( .A(p_input[1896]), .B(p_input[11896]), .Z(n18012) );
  AND U27018 ( .A(p_input[31896]), .B(p_input[21896]), .Z(n18011) );
  AND U27019 ( .A(n18013), .B(n18014), .Z(o[1895]) );
  AND U27020 ( .A(p_input[1895]), .B(p_input[11895]), .Z(n18014) );
  AND U27021 ( .A(p_input[31895]), .B(p_input[21895]), .Z(n18013) );
  AND U27022 ( .A(n18015), .B(n18016), .Z(o[1894]) );
  AND U27023 ( .A(p_input[1894]), .B(p_input[11894]), .Z(n18016) );
  AND U27024 ( .A(p_input[31894]), .B(p_input[21894]), .Z(n18015) );
  AND U27025 ( .A(n18017), .B(n18018), .Z(o[1893]) );
  AND U27026 ( .A(p_input[1893]), .B(p_input[11893]), .Z(n18018) );
  AND U27027 ( .A(p_input[31893]), .B(p_input[21893]), .Z(n18017) );
  AND U27028 ( .A(n18019), .B(n18020), .Z(o[1892]) );
  AND U27029 ( .A(p_input[1892]), .B(p_input[11892]), .Z(n18020) );
  AND U27030 ( .A(p_input[31892]), .B(p_input[21892]), .Z(n18019) );
  AND U27031 ( .A(n18021), .B(n18022), .Z(o[1891]) );
  AND U27032 ( .A(p_input[1891]), .B(p_input[11891]), .Z(n18022) );
  AND U27033 ( .A(p_input[31891]), .B(p_input[21891]), .Z(n18021) );
  AND U27034 ( .A(n18023), .B(n18024), .Z(o[1890]) );
  AND U27035 ( .A(p_input[1890]), .B(p_input[11890]), .Z(n18024) );
  AND U27036 ( .A(p_input[31890]), .B(p_input[21890]), .Z(n18023) );
  AND U27037 ( .A(n18025), .B(n18026), .Z(o[188]) );
  AND U27038 ( .A(p_input[188]), .B(p_input[10188]), .Z(n18026) );
  AND U27039 ( .A(p_input[30188]), .B(p_input[20188]), .Z(n18025) );
  AND U27040 ( .A(n18027), .B(n18028), .Z(o[1889]) );
  AND U27041 ( .A(p_input[1889]), .B(p_input[11889]), .Z(n18028) );
  AND U27042 ( .A(p_input[31889]), .B(p_input[21889]), .Z(n18027) );
  AND U27043 ( .A(n18029), .B(n18030), .Z(o[1888]) );
  AND U27044 ( .A(p_input[1888]), .B(p_input[11888]), .Z(n18030) );
  AND U27045 ( .A(p_input[31888]), .B(p_input[21888]), .Z(n18029) );
  AND U27046 ( .A(n18031), .B(n18032), .Z(o[1887]) );
  AND U27047 ( .A(p_input[1887]), .B(p_input[11887]), .Z(n18032) );
  AND U27048 ( .A(p_input[31887]), .B(p_input[21887]), .Z(n18031) );
  AND U27049 ( .A(n18033), .B(n18034), .Z(o[1886]) );
  AND U27050 ( .A(p_input[1886]), .B(p_input[11886]), .Z(n18034) );
  AND U27051 ( .A(p_input[31886]), .B(p_input[21886]), .Z(n18033) );
  AND U27052 ( .A(n18035), .B(n18036), .Z(o[1885]) );
  AND U27053 ( .A(p_input[1885]), .B(p_input[11885]), .Z(n18036) );
  AND U27054 ( .A(p_input[31885]), .B(p_input[21885]), .Z(n18035) );
  AND U27055 ( .A(n18037), .B(n18038), .Z(o[1884]) );
  AND U27056 ( .A(p_input[1884]), .B(p_input[11884]), .Z(n18038) );
  AND U27057 ( .A(p_input[31884]), .B(p_input[21884]), .Z(n18037) );
  AND U27058 ( .A(n18039), .B(n18040), .Z(o[1883]) );
  AND U27059 ( .A(p_input[1883]), .B(p_input[11883]), .Z(n18040) );
  AND U27060 ( .A(p_input[31883]), .B(p_input[21883]), .Z(n18039) );
  AND U27061 ( .A(n18041), .B(n18042), .Z(o[1882]) );
  AND U27062 ( .A(p_input[1882]), .B(p_input[11882]), .Z(n18042) );
  AND U27063 ( .A(p_input[31882]), .B(p_input[21882]), .Z(n18041) );
  AND U27064 ( .A(n18043), .B(n18044), .Z(o[1881]) );
  AND U27065 ( .A(p_input[1881]), .B(p_input[11881]), .Z(n18044) );
  AND U27066 ( .A(p_input[31881]), .B(p_input[21881]), .Z(n18043) );
  AND U27067 ( .A(n18045), .B(n18046), .Z(o[1880]) );
  AND U27068 ( .A(p_input[1880]), .B(p_input[11880]), .Z(n18046) );
  AND U27069 ( .A(p_input[31880]), .B(p_input[21880]), .Z(n18045) );
  AND U27070 ( .A(n18047), .B(n18048), .Z(o[187]) );
  AND U27071 ( .A(p_input[187]), .B(p_input[10187]), .Z(n18048) );
  AND U27072 ( .A(p_input[30187]), .B(p_input[20187]), .Z(n18047) );
  AND U27073 ( .A(n18049), .B(n18050), .Z(o[1879]) );
  AND U27074 ( .A(p_input[1879]), .B(p_input[11879]), .Z(n18050) );
  AND U27075 ( .A(p_input[31879]), .B(p_input[21879]), .Z(n18049) );
  AND U27076 ( .A(n18051), .B(n18052), .Z(o[1878]) );
  AND U27077 ( .A(p_input[1878]), .B(p_input[11878]), .Z(n18052) );
  AND U27078 ( .A(p_input[31878]), .B(p_input[21878]), .Z(n18051) );
  AND U27079 ( .A(n18053), .B(n18054), .Z(o[1877]) );
  AND U27080 ( .A(p_input[1877]), .B(p_input[11877]), .Z(n18054) );
  AND U27081 ( .A(p_input[31877]), .B(p_input[21877]), .Z(n18053) );
  AND U27082 ( .A(n18055), .B(n18056), .Z(o[1876]) );
  AND U27083 ( .A(p_input[1876]), .B(p_input[11876]), .Z(n18056) );
  AND U27084 ( .A(p_input[31876]), .B(p_input[21876]), .Z(n18055) );
  AND U27085 ( .A(n18057), .B(n18058), .Z(o[1875]) );
  AND U27086 ( .A(p_input[1875]), .B(p_input[11875]), .Z(n18058) );
  AND U27087 ( .A(p_input[31875]), .B(p_input[21875]), .Z(n18057) );
  AND U27088 ( .A(n18059), .B(n18060), .Z(o[1874]) );
  AND U27089 ( .A(p_input[1874]), .B(p_input[11874]), .Z(n18060) );
  AND U27090 ( .A(p_input[31874]), .B(p_input[21874]), .Z(n18059) );
  AND U27091 ( .A(n18061), .B(n18062), .Z(o[1873]) );
  AND U27092 ( .A(p_input[1873]), .B(p_input[11873]), .Z(n18062) );
  AND U27093 ( .A(p_input[31873]), .B(p_input[21873]), .Z(n18061) );
  AND U27094 ( .A(n18063), .B(n18064), .Z(o[1872]) );
  AND U27095 ( .A(p_input[1872]), .B(p_input[11872]), .Z(n18064) );
  AND U27096 ( .A(p_input[31872]), .B(p_input[21872]), .Z(n18063) );
  AND U27097 ( .A(n18065), .B(n18066), .Z(o[1871]) );
  AND U27098 ( .A(p_input[1871]), .B(p_input[11871]), .Z(n18066) );
  AND U27099 ( .A(p_input[31871]), .B(p_input[21871]), .Z(n18065) );
  AND U27100 ( .A(n18067), .B(n18068), .Z(o[1870]) );
  AND U27101 ( .A(p_input[1870]), .B(p_input[11870]), .Z(n18068) );
  AND U27102 ( .A(p_input[31870]), .B(p_input[21870]), .Z(n18067) );
  AND U27103 ( .A(n18069), .B(n18070), .Z(o[186]) );
  AND U27104 ( .A(p_input[186]), .B(p_input[10186]), .Z(n18070) );
  AND U27105 ( .A(p_input[30186]), .B(p_input[20186]), .Z(n18069) );
  AND U27106 ( .A(n18071), .B(n18072), .Z(o[1869]) );
  AND U27107 ( .A(p_input[1869]), .B(p_input[11869]), .Z(n18072) );
  AND U27108 ( .A(p_input[31869]), .B(p_input[21869]), .Z(n18071) );
  AND U27109 ( .A(n18073), .B(n18074), .Z(o[1868]) );
  AND U27110 ( .A(p_input[1868]), .B(p_input[11868]), .Z(n18074) );
  AND U27111 ( .A(p_input[31868]), .B(p_input[21868]), .Z(n18073) );
  AND U27112 ( .A(n18075), .B(n18076), .Z(o[1867]) );
  AND U27113 ( .A(p_input[1867]), .B(p_input[11867]), .Z(n18076) );
  AND U27114 ( .A(p_input[31867]), .B(p_input[21867]), .Z(n18075) );
  AND U27115 ( .A(n18077), .B(n18078), .Z(o[1866]) );
  AND U27116 ( .A(p_input[1866]), .B(p_input[11866]), .Z(n18078) );
  AND U27117 ( .A(p_input[31866]), .B(p_input[21866]), .Z(n18077) );
  AND U27118 ( .A(n18079), .B(n18080), .Z(o[1865]) );
  AND U27119 ( .A(p_input[1865]), .B(p_input[11865]), .Z(n18080) );
  AND U27120 ( .A(p_input[31865]), .B(p_input[21865]), .Z(n18079) );
  AND U27121 ( .A(n18081), .B(n18082), .Z(o[1864]) );
  AND U27122 ( .A(p_input[1864]), .B(p_input[11864]), .Z(n18082) );
  AND U27123 ( .A(p_input[31864]), .B(p_input[21864]), .Z(n18081) );
  AND U27124 ( .A(n18083), .B(n18084), .Z(o[1863]) );
  AND U27125 ( .A(p_input[1863]), .B(p_input[11863]), .Z(n18084) );
  AND U27126 ( .A(p_input[31863]), .B(p_input[21863]), .Z(n18083) );
  AND U27127 ( .A(n18085), .B(n18086), .Z(o[1862]) );
  AND U27128 ( .A(p_input[1862]), .B(p_input[11862]), .Z(n18086) );
  AND U27129 ( .A(p_input[31862]), .B(p_input[21862]), .Z(n18085) );
  AND U27130 ( .A(n18087), .B(n18088), .Z(o[1861]) );
  AND U27131 ( .A(p_input[1861]), .B(p_input[11861]), .Z(n18088) );
  AND U27132 ( .A(p_input[31861]), .B(p_input[21861]), .Z(n18087) );
  AND U27133 ( .A(n18089), .B(n18090), .Z(o[1860]) );
  AND U27134 ( .A(p_input[1860]), .B(p_input[11860]), .Z(n18090) );
  AND U27135 ( .A(p_input[31860]), .B(p_input[21860]), .Z(n18089) );
  AND U27136 ( .A(n18091), .B(n18092), .Z(o[185]) );
  AND U27137 ( .A(p_input[185]), .B(p_input[10185]), .Z(n18092) );
  AND U27138 ( .A(p_input[30185]), .B(p_input[20185]), .Z(n18091) );
  AND U27139 ( .A(n18093), .B(n18094), .Z(o[1859]) );
  AND U27140 ( .A(p_input[1859]), .B(p_input[11859]), .Z(n18094) );
  AND U27141 ( .A(p_input[31859]), .B(p_input[21859]), .Z(n18093) );
  AND U27142 ( .A(n18095), .B(n18096), .Z(o[1858]) );
  AND U27143 ( .A(p_input[1858]), .B(p_input[11858]), .Z(n18096) );
  AND U27144 ( .A(p_input[31858]), .B(p_input[21858]), .Z(n18095) );
  AND U27145 ( .A(n18097), .B(n18098), .Z(o[1857]) );
  AND U27146 ( .A(p_input[1857]), .B(p_input[11857]), .Z(n18098) );
  AND U27147 ( .A(p_input[31857]), .B(p_input[21857]), .Z(n18097) );
  AND U27148 ( .A(n18099), .B(n18100), .Z(o[1856]) );
  AND U27149 ( .A(p_input[1856]), .B(p_input[11856]), .Z(n18100) );
  AND U27150 ( .A(p_input[31856]), .B(p_input[21856]), .Z(n18099) );
  AND U27151 ( .A(n18101), .B(n18102), .Z(o[1855]) );
  AND U27152 ( .A(p_input[1855]), .B(p_input[11855]), .Z(n18102) );
  AND U27153 ( .A(p_input[31855]), .B(p_input[21855]), .Z(n18101) );
  AND U27154 ( .A(n18103), .B(n18104), .Z(o[1854]) );
  AND U27155 ( .A(p_input[1854]), .B(p_input[11854]), .Z(n18104) );
  AND U27156 ( .A(p_input[31854]), .B(p_input[21854]), .Z(n18103) );
  AND U27157 ( .A(n18105), .B(n18106), .Z(o[1853]) );
  AND U27158 ( .A(p_input[1853]), .B(p_input[11853]), .Z(n18106) );
  AND U27159 ( .A(p_input[31853]), .B(p_input[21853]), .Z(n18105) );
  AND U27160 ( .A(n18107), .B(n18108), .Z(o[1852]) );
  AND U27161 ( .A(p_input[1852]), .B(p_input[11852]), .Z(n18108) );
  AND U27162 ( .A(p_input[31852]), .B(p_input[21852]), .Z(n18107) );
  AND U27163 ( .A(n18109), .B(n18110), .Z(o[1851]) );
  AND U27164 ( .A(p_input[1851]), .B(p_input[11851]), .Z(n18110) );
  AND U27165 ( .A(p_input[31851]), .B(p_input[21851]), .Z(n18109) );
  AND U27166 ( .A(n18111), .B(n18112), .Z(o[1850]) );
  AND U27167 ( .A(p_input[1850]), .B(p_input[11850]), .Z(n18112) );
  AND U27168 ( .A(p_input[31850]), .B(p_input[21850]), .Z(n18111) );
  AND U27169 ( .A(n18113), .B(n18114), .Z(o[184]) );
  AND U27170 ( .A(p_input[184]), .B(p_input[10184]), .Z(n18114) );
  AND U27171 ( .A(p_input[30184]), .B(p_input[20184]), .Z(n18113) );
  AND U27172 ( .A(n18115), .B(n18116), .Z(o[1849]) );
  AND U27173 ( .A(p_input[1849]), .B(p_input[11849]), .Z(n18116) );
  AND U27174 ( .A(p_input[31849]), .B(p_input[21849]), .Z(n18115) );
  AND U27175 ( .A(n18117), .B(n18118), .Z(o[1848]) );
  AND U27176 ( .A(p_input[1848]), .B(p_input[11848]), .Z(n18118) );
  AND U27177 ( .A(p_input[31848]), .B(p_input[21848]), .Z(n18117) );
  AND U27178 ( .A(n18119), .B(n18120), .Z(o[1847]) );
  AND U27179 ( .A(p_input[1847]), .B(p_input[11847]), .Z(n18120) );
  AND U27180 ( .A(p_input[31847]), .B(p_input[21847]), .Z(n18119) );
  AND U27181 ( .A(n18121), .B(n18122), .Z(o[1846]) );
  AND U27182 ( .A(p_input[1846]), .B(p_input[11846]), .Z(n18122) );
  AND U27183 ( .A(p_input[31846]), .B(p_input[21846]), .Z(n18121) );
  AND U27184 ( .A(n18123), .B(n18124), .Z(o[1845]) );
  AND U27185 ( .A(p_input[1845]), .B(p_input[11845]), .Z(n18124) );
  AND U27186 ( .A(p_input[31845]), .B(p_input[21845]), .Z(n18123) );
  AND U27187 ( .A(n18125), .B(n18126), .Z(o[1844]) );
  AND U27188 ( .A(p_input[1844]), .B(p_input[11844]), .Z(n18126) );
  AND U27189 ( .A(p_input[31844]), .B(p_input[21844]), .Z(n18125) );
  AND U27190 ( .A(n18127), .B(n18128), .Z(o[1843]) );
  AND U27191 ( .A(p_input[1843]), .B(p_input[11843]), .Z(n18128) );
  AND U27192 ( .A(p_input[31843]), .B(p_input[21843]), .Z(n18127) );
  AND U27193 ( .A(n18129), .B(n18130), .Z(o[1842]) );
  AND U27194 ( .A(p_input[1842]), .B(p_input[11842]), .Z(n18130) );
  AND U27195 ( .A(p_input[31842]), .B(p_input[21842]), .Z(n18129) );
  AND U27196 ( .A(n18131), .B(n18132), .Z(o[1841]) );
  AND U27197 ( .A(p_input[1841]), .B(p_input[11841]), .Z(n18132) );
  AND U27198 ( .A(p_input[31841]), .B(p_input[21841]), .Z(n18131) );
  AND U27199 ( .A(n18133), .B(n18134), .Z(o[1840]) );
  AND U27200 ( .A(p_input[1840]), .B(p_input[11840]), .Z(n18134) );
  AND U27201 ( .A(p_input[31840]), .B(p_input[21840]), .Z(n18133) );
  AND U27202 ( .A(n18135), .B(n18136), .Z(o[183]) );
  AND U27203 ( .A(p_input[183]), .B(p_input[10183]), .Z(n18136) );
  AND U27204 ( .A(p_input[30183]), .B(p_input[20183]), .Z(n18135) );
  AND U27205 ( .A(n18137), .B(n18138), .Z(o[1839]) );
  AND U27206 ( .A(p_input[1839]), .B(p_input[11839]), .Z(n18138) );
  AND U27207 ( .A(p_input[31839]), .B(p_input[21839]), .Z(n18137) );
  AND U27208 ( .A(n18139), .B(n18140), .Z(o[1838]) );
  AND U27209 ( .A(p_input[1838]), .B(p_input[11838]), .Z(n18140) );
  AND U27210 ( .A(p_input[31838]), .B(p_input[21838]), .Z(n18139) );
  AND U27211 ( .A(n18141), .B(n18142), .Z(o[1837]) );
  AND U27212 ( .A(p_input[1837]), .B(p_input[11837]), .Z(n18142) );
  AND U27213 ( .A(p_input[31837]), .B(p_input[21837]), .Z(n18141) );
  AND U27214 ( .A(n18143), .B(n18144), .Z(o[1836]) );
  AND U27215 ( .A(p_input[1836]), .B(p_input[11836]), .Z(n18144) );
  AND U27216 ( .A(p_input[31836]), .B(p_input[21836]), .Z(n18143) );
  AND U27217 ( .A(n18145), .B(n18146), .Z(o[1835]) );
  AND U27218 ( .A(p_input[1835]), .B(p_input[11835]), .Z(n18146) );
  AND U27219 ( .A(p_input[31835]), .B(p_input[21835]), .Z(n18145) );
  AND U27220 ( .A(n18147), .B(n18148), .Z(o[1834]) );
  AND U27221 ( .A(p_input[1834]), .B(p_input[11834]), .Z(n18148) );
  AND U27222 ( .A(p_input[31834]), .B(p_input[21834]), .Z(n18147) );
  AND U27223 ( .A(n18149), .B(n18150), .Z(o[1833]) );
  AND U27224 ( .A(p_input[1833]), .B(p_input[11833]), .Z(n18150) );
  AND U27225 ( .A(p_input[31833]), .B(p_input[21833]), .Z(n18149) );
  AND U27226 ( .A(n18151), .B(n18152), .Z(o[1832]) );
  AND U27227 ( .A(p_input[1832]), .B(p_input[11832]), .Z(n18152) );
  AND U27228 ( .A(p_input[31832]), .B(p_input[21832]), .Z(n18151) );
  AND U27229 ( .A(n18153), .B(n18154), .Z(o[1831]) );
  AND U27230 ( .A(p_input[1831]), .B(p_input[11831]), .Z(n18154) );
  AND U27231 ( .A(p_input[31831]), .B(p_input[21831]), .Z(n18153) );
  AND U27232 ( .A(n18155), .B(n18156), .Z(o[1830]) );
  AND U27233 ( .A(p_input[1830]), .B(p_input[11830]), .Z(n18156) );
  AND U27234 ( .A(p_input[31830]), .B(p_input[21830]), .Z(n18155) );
  AND U27235 ( .A(n18157), .B(n18158), .Z(o[182]) );
  AND U27236 ( .A(p_input[182]), .B(p_input[10182]), .Z(n18158) );
  AND U27237 ( .A(p_input[30182]), .B(p_input[20182]), .Z(n18157) );
  AND U27238 ( .A(n18159), .B(n18160), .Z(o[1829]) );
  AND U27239 ( .A(p_input[1829]), .B(p_input[11829]), .Z(n18160) );
  AND U27240 ( .A(p_input[31829]), .B(p_input[21829]), .Z(n18159) );
  AND U27241 ( .A(n18161), .B(n18162), .Z(o[1828]) );
  AND U27242 ( .A(p_input[1828]), .B(p_input[11828]), .Z(n18162) );
  AND U27243 ( .A(p_input[31828]), .B(p_input[21828]), .Z(n18161) );
  AND U27244 ( .A(n18163), .B(n18164), .Z(o[1827]) );
  AND U27245 ( .A(p_input[1827]), .B(p_input[11827]), .Z(n18164) );
  AND U27246 ( .A(p_input[31827]), .B(p_input[21827]), .Z(n18163) );
  AND U27247 ( .A(n18165), .B(n18166), .Z(o[1826]) );
  AND U27248 ( .A(p_input[1826]), .B(p_input[11826]), .Z(n18166) );
  AND U27249 ( .A(p_input[31826]), .B(p_input[21826]), .Z(n18165) );
  AND U27250 ( .A(n18167), .B(n18168), .Z(o[1825]) );
  AND U27251 ( .A(p_input[1825]), .B(p_input[11825]), .Z(n18168) );
  AND U27252 ( .A(p_input[31825]), .B(p_input[21825]), .Z(n18167) );
  AND U27253 ( .A(n18169), .B(n18170), .Z(o[1824]) );
  AND U27254 ( .A(p_input[1824]), .B(p_input[11824]), .Z(n18170) );
  AND U27255 ( .A(p_input[31824]), .B(p_input[21824]), .Z(n18169) );
  AND U27256 ( .A(n18171), .B(n18172), .Z(o[1823]) );
  AND U27257 ( .A(p_input[1823]), .B(p_input[11823]), .Z(n18172) );
  AND U27258 ( .A(p_input[31823]), .B(p_input[21823]), .Z(n18171) );
  AND U27259 ( .A(n18173), .B(n18174), .Z(o[1822]) );
  AND U27260 ( .A(p_input[1822]), .B(p_input[11822]), .Z(n18174) );
  AND U27261 ( .A(p_input[31822]), .B(p_input[21822]), .Z(n18173) );
  AND U27262 ( .A(n18175), .B(n18176), .Z(o[1821]) );
  AND U27263 ( .A(p_input[1821]), .B(p_input[11821]), .Z(n18176) );
  AND U27264 ( .A(p_input[31821]), .B(p_input[21821]), .Z(n18175) );
  AND U27265 ( .A(n18177), .B(n18178), .Z(o[1820]) );
  AND U27266 ( .A(p_input[1820]), .B(p_input[11820]), .Z(n18178) );
  AND U27267 ( .A(p_input[31820]), .B(p_input[21820]), .Z(n18177) );
  AND U27268 ( .A(n18179), .B(n18180), .Z(o[181]) );
  AND U27269 ( .A(p_input[181]), .B(p_input[10181]), .Z(n18180) );
  AND U27270 ( .A(p_input[30181]), .B(p_input[20181]), .Z(n18179) );
  AND U27271 ( .A(n18181), .B(n18182), .Z(o[1819]) );
  AND U27272 ( .A(p_input[1819]), .B(p_input[11819]), .Z(n18182) );
  AND U27273 ( .A(p_input[31819]), .B(p_input[21819]), .Z(n18181) );
  AND U27274 ( .A(n18183), .B(n18184), .Z(o[1818]) );
  AND U27275 ( .A(p_input[1818]), .B(p_input[11818]), .Z(n18184) );
  AND U27276 ( .A(p_input[31818]), .B(p_input[21818]), .Z(n18183) );
  AND U27277 ( .A(n18185), .B(n18186), .Z(o[1817]) );
  AND U27278 ( .A(p_input[1817]), .B(p_input[11817]), .Z(n18186) );
  AND U27279 ( .A(p_input[31817]), .B(p_input[21817]), .Z(n18185) );
  AND U27280 ( .A(n18187), .B(n18188), .Z(o[1816]) );
  AND U27281 ( .A(p_input[1816]), .B(p_input[11816]), .Z(n18188) );
  AND U27282 ( .A(p_input[31816]), .B(p_input[21816]), .Z(n18187) );
  AND U27283 ( .A(n18189), .B(n18190), .Z(o[1815]) );
  AND U27284 ( .A(p_input[1815]), .B(p_input[11815]), .Z(n18190) );
  AND U27285 ( .A(p_input[31815]), .B(p_input[21815]), .Z(n18189) );
  AND U27286 ( .A(n18191), .B(n18192), .Z(o[1814]) );
  AND U27287 ( .A(p_input[1814]), .B(p_input[11814]), .Z(n18192) );
  AND U27288 ( .A(p_input[31814]), .B(p_input[21814]), .Z(n18191) );
  AND U27289 ( .A(n18193), .B(n18194), .Z(o[1813]) );
  AND U27290 ( .A(p_input[1813]), .B(p_input[11813]), .Z(n18194) );
  AND U27291 ( .A(p_input[31813]), .B(p_input[21813]), .Z(n18193) );
  AND U27292 ( .A(n18195), .B(n18196), .Z(o[1812]) );
  AND U27293 ( .A(p_input[1812]), .B(p_input[11812]), .Z(n18196) );
  AND U27294 ( .A(p_input[31812]), .B(p_input[21812]), .Z(n18195) );
  AND U27295 ( .A(n18197), .B(n18198), .Z(o[1811]) );
  AND U27296 ( .A(p_input[1811]), .B(p_input[11811]), .Z(n18198) );
  AND U27297 ( .A(p_input[31811]), .B(p_input[21811]), .Z(n18197) );
  AND U27298 ( .A(n18199), .B(n18200), .Z(o[1810]) );
  AND U27299 ( .A(p_input[1810]), .B(p_input[11810]), .Z(n18200) );
  AND U27300 ( .A(p_input[31810]), .B(p_input[21810]), .Z(n18199) );
  AND U27301 ( .A(n18201), .B(n18202), .Z(o[180]) );
  AND U27302 ( .A(p_input[180]), .B(p_input[10180]), .Z(n18202) );
  AND U27303 ( .A(p_input[30180]), .B(p_input[20180]), .Z(n18201) );
  AND U27304 ( .A(n18203), .B(n18204), .Z(o[1809]) );
  AND U27305 ( .A(p_input[1809]), .B(p_input[11809]), .Z(n18204) );
  AND U27306 ( .A(p_input[31809]), .B(p_input[21809]), .Z(n18203) );
  AND U27307 ( .A(n18205), .B(n18206), .Z(o[1808]) );
  AND U27308 ( .A(p_input[1808]), .B(p_input[11808]), .Z(n18206) );
  AND U27309 ( .A(p_input[31808]), .B(p_input[21808]), .Z(n18205) );
  AND U27310 ( .A(n18207), .B(n18208), .Z(o[1807]) );
  AND U27311 ( .A(p_input[1807]), .B(p_input[11807]), .Z(n18208) );
  AND U27312 ( .A(p_input[31807]), .B(p_input[21807]), .Z(n18207) );
  AND U27313 ( .A(n18209), .B(n18210), .Z(o[1806]) );
  AND U27314 ( .A(p_input[1806]), .B(p_input[11806]), .Z(n18210) );
  AND U27315 ( .A(p_input[31806]), .B(p_input[21806]), .Z(n18209) );
  AND U27316 ( .A(n18211), .B(n18212), .Z(o[1805]) );
  AND U27317 ( .A(p_input[1805]), .B(p_input[11805]), .Z(n18212) );
  AND U27318 ( .A(p_input[31805]), .B(p_input[21805]), .Z(n18211) );
  AND U27319 ( .A(n18213), .B(n18214), .Z(o[1804]) );
  AND U27320 ( .A(p_input[1804]), .B(p_input[11804]), .Z(n18214) );
  AND U27321 ( .A(p_input[31804]), .B(p_input[21804]), .Z(n18213) );
  AND U27322 ( .A(n18215), .B(n18216), .Z(o[1803]) );
  AND U27323 ( .A(p_input[1803]), .B(p_input[11803]), .Z(n18216) );
  AND U27324 ( .A(p_input[31803]), .B(p_input[21803]), .Z(n18215) );
  AND U27325 ( .A(n18217), .B(n18218), .Z(o[1802]) );
  AND U27326 ( .A(p_input[1802]), .B(p_input[11802]), .Z(n18218) );
  AND U27327 ( .A(p_input[31802]), .B(p_input[21802]), .Z(n18217) );
  AND U27328 ( .A(n18219), .B(n18220), .Z(o[1801]) );
  AND U27329 ( .A(p_input[1801]), .B(p_input[11801]), .Z(n18220) );
  AND U27330 ( .A(p_input[31801]), .B(p_input[21801]), .Z(n18219) );
  AND U27331 ( .A(n18221), .B(n18222), .Z(o[1800]) );
  AND U27332 ( .A(p_input[1800]), .B(p_input[11800]), .Z(n18222) );
  AND U27333 ( .A(p_input[31800]), .B(p_input[21800]), .Z(n18221) );
  AND U27334 ( .A(n18223), .B(n18224), .Z(o[17]) );
  AND U27335 ( .A(p_input[17]), .B(p_input[10017]), .Z(n18224) );
  AND U27336 ( .A(p_input[30017]), .B(p_input[20017]), .Z(n18223) );
  AND U27337 ( .A(n18225), .B(n18226), .Z(o[179]) );
  AND U27338 ( .A(p_input[179]), .B(p_input[10179]), .Z(n18226) );
  AND U27339 ( .A(p_input[30179]), .B(p_input[20179]), .Z(n18225) );
  AND U27340 ( .A(n18227), .B(n18228), .Z(o[1799]) );
  AND U27341 ( .A(p_input[1799]), .B(p_input[11799]), .Z(n18228) );
  AND U27342 ( .A(p_input[31799]), .B(p_input[21799]), .Z(n18227) );
  AND U27343 ( .A(n18229), .B(n18230), .Z(o[1798]) );
  AND U27344 ( .A(p_input[1798]), .B(p_input[11798]), .Z(n18230) );
  AND U27345 ( .A(p_input[31798]), .B(p_input[21798]), .Z(n18229) );
  AND U27346 ( .A(n18231), .B(n18232), .Z(o[1797]) );
  AND U27347 ( .A(p_input[1797]), .B(p_input[11797]), .Z(n18232) );
  AND U27348 ( .A(p_input[31797]), .B(p_input[21797]), .Z(n18231) );
  AND U27349 ( .A(n18233), .B(n18234), .Z(o[1796]) );
  AND U27350 ( .A(p_input[1796]), .B(p_input[11796]), .Z(n18234) );
  AND U27351 ( .A(p_input[31796]), .B(p_input[21796]), .Z(n18233) );
  AND U27352 ( .A(n18235), .B(n18236), .Z(o[1795]) );
  AND U27353 ( .A(p_input[1795]), .B(p_input[11795]), .Z(n18236) );
  AND U27354 ( .A(p_input[31795]), .B(p_input[21795]), .Z(n18235) );
  AND U27355 ( .A(n18237), .B(n18238), .Z(o[1794]) );
  AND U27356 ( .A(p_input[1794]), .B(p_input[11794]), .Z(n18238) );
  AND U27357 ( .A(p_input[31794]), .B(p_input[21794]), .Z(n18237) );
  AND U27358 ( .A(n18239), .B(n18240), .Z(o[1793]) );
  AND U27359 ( .A(p_input[1793]), .B(p_input[11793]), .Z(n18240) );
  AND U27360 ( .A(p_input[31793]), .B(p_input[21793]), .Z(n18239) );
  AND U27361 ( .A(n18241), .B(n18242), .Z(o[1792]) );
  AND U27362 ( .A(p_input[1792]), .B(p_input[11792]), .Z(n18242) );
  AND U27363 ( .A(p_input[31792]), .B(p_input[21792]), .Z(n18241) );
  AND U27364 ( .A(n18243), .B(n18244), .Z(o[1791]) );
  AND U27365 ( .A(p_input[1791]), .B(p_input[11791]), .Z(n18244) );
  AND U27366 ( .A(p_input[31791]), .B(p_input[21791]), .Z(n18243) );
  AND U27367 ( .A(n18245), .B(n18246), .Z(o[1790]) );
  AND U27368 ( .A(p_input[1790]), .B(p_input[11790]), .Z(n18246) );
  AND U27369 ( .A(p_input[31790]), .B(p_input[21790]), .Z(n18245) );
  AND U27370 ( .A(n18247), .B(n18248), .Z(o[178]) );
  AND U27371 ( .A(p_input[178]), .B(p_input[10178]), .Z(n18248) );
  AND U27372 ( .A(p_input[30178]), .B(p_input[20178]), .Z(n18247) );
  AND U27373 ( .A(n18249), .B(n18250), .Z(o[1789]) );
  AND U27374 ( .A(p_input[1789]), .B(p_input[11789]), .Z(n18250) );
  AND U27375 ( .A(p_input[31789]), .B(p_input[21789]), .Z(n18249) );
  AND U27376 ( .A(n18251), .B(n18252), .Z(o[1788]) );
  AND U27377 ( .A(p_input[1788]), .B(p_input[11788]), .Z(n18252) );
  AND U27378 ( .A(p_input[31788]), .B(p_input[21788]), .Z(n18251) );
  AND U27379 ( .A(n18253), .B(n18254), .Z(o[1787]) );
  AND U27380 ( .A(p_input[1787]), .B(p_input[11787]), .Z(n18254) );
  AND U27381 ( .A(p_input[31787]), .B(p_input[21787]), .Z(n18253) );
  AND U27382 ( .A(n18255), .B(n18256), .Z(o[1786]) );
  AND U27383 ( .A(p_input[1786]), .B(p_input[11786]), .Z(n18256) );
  AND U27384 ( .A(p_input[31786]), .B(p_input[21786]), .Z(n18255) );
  AND U27385 ( .A(n18257), .B(n18258), .Z(o[1785]) );
  AND U27386 ( .A(p_input[1785]), .B(p_input[11785]), .Z(n18258) );
  AND U27387 ( .A(p_input[31785]), .B(p_input[21785]), .Z(n18257) );
  AND U27388 ( .A(n18259), .B(n18260), .Z(o[1784]) );
  AND U27389 ( .A(p_input[1784]), .B(p_input[11784]), .Z(n18260) );
  AND U27390 ( .A(p_input[31784]), .B(p_input[21784]), .Z(n18259) );
  AND U27391 ( .A(n18261), .B(n18262), .Z(o[1783]) );
  AND U27392 ( .A(p_input[1783]), .B(p_input[11783]), .Z(n18262) );
  AND U27393 ( .A(p_input[31783]), .B(p_input[21783]), .Z(n18261) );
  AND U27394 ( .A(n18263), .B(n18264), .Z(o[1782]) );
  AND U27395 ( .A(p_input[1782]), .B(p_input[11782]), .Z(n18264) );
  AND U27396 ( .A(p_input[31782]), .B(p_input[21782]), .Z(n18263) );
  AND U27397 ( .A(n18265), .B(n18266), .Z(o[1781]) );
  AND U27398 ( .A(p_input[1781]), .B(p_input[11781]), .Z(n18266) );
  AND U27399 ( .A(p_input[31781]), .B(p_input[21781]), .Z(n18265) );
  AND U27400 ( .A(n18267), .B(n18268), .Z(o[1780]) );
  AND U27401 ( .A(p_input[1780]), .B(p_input[11780]), .Z(n18268) );
  AND U27402 ( .A(p_input[31780]), .B(p_input[21780]), .Z(n18267) );
  AND U27403 ( .A(n18269), .B(n18270), .Z(o[177]) );
  AND U27404 ( .A(p_input[177]), .B(p_input[10177]), .Z(n18270) );
  AND U27405 ( .A(p_input[30177]), .B(p_input[20177]), .Z(n18269) );
  AND U27406 ( .A(n18271), .B(n18272), .Z(o[1779]) );
  AND U27407 ( .A(p_input[1779]), .B(p_input[11779]), .Z(n18272) );
  AND U27408 ( .A(p_input[31779]), .B(p_input[21779]), .Z(n18271) );
  AND U27409 ( .A(n18273), .B(n18274), .Z(o[1778]) );
  AND U27410 ( .A(p_input[1778]), .B(p_input[11778]), .Z(n18274) );
  AND U27411 ( .A(p_input[31778]), .B(p_input[21778]), .Z(n18273) );
  AND U27412 ( .A(n18275), .B(n18276), .Z(o[1777]) );
  AND U27413 ( .A(p_input[1777]), .B(p_input[11777]), .Z(n18276) );
  AND U27414 ( .A(p_input[31777]), .B(p_input[21777]), .Z(n18275) );
  AND U27415 ( .A(n18277), .B(n18278), .Z(o[1776]) );
  AND U27416 ( .A(p_input[1776]), .B(p_input[11776]), .Z(n18278) );
  AND U27417 ( .A(p_input[31776]), .B(p_input[21776]), .Z(n18277) );
  AND U27418 ( .A(n18279), .B(n18280), .Z(o[1775]) );
  AND U27419 ( .A(p_input[1775]), .B(p_input[11775]), .Z(n18280) );
  AND U27420 ( .A(p_input[31775]), .B(p_input[21775]), .Z(n18279) );
  AND U27421 ( .A(n18281), .B(n18282), .Z(o[1774]) );
  AND U27422 ( .A(p_input[1774]), .B(p_input[11774]), .Z(n18282) );
  AND U27423 ( .A(p_input[31774]), .B(p_input[21774]), .Z(n18281) );
  AND U27424 ( .A(n18283), .B(n18284), .Z(o[1773]) );
  AND U27425 ( .A(p_input[1773]), .B(p_input[11773]), .Z(n18284) );
  AND U27426 ( .A(p_input[31773]), .B(p_input[21773]), .Z(n18283) );
  AND U27427 ( .A(n18285), .B(n18286), .Z(o[1772]) );
  AND U27428 ( .A(p_input[1772]), .B(p_input[11772]), .Z(n18286) );
  AND U27429 ( .A(p_input[31772]), .B(p_input[21772]), .Z(n18285) );
  AND U27430 ( .A(n18287), .B(n18288), .Z(o[1771]) );
  AND U27431 ( .A(p_input[1771]), .B(p_input[11771]), .Z(n18288) );
  AND U27432 ( .A(p_input[31771]), .B(p_input[21771]), .Z(n18287) );
  AND U27433 ( .A(n18289), .B(n18290), .Z(o[1770]) );
  AND U27434 ( .A(p_input[1770]), .B(p_input[11770]), .Z(n18290) );
  AND U27435 ( .A(p_input[31770]), .B(p_input[21770]), .Z(n18289) );
  AND U27436 ( .A(n18291), .B(n18292), .Z(o[176]) );
  AND U27437 ( .A(p_input[176]), .B(p_input[10176]), .Z(n18292) );
  AND U27438 ( .A(p_input[30176]), .B(p_input[20176]), .Z(n18291) );
  AND U27439 ( .A(n18293), .B(n18294), .Z(o[1769]) );
  AND U27440 ( .A(p_input[1769]), .B(p_input[11769]), .Z(n18294) );
  AND U27441 ( .A(p_input[31769]), .B(p_input[21769]), .Z(n18293) );
  AND U27442 ( .A(n18295), .B(n18296), .Z(o[1768]) );
  AND U27443 ( .A(p_input[1768]), .B(p_input[11768]), .Z(n18296) );
  AND U27444 ( .A(p_input[31768]), .B(p_input[21768]), .Z(n18295) );
  AND U27445 ( .A(n18297), .B(n18298), .Z(o[1767]) );
  AND U27446 ( .A(p_input[1767]), .B(p_input[11767]), .Z(n18298) );
  AND U27447 ( .A(p_input[31767]), .B(p_input[21767]), .Z(n18297) );
  AND U27448 ( .A(n18299), .B(n18300), .Z(o[1766]) );
  AND U27449 ( .A(p_input[1766]), .B(p_input[11766]), .Z(n18300) );
  AND U27450 ( .A(p_input[31766]), .B(p_input[21766]), .Z(n18299) );
  AND U27451 ( .A(n18301), .B(n18302), .Z(o[1765]) );
  AND U27452 ( .A(p_input[1765]), .B(p_input[11765]), .Z(n18302) );
  AND U27453 ( .A(p_input[31765]), .B(p_input[21765]), .Z(n18301) );
  AND U27454 ( .A(n18303), .B(n18304), .Z(o[1764]) );
  AND U27455 ( .A(p_input[1764]), .B(p_input[11764]), .Z(n18304) );
  AND U27456 ( .A(p_input[31764]), .B(p_input[21764]), .Z(n18303) );
  AND U27457 ( .A(n18305), .B(n18306), .Z(o[1763]) );
  AND U27458 ( .A(p_input[1763]), .B(p_input[11763]), .Z(n18306) );
  AND U27459 ( .A(p_input[31763]), .B(p_input[21763]), .Z(n18305) );
  AND U27460 ( .A(n18307), .B(n18308), .Z(o[1762]) );
  AND U27461 ( .A(p_input[1762]), .B(p_input[11762]), .Z(n18308) );
  AND U27462 ( .A(p_input[31762]), .B(p_input[21762]), .Z(n18307) );
  AND U27463 ( .A(n18309), .B(n18310), .Z(o[1761]) );
  AND U27464 ( .A(p_input[1761]), .B(p_input[11761]), .Z(n18310) );
  AND U27465 ( .A(p_input[31761]), .B(p_input[21761]), .Z(n18309) );
  AND U27466 ( .A(n18311), .B(n18312), .Z(o[1760]) );
  AND U27467 ( .A(p_input[1760]), .B(p_input[11760]), .Z(n18312) );
  AND U27468 ( .A(p_input[31760]), .B(p_input[21760]), .Z(n18311) );
  AND U27469 ( .A(n18313), .B(n18314), .Z(o[175]) );
  AND U27470 ( .A(p_input[175]), .B(p_input[10175]), .Z(n18314) );
  AND U27471 ( .A(p_input[30175]), .B(p_input[20175]), .Z(n18313) );
  AND U27472 ( .A(n18315), .B(n18316), .Z(o[1759]) );
  AND U27473 ( .A(p_input[1759]), .B(p_input[11759]), .Z(n18316) );
  AND U27474 ( .A(p_input[31759]), .B(p_input[21759]), .Z(n18315) );
  AND U27475 ( .A(n18317), .B(n18318), .Z(o[1758]) );
  AND U27476 ( .A(p_input[1758]), .B(p_input[11758]), .Z(n18318) );
  AND U27477 ( .A(p_input[31758]), .B(p_input[21758]), .Z(n18317) );
  AND U27478 ( .A(n18319), .B(n18320), .Z(o[1757]) );
  AND U27479 ( .A(p_input[1757]), .B(p_input[11757]), .Z(n18320) );
  AND U27480 ( .A(p_input[31757]), .B(p_input[21757]), .Z(n18319) );
  AND U27481 ( .A(n18321), .B(n18322), .Z(o[1756]) );
  AND U27482 ( .A(p_input[1756]), .B(p_input[11756]), .Z(n18322) );
  AND U27483 ( .A(p_input[31756]), .B(p_input[21756]), .Z(n18321) );
  AND U27484 ( .A(n18323), .B(n18324), .Z(o[1755]) );
  AND U27485 ( .A(p_input[1755]), .B(p_input[11755]), .Z(n18324) );
  AND U27486 ( .A(p_input[31755]), .B(p_input[21755]), .Z(n18323) );
  AND U27487 ( .A(n18325), .B(n18326), .Z(o[1754]) );
  AND U27488 ( .A(p_input[1754]), .B(p_input[11754]), .Z(n18326) );
  AND U27489 ( .A(p_input[31754]), .B(p_input[21754]), .Z(n18325) );
  AND U27490 ( .A(n18327), .B(n18328), .Z(o[1753]) );
  AND U27491 ( .A(p_input[1753]), .B(p_input[11753]), .Z(n18328) );
  AND U27492 ( .A(p_input[31753]), .B(p_input[21753]), .Z(n18327) );
  AND U27493 ( .A(n18329), .B(n18330), .Z(o[1752]) );
  AND U27494 ( .A(p_input[1752]), .B(p_input[11752]), .Z(n18330) );
  AND U27495 ( .A(p_input[31752]), .B(p_input[21752]), .Z(n18329) );
  AND U27496 ( .A(n18331), .B(n18332), .Z(o[1751]) );
  AND U27497 ( .A(p_input[1751]), .B(p_input[11751]), .Z(n18332) );
  AND U27498 ( .A(p_input[31751]), .B(p_input[21751]), .Z(n18331) );
  AND U27499 ( .A(n18333), .B(n18334), .Z(o[1750]) );
  AND U27500 ( .A(p_input[1750]), .B(p_input[11750]), .Z(n18334) );
  AND U27501 ( .A(p_input[31750]), .B(p_input[21750]), .Z(n18333) );
  AND U27502 ( .A(n18335), .B(n18336), .Z(o[174]) );
  AND U27503 ( .A(p_input[174]), .B(p_input[10174]), .Z(n18336) );
  AND U27504 ( .A(p_input[30174]), .B(p_input[20174]), .Z(n18335) );
  AND U27505 ( .A(n18337), .B(n18338), .Z(o[1749]) );
  AND U27506 ( .A(p_input[1749]), .B(p_input[11749]), .Z(n18338) );
  AND U27507 ( .A(p_input[31749]), .B(p_input[21749]), .Z(n18337) );
  AND U27508 ( .A(n18339), .B(n18340), .Z(o[1748]) );
  AND U27509 ( .A(p_input[1748]), .B(p_input[11748]), .Z(n18340) );
  AND U27510 ( .A(p_input[31748]), .B(p_input[21748]), .Z(n18339) );
  AND U27511 ( .A(n18341), .B(n18342), .Z(o[1747]) );
  AND U27512 ( .A(p_input[1747]), .B(p_input[11747]), .Z(n18342) );
  AND U27513 ( .A(p_input[31747]), .B(p_input[21747]), .Z(n18341) );
  AND U27514 ( .A(n18343), .B(n18344), .Z(o[1746]) );
  AND U27515 ( .A(p_input[1746]), .B(p_input[11746]), .Z(n18344) );
  AND U27516 ( .A(p_input[31746]), .B(p_input[21746]), .Z(n18343) );
  AND U27517 ( .A(n18345), .B(n18346), .Z(o[1745]) );
  AND U27518 ( .A(p_input[1745]), .B(p_input[11745]), .Z(n18346) );
  AND U27519 ( .A(p_input[31745]), .B(p_input[21745]), .Z(n18345) );
  AND U27520 ( .A(n18347), .B(n18348), .Z(o[1744]) );
  AND U27521 ( .A(p_input[1744]), .B(p_input[11744]), .Z(n18348) );
  AND U27522 ( .A(p_input[31744]), .B(p_input[21744]), .Z(n18347) );
  AND U27523 ( .A(n18349), .B(n18350), .Z(o[1743]) );
  AND U27524 ( .A(p_input[1743]), .B(p_input[11743]), .Z(n18350) );
  AND U27525 ( .A(p_input[31743]), .B(p_input[21743]), .Z(n18349) );
  AND U27526 ( .A(n18351), .B(n18352), .Z(o[1742]) );
  AND U27527 ( .A(p_input[1742]), .B(p_input[11742]), .Z(n18352) );
  AND U27528 ( .A(p_input[31742]), .B(p_input[21742]), .Z(n18351) );
  AND U27529 ( .A(n18353), .B(n18354), .Z(o[1741]) );
  AND U27530 ( .A(p_input[1741]), .B(p_input[11741]), .Z(n18354) );
  AND U27531 ( .A(p_input[31741]), .B(p_input[21741]), .Z(n18353) );
  AND U27532 ( .A(n18355), .B(n18356), .Z(o[1740]) );
  AND U27533 ( .A(p_input[1740]), .B(p_input[11740]), .Z(n18356) );
  AND U27534 ( .A(p_input[31740]), .B(p_input[21740]), .Z(n18355) );
  AND U27535 ( .A(n18357), .B(n18358), .Z(o[173]) );
  AND U27536 ( .A(p_input[173]), .B(p_input[10173]), .Z(n18358) );
  AND U27537 ( .A(p_input[30173]), .B(p_input[20173]), .Z(n18357) );
  AND U27538 ( .A(n18359), .B(n18360), .Z(o[1739]) );
  AND U27539 ( .A(p_input[1739]), .B(p_input[11739]), .Z(n18360) );
  AND U27540 ( .A(p_input[31739]), .B(p_input[21739]), .Z(n18359) );
  AND U27541 ( .A(n18361), .B(n18362), .Z(o[1738]) );
  AND U27542 ( .A(p_input[1738]), .B(p_input[11738]), .Z(n18362) );
  AND U27543 ( .A(p_input[31738]), .B(p_input[21738]), .Z(n18361) );
  AND U27544 ( .A(n18363), .B(n18364), .Z(o[1737]) );
  AND U27545 ( .A(p_input[1737]), .B(p_input[11737]), .Z(n18364) );
  AND U27546 ( .A(p_input[31737]), .B(p_input[21737]), .Z(n18363) );
  AND U27547 ( .A(n18365), .B(n18366), .Z(o[1736]) );
  AND U27548 ( .A(p_input[1736]), .B(p_input[11736]), .Z(n18366) );
  AND U27549 ( .A(p_input[31736]), .B(p_input[21736]), .Z(n18365) );
  AND U27550 ( .A(n18367), .B(n18368), .Z(o[1735]) );
  AND U27551 ( .A(p_input[1735]), .B(p_input[11735]), .Z(n18368) );
  AND U27552 ( .A(p_input[31735]), .B(p_input[21735]), .Z(n18367) );
  AND U27553 ( .A(n18369), .B(n18370), .Z(o[1734]) );
  AND U27554 ( .A(p_input[1734]), .B(p_input[11734]), .Z(n18370) );
  AND U27555 ( .A(p_input[31734]), .B(p_input[21734]), .Z(n18369) );
  AND U27556 ( .A(n18371), .B(n18372), .Z(o[1733]) );
  AND U27557 ( .A(p_input[1733]), .B(p_input[11733]), .Z(n18372) );
  AND U27558 ( .A(p_input[31733]), .B(p_input[21733]), .Z(n18371) );
  AND U27559 ( .A(n18373), .B(n18374), .Z(o[1732]) );
  AND U27560 ( .A(p_input[1732]), .B(p_input[11732]), .Z(n18374) );
  AND U27561 ( .A(p_input[31732]), .B(p_input[21732]), .Z(n18373) );
  AND U27562 ( .A(n18375), .B(n18376), .Z(o[1731]) );
  AND U27563 ( .A(p_input[1731]), .B(p_input[11731]), .Z(n18376) );
  AND U27564 ( .A(p_input[31731]), .B(p_input[21731]), .Z(n18375) );
  AND U27565 ( .A(n18377), .B(n18378), .Z(o[1730]) );
  AND U27566 ( .A(p_input[1730]), .B(p_input[11730]), .Z(n18378) );
  AND U27567 ( .A(p_input[31730]), .B(p_input[21730]), .Z(n18377) );
  AND U27568 ( .A(n18379), .B(n18380), .Z(o[172]) );
  AND U27569 ( .A(p_input[172]), .B(p_input[10172]), .Z(n18380) );
  AND U27570 ( .A(p_input[30172]), .B(p_input[20172]), .Z(n18379) );
  AND U27571 ( .A(n18381), .B(n18382), .Z(o[1729]) );
  AND U27572 ( .A(p_input[1729]), .B(p_input[11729]), .Z(n18382) );
  AND U27573 ( .A(p_input[31729]), .B(p_input[21729]), .Z(n18381) );
  AND U27574 ( .A(n18383), .B(n18384), .Z(o[1728]) );
  AND U27575 ( .A(p_input[1728]), .B(p_input[11728]), .Z(n18384) );
  AND U27576 ( .A(p_input[31728]), .B(p_input[21728]), .Z(n18383) );
  AND U27577 ( .A(n18385), .B(n18386), .Z(o[1727]) );
  AND U27578 ( .A(p_input[1727]), .B(p_input[11727]), .Z(n18386) );
  AND U27579 ( .A(p_input[31727]), .B(p_input[21727]), .Z(n18385) );
  AND U27580 ( .A(n18387), .B(n18388), .Z(o[1726]) );
  AND U27581 ( .A(p_input[1726]), .B(p_input[11726]), .Z(n18388) );
  AND U27582 ( .A(p_input[31726]), .B(p_input[21726]), .Z(n18387) );
  AND U27583 ( .A(n18389), .B(n18390), .Z(o[1725]) );
  AND U27584 ( .A(p_input[1725]), .B(p_input[11725]), .Z(n18390) );
  AND U27585 ( .A(p_input[31725]), .B(p_input[21725]), .Z(n18389) );
  AND U27586 ( .A(n18391), .B(n18392), .Z(o[1724]) );
  AND U27587 ( .A(p_input[1724]), .B(p_input[11724]), .Z(n18392) );
  AND U27588 ( .A(p_input[31724]), .B(p_input[21724]), .Z(n18391) );
  AND U27589 ( .A(n18393), .B(n18394), .Z(o[1723]) );
  AND U27590 ( .A(p_input[1723]), .B(p_input[11723]), .Z(n18394) );
  AND U27591 ( .A(p_input[31723]), .B(p_input[21723]), .Z(n18393) );
  AND U27592 ( .A(n18395), .B(n18396), .Z(o[1722]) );
  AND U27593 ( .A(p_input[1722]), .B(p_input[11722]), .Z(n18396) );
  AND U27594 ( .A(p_input[31722]), .B(p_input[21722]), .Z(n18395) );
  AND U27595 ( .A(n18397), .B(n18398), .Z(o[1721]) );
  AND U27596 ( .A(p_input[1721]), .B(p_input[11721]), .Z(n18398) );
  AND U27597 ( .A(p_input[31721]), .B(p_input[21721]), .Z(n18397) );
  AND U27598 ( .A(n18399), .B(n18400), .Z(o[1720]) );
  AND U27599 ( .A(p_input[1720]), .B(p_input[11720]), .Z(n18400) );
  AND U27600 ( .A(p_input[31720]), .B(p_input[21720]), .Z(n18399) );
  AND U27601 ( .A(n18401), .B(n18402), .Z(o[171]) );
  AND U27602 ( .A(p_input[171]), .B(p_input[10171]), .Z(n18402) );
  AND U27603 ( .A(p_input[30171]), .B(p_input[20171]), .Z(n18401) );
  AND U27604 ( .A(n18403), .B(n18404), .Z(o[1719]) );
  AND U27605 ( .A(p_input[1719]), .B(p_input[11719]), .Z(n18404) );
  AND U27606 ( .A(p_input[31719]), .B(p_input[21719]), .Z(n18403) );
  AND U27607 ( .A(n18405), .B(n18406), .Z(o[1718]) );
  AND U27608 ( .A(p_input[1718]), .B(p_input[11718]), .Z(n18406) );
  AND U27609 ( .A(p_input[31718]), .B(p_input[21718]), .Z(n18405) );
  AND U27610 ( .A(n18407), .B(n18408), .Z(o[1717]) );
  AND U27611 ( .A(p_input[1717]), .B(p_input[11717]), .Z(n18408) );
  AND U27612 ( .A(p_input[31717]), .B(p_input[21717]), .Z(n18407) );
  AND U27613 ( .A(n18409), .B(n18410), .Z(o[1716]) );
  AND U27614 ( .A(p_input[1716]), .B(p_input[11716]), .Z(n18410) );
  AND U27615 ( .A(p_input[31716]), .B(p_input[21716]), .Z(n18409) );
  AND U27616 ( .A(n18411), .B(n18412), .Z(o[1715]) );
  AND U27617 ( .A(p_input[1715]), .B(p_input[11715]), .Z(n18412) );
  AND U27618 ( .A(p_input[31715]), .B(p_input[21715]), .Z(n18411) );
  AND U27619 ( .A(n18413), .B(n18414), .Z(o[1714]) );
  AND U27620 ( .A(p_input[1714]), .B(p_input[11714]), .Z(n18414) );
  AND U27621 ( .A(p_input[31714]), .B(p_input[21714]), .Z(n18413) );
  AND U27622 ( .A(n18415), .B(n18416), .Z(o[1713]) );
  AND U27623 ( .A(p_input[1713]), .B(p_input[11713]), .Z(n18416) );
  AND U27624 ( .A(p_input[31713]), .B(p_input[21713]), .Z(n18415) );
  AND U27625 ( .A(n18417), .B(n18418), .Z(o[1712]) );
  AND U27626 ( .A(p_input[1712]), .B(p_input[11712]), .Z(n18418) );
  AND U27627 ( .A(p_input[31712]), .B(p_input[21712]), .Z(n18417) );
  AND U27628 ( .A(n18419), .B(n18420), .Z(o[1711]) );
  AND U27629 ( .A(p_input[1711]), .B(p_input[11711]), .Z(n18420) );
  AND U27630 ( .A(p_input[31711]), .B(p_input[21711]), .Z(n18419) );
  AND U27631 ( .A(n18421), .B(n18422), .Z(o[1710]) );
  AND U27632 ( .A(p_input[1710]), .B(p_input[11710]), .Z(n18422) );
  AND U27633 ( .A(p_input[31710]), .B(p_input[21710]), .Z(n18421) );
  AND U27634 ( .A(n18423), .B(n18424), .Z(o[170]) );
  AND U27635 ( .A(p_input[170]), .B(p_input[10170]), .Z(n18424) );
  AND U27636 ( .A(p_input[30170]), .B(p_input[20170]), .Z(n18423) );
  AND U27637 ( .A(n18425), .B(n18426), .Z(o[1709]) );
  AND U27638 ( .A(p_input[1709]), .B(p_input[11709]), .Z(n18426) );
  AND U27639 ( .A(p_input[31709]), .B(p_input[21709]), .Z(n18425) );
  AND U27640 ( .A(n18427), .B(n18428), .Z(o[1708]) );
  AND U27641 ( .A(p_input[1708]), .B(p_input[11708]), .Z(n18428) );
  AND U27642 ( .A(p_input[31708]), .B(p_input[21708]), .Z(n18427) );
  AND U27643 ( .A(n18429), .B(n18430), .Z(o[1707]) );
  AND U27644 ( .A(p_input[1707]), .B(p_input[11707]), .Z(n18430) );
  AND U27645 ( .A(p_input[31707]), .B(p_input[21707]), .Z(n18429) );
  AND U27646 ( .A(n18431), .B(n18432), .Z(o[1706]) );
  AND U27647 ( .A(p_input[1706]), .B(p_input[11706]), .Z(n18432) );
  AND U27648 ( .A(p_input[31706]), .B(p_input[21706]), .Z(n18431) );
  AND U27649 ( .A(n18433), .B(n18434), .Z(o[1705]) );
  AND U27650 ( .A(p_input[1705]), .B(p_input[11705]), .Z(n18434) );
  AND U27651 ( .A(p_input[31705]), .B(p_input[21705]), .Z(n18433) );
  AND U27652 ( .A(n18435), .B(n18436), .Z(o[1704]) );
  AND U27653 ( .A(p_input[1704]), .B(p_input[11704]), .Z(n18436) );
  AND U27654 ( .A(p_input[31704]), .B(p_input[21704]), .Z(n18435) );
  AND U27655 ( .A(n18437), .B(n18438), .Z(o[1703]) );
  AND U27656 ( .A(p_input[1703]), .B(p_input[11703]), .Z(n18438) );
  AND U27657 ( .A(p_input[31703]), .B(p_input[21703]), .Z(n18437) );
  AND U27658 ( .A(n18439), .B(n18440), .Z(o[1702]) );
  AND U27659 ( .A(p_input[1702]), .B(p_input[11702]), .Z(n18440) );
  AND U27660 ( .A(p_input[31702]), .B(p_input[21702]), .Z(n18439) );
  AND U27661 ( .A(n18441), .B(n18442), .Z(o[1701]) );
  AND U27662 ( .A(p_input[1701]), .B(p_input[11701]), .Z(n18442) );
  AND U27663 ( .A(p_input[31701]), .B(p_input[21701]), .Z(n18441) );
  AND U27664 ( .A(n18443), .B(n18444), .Z(o[1700]) );
  AND U27665 ( .A(p_input[1700]), .B(p_input[11700]), .Z(n18444) );
  AND U27666 ( .A(p_input[31700]), .B(p_input[21700]), .Z(n18443) );
  AND U27667 ( .A(n18445), .B(n18446), .Z(o[16]) );
  AND U27668 ( .A(p_input[16]), .B(p_input[10016]), .Z(n18446) );
  AND U27669 ( .A(p_input[30016]), .B(p_input[20016]), .Z(n18445) );
  AND U27670 ( .A(n18447), .B(n18448), .Z(o[169]) );
  AND U27671 ( .A(p_input[169]), .B(p_input[10169]), .Z(n18448) );
  AND U27672 ( .A(p_input[30169]), .B(p_input[20169]), .Z(n18447) );
  AND U27673 ( .A(n18449), .B(n18450), .Z(o[1699]) );
  AND U27674 ( .A(p_input[1699]), .B(p_input[11699]), .Z(n18450) );
  AND U27675 ( .A(p_input[31699]), .B(p_input[21699]), .Z(n18449) );
  AND U27676 ( .A(n18451), .B(n18452), .Z(o[1698]) );
  AND U27677 ( .A(p_input[1698]), .B(p_input[11698]), .Z(n18452) );
  AND U27678 ( .A(p_input[31698]), .B(p_input[21698]), .Z(n18451) );
  AND U27679 ( .A(n18453), .B(n18454), .Z(o[1697]) );
  AND U27680 ( .A(p_input[1697]), .B(p_input[11697]), .Z(n18454) );
  AND U27681 ( .A(p_input[31697]), .B(p_input[21697]), .Z(n18453) );
  AND U27682 ( .A(n18455), .B(n18456), .Z(o[1696]) );
  AND U27683 ( .A(p_input[1696]), .B(p_input[11696]), .Z(n18456) );
  AND U27684 ( .A(p_input[31696]), .B(p_input[21696]), .Z(n18455) );
  AND U27685 ( .A(n18457), .B(n18458), .Z(o[1695]) );
  AND U27686 ( .A(p_input[1695]), .B(p_input[11695]), .Z(n18458) );
  AND U27687 ( .A(p_input[31695]), .B(p_input[21695]), .Z(n18457) );
  AND U27688 ( .A(n18459), .B(n18460), .Z(o[1694]) );
  AND U27689 ( .A(p_input[1694]), .B(p_input[11694]), .Z(n18460) );
  AND U27690 ( .A(p_input[31694]), .B(p_input[21694]), .Z(n18459) );
  AND U27691 ( .A(n18461), .B(n18462), .Z(o[1693]) );
  AND U27692 ( .A(p_input[1693]), .B(p_input[11693]), .Z(n18462) );
  AND U27693 ( .A(p_input[31693]), .B(p_input[21693]), .Z(n18461) );
  AND U27694 ( .A(n18463), .B(n18464), .Z(o[1692]) );
  AND U27695 ( .A(p_input[1692]), .B(p_input[11692]), .Z(n18464) );
  AND U27696 ( .A(p_input[31692]), .B(p_input[21692]), .Z(n18463) );
  AND U27697 ( .A(n18465), .B(n18466), .Z(o[1691]) );
  AND U27698 ( .A(p_input[1691]), .B(p_input[11691]), .Z(n18466) );
  AND U27699 ( .A(p_input[31691]), .B(p_input[21691]), .Z(n18465) );
  AND U27700 ( .A(n18467), .B(n18468), .Z(o[1690]) );
  AND U27701 ( .A(p_input[1690]), .B(p_input[11690]), .Z(n18468) );
  AND U27702 ( .A(p_input[31690]), .B(p_input[21690]), .Z(n18467) );
  AND U27703 ( .A(n18469), .B(n18470), .Z(o[168]) );
  AND U27704 ( .A(p_input[168]), .B(p_input[10168]), .Z(n18470) );
  AND U27705 ( .A(p_input[30168]), .B(p_input[20168]), .Z(n18469) );
  AND U27706 ( .A(n18471), .B(n18472), .Z(o[1689]) );
  AND U27707 ( .A(p_input[1689]), .B(p_input[11689]), .Z(n18472) );
  AND U27708 ( .A(p_input[31689]), .B(p_input[21689]), .Z(n18471) );
  AND U27709 ( .A(n18473), .B(n18474), .Z(o[1688]) );
  AND U27710 ( .A(p_input[1688]), .B(p_input[11688]), .Z(n18474) );
  AND U27711 ( .A(p_input[31688]), .B(p_input[21688]), .Z(n18473) );
  AND U27712 ( .A(n18475), .B(n18476), .Z(o[1687]) );
  AND U27713 ( .A(p_input[1687]), .B(p_input[11687]), .Z(n18476) );
  AND U27714 ( .A(p_input[31687]), .B(p_input[21687]), .Z(n18475) );
  AND U27715 ( .A(n18477), .B(n18478), .Z(o[1686]) );
  AND U27716 ( .A(p_input[1686]), .B(p_input[11686]), .Z(n18478) );
  AND U27717 ( .A(p_input[31686]), .B(p_input[21686]), .Z(n18477) );
  AND U27718 ( .A(n18479), .B(n18480), .Z(o[1685]) );
  AND U27719 ( .A(p_input[1685]), .B(p_input[11685]), .Z(n18480) );
  AND U27720 ( .A(p_input[31685]), .B(p_input[21685]), .Z(n18479) );
  AND U27721 ( .A(n18481), .B(n18482), .Z(o[1684]) );
  AND U27722 ( .A(p_input[1684]), .B(p_input[11684]), .Z(n18482) );
  AND U27723 ( .A(p_input[31684]), .B(p_input[21684]), .Z(n18481) );
  AND U27724 ( .A(n18483), .B(n18484), .Z(o[1683]) );
  AND U27725 ( .A(p_input[1683]), .B(p_input[11683]), .Z(n18484) );
  AND U27726 ( .A(p_input[31683]), .B(p_input[21683]), .Z(n18483) );
  AND U27727 ( .A(n18485), .B(n18486), .Z(o[1682]) );
  AND U27728 ( .A(p_input[1682]), .B(p_input[11682]), .Z(n18486) );
  AND U27729 ( .A(p_input[31682]), .B(p_input[21682]), .Z(n18485) );
  AND U27730 ( .A(n18487), .B(n18488), .Z(o[1681]) );
  AND U27731 ( .A(p_input[1681]), .B(p_input[11681]), .Z(n18488) );
  AND U27732 ( .A(p_input[31681]), .B(p_input[21681]), .Z(n18487) );
  AND U27733 ( .A(n18489), .B(n18490), .Z(o[1680]) );
  AND U27734 ( .A(p_input[1680]), .B(p_input[11680]), .Z(n18490) );
  AND U27735 ( .A(p_input[31680]), .B(p_input[21680]), .Z(n18489) );
  AND U27736 ( .A(n18491), .B(n18492), .Z(o[167]) );
  AND U27737 ( .A(p_input[167]), .B(p_input[10167]), .Z(n18492) );
  AND U27738 ( .A(p_input[30167]), .B(p_input[20167]), .Z(n18491) );
  AND U27739 ( .A(n18493), .B(n18494), .Z(o[1679]) );
  AND U27740 ( .A(p_input[1679]), .B(p_input[11679]), .Z(n18494) );
  AND U27741 ( .A(p_input[31679]), .B(p_input[21679]), .Z(n18493) );
  AND U27742 ( .A(n18495), .B(n18496), .Z(o[1678]) );
  AND U27743 ( .A(p_input[1678]), .B(p_input[11678]), .Z(n18496) );
  AND U27744 ( .A(p_input[31678]), .B(p_input[21678]), .Z(n18495) );
  AND U27745 ( .A(n18497), .B(n18498), .Z(o[1677]) );
  AND U27746 ( .A(p_input[1677]), .B(p_input[11677]), .Z(n18498) );
  AND U27747 ( .A(p_input[31677]), .B(p_input[21677]), .Z(n18497) );
  AND U27748 ( .A(n18499), .B(n18500), .Z(o[1676]) );
  AND U27749 ( .A(p_input[1676]), .B(p_input[11676]), .Z(n18500) );
  AND U27750 ( .A(p_input[31676]), .B(p_input[21676]), .Z(n18499) );
  AND U27751 ( .A(n18501), .B(n18502), .Z(o[1675]) );
  AND U27752 ( .A(p_input[1675]), .B(p_input[11675]), .Z(n18502) );
  AND U27753 ( .A(p_input[31675]), .B(p_input[21675]), .Z(n18501) );
  AND U27754 ( .A(n18503), .B(n18504), .Z(o[1674]) );
  AND U27755 ( .A(p_input[1674]), .B(p_input[11674]), .Z(n18504) );
  AND U27756 ( .A(p_input[31674]), .B(p_input[21674]), .Z(n18503) );
  AND U27757 ( .A(n18505), .B(n18506), .Z(o[1673]) );
  AND U27758 ( .A(p_input[1673]), .B(p_input[11673]), .Z(n18506) );
  AND U27759 ( .A(p_input[31673]), .B(p_input[21673]), .Z(n18505) );
  AND U27760 ( .A(n18507), .B(n18508), .Z(o[1672]) );
  AND U27761 ( .A(p_input[1672]), .B(p_input[11672]), .Z(n18508) );
  AND U27762 ( .A(p_input[31672]), .B(p_input[21672]), .Z(n18507) );
  AND U27763 ( .A(n18509), .B(n18510), .Z(o[1671]) );
  AND U27764 ( .A(p_input[1671]), .B(p_input[11671]), .Z(n18510) );
  AND U27765 ( .A(p_input[31671]), .B(p_input[21671]), .Z(n18509) );
  AND U27766 ( .A(n18511), .B(n18512), .Z(o[1670]) );
  AND U27767 ( .A(p_input[1670]), .B(p_input[11670]), .Z(n18512) );
  AND U27768 ( .A(p_input[31670]), .B(p_input[21670]), .Z(n18511) );
  AND U27769 ( .A(n18513), .B(n18514), .Z(o[166]) );
  AND U27770 ( .A(p_input[166]), .B(p_input[10166]), .Z(n18514) );
  AND U27771 ( .A(p_input[30166]), .B(p_input[20166]), .Z(n18513) );
  AND U27772 ( .A(n18515), .B(n18516), .Z(o[1669]) );
  AND U27773 ( .A(p_input[1669]), .B(p_input[11669]), .Z(n18516) );
  AND U27774 ( .A(p_input[31669]), .B(p_input[21669]), .Z(n18515) );
  AND U27775 ( .A(n18517), .B(n18518), .Z(o[1668]) );
  AND U27776 ( .A(p_input[1668]), .B(p_input[11668]), .Z(n18518) );
  AND U27777 ( .A(p_input[31668]), .B(p_input[21668]), .Z(n18517) );
  AND U27778 ( .A(n18519), .B(n18520), .Z(o[1667]) );
  AND U27779 ( .A(p_input[1667]), .B(p_input[11667]), .Z(n18520) );
  AND U27780 ( .A(p_input[31667]), .B(p_input[21667]), .Z(n18519) );
  AND U27781 ( .A(n18521), .B(n18522), .Z(o[1666]) );
  AND U27782 ( .A(p_input[1666]), .B(p_input[11666]), .Z(n18522) );
  AND U27783 ( .A(p_input[31666]), .B(p_input[21666]), .Z(n18521) );
  AND U27784 ( .A(n18523), .B(n18524), .Z(o[1665]) );
  AND U27785 ( .A(p_input[1665]), .B(p_input[11665]), .Z(n18524) );
  AND U27786 ( .A(p_input[31665]), .B(p_input[21665]), .Z(n18523) );
  AND U27787 ( .A(n18525), .B(n18526), .Z(o[1664]) );
  AND U27788 ( .A(p_input[1664]), .B(p_input[11664]), .Z(n18526) );
  AND U27789 ( .A(p_input[31664]), .B(p_input[21664]), .Z(n18525) );
  AND U27790 ( .A(n18527), .B(n18528), .Z(o[1663]) );
  AND U27791 ( .A(p_input[1663]), .B(p_input[11663]), .Z(n18528) );
  AND U27792 ( .A(p_input[31663]), .B(p_input[21663]), .Z(n18527) );
  AND U27793 ( .A(n18529), .B(n18530), .Z(o[1662]) );
  AND U27794 ( .A(p_input[1662]), .B(p_input[11662]), .Z(n18530) );
  AND U27795 ( .A(p_input[31662]), .B(p_input[21662]), .Z(n18529) );
  AND U27796 ( .A(n18531), .B(n18532), .Z(o[1661]) );
  AND U27797 ( .A(p_input[1661]), .B(p_input[11661]), .Z(n18532) );
  AND U27798 ( .A(p_input[31661]), .B(p_input[21661]), .Z(n18531) );
  AND U27799 ( .A(n18533), .B(n18534), .Z(o[1660]) );
  AND U27800 ( .A(p_input[1660]), .B(p_input[11660]), .Z(n18534) );
  AND U27801 ( .A(p_input[31660]), .B(p_input[21660]), .Z(n18533) );
  AND U27802 ( .A(n18535), .B(n18536), .Z(o[165]) );
  AND U27803 ( .A(p_input[165]), .B(p_input[10165]), .Z(n18536) );
  AND U27804 ( .A(p_input[30165]), .B(p_input[20165]), .Z(n18535) );
  AND U27805 ( .A(n18537), .B(n18538), .Z(o[1659]) );
  AND U27806 ( .A(p_input[1659]), .B(p_input[11659]), .Z(n18538) );
  AND U27807 ( .A(p_input[31659]), .B(p_input[21659]), .Z(n18537) );
  AND U27808 ( .A(n18539), .B(n18540), .Z(o[1658]) );
  AND U27809 ( .A(p_input[1658]), .B(p_input[11658]), .Z(n18540) );
  AND U27810 ( .A(p_input[31658]), .B(p_input[21658]), .Z(n18539) );
  AND U27811 ( .A(n18541), .B(n18542), .Z(o[1657]) );
  AND U27812 ( .A(p_input[1657]), .B(p_input[11657]), .Z(n18542) );
  AND U27813 ( .A(p_input[31657]), .B(p_input[21657]), .Z(n18541) );
  AND U27814 ( .A(n18543), .B(n18544), .Z(o[1656]) );
  AND U27815 ( .A(p_input[1656]), .B(p_input[11656]), .Z(n18544) );
  AND U27816 ( .A(p_input[31656]), .B(p_input[21656]), .Z(n18543) );
  AND U27817 ( .A(n18545), .B(n18546), .Z(o[1655]) );
  AND U27818 ( .A(p_input[1655]), .B(p_input[11655]), .Z(n18546) );
  AND U27819 ( .A(p_input[31655]), .B(p_input[21655]), .Z(n18545) );
  AND U27820 ( .A(n18547), .B(n18548), .Z(o[1654]) );
  AND U27821 ( .A(p_input[1654]), .B(p_input[11654]), .Z(n18548) );
  AND U27822 ( .A(p_input[31654]), .B(p_input[21654]), .Z(n18547) );
  AND U27823 ( .A(n18549), .B(n18550), .Z(o[1653]) );
  AND U27824 ( .A(p_input[1653]), .B(p_input[11653]), .Z(n18550) );
  AND U27825 ( .A(p_input[31653]), .B(p_input[21653]), .Z(n18549) );
  AND U27826 ( .A(n18551), .B(n18552), .Z(o[1652]) );
  AND U27827 ( .A(p_input[1652]), .B(p_input[11652]), .Z(n18552) );
  AND U27828 ( .A(p_input[31652]), .B(p_input[21652]), .Z(n18551) );
  AND U27829 ( .A(n18553), .B(n18554), .Z(o[1651]) );
  AND U27830 ( .A(p_input[1651]), .B(p_input[11651]), .Z(n18554) );
  AND U27831 ( .A(p_input[31651]), .B(p_input[21651]), .Z(n18553) );
  AND U27832 ( .A(n18555), .B(n18556), .Z(o[1650]) );
  AND U27833 ( .A(p_input[1650]), .B(p_input[11650]), .Z(n18556) );
  AND U27834 ( .A(p_input[31650]), .B(p_input[21650]), .Z(n18555) );
  AND U27835 ( .A(n18557), .B(n18558), .Z(o[164]) );
  AND U27836 ( .A(p_input[164]), .B(p_input[10164]), .Z(n18558) );
  AND U27837 ( .A(p_input[30164]), .B(p_input[20164]), .Z(n18557) );
  AND U27838 ( .A(n18559), .B(n18560), .Z(o[1649]) );
  AND U27839 ( .A(p_input[1649]), .B(p_input[11649]), .Z(n18560) );
  AND U27840 ( .A(p_input[31649]), .B(p_input[21649]), .Z(n18559) );
  AND U27841 ( .A(n18561), .B(n18562), .Z(o[1648]) );
  AND U27842 ( .A(p_input[1648]), .B(p_input[11648]), .Z(n18562) );
  AND U27843 ( .A(p_input[31648]), .B(p_input[21648]), .Z(n18561) );
  AND U27844 ( .A(n18563), .B(n18564), .Z(o[1647]) );
  AND U27845 ( .A(p_input[1647]), .B(p_input[11647]), .Z(n18564) );
  AND U27846 ( .A(p_input[31647]), .B(p_input[21647]), .Z(n18563) );
  AND U27847 ( .A(n18565), .B(n18566), .Z(o[1646]) );
  AND U27848 ( .A(p_input[1646]), .B(p_input[11646]), .Z(n18566) );
  AND U27849 ( .A(p_input[31646]), .B(p_input[21646]), .Z(n18565) );
  AND U27850 ( .A(n18567), .B(n18568), .Z(o[1645]) );
  AND U27851 ( .A(p_input[1645]), .B(p_input[11645]), .Z(n18568) );
  AND U27852 ( .A(p_input[31645]), .B(p_input[21645]), .Z(n18567) );
  AND U27853 ( .A(n18569), .B(n18570), .Z(o[1644]) );
  AND U27854 ( .A(p_input[1644]), .B(p_input[11644]), .Z(n18570) );
  AND U27855 ( .A(p_input[31644]), .B(p_input[21644]), .Z(n18569) );
  AND U27856 ( .A(n18571), .B(n18572), .Z(o[1643]) );
  AND U27857 ( .A(p_input[1643]), .B(p_input[11643]), .Z(n18572) );
  AND U27858 ( .A(p_input[31643]), .B(p_input[21643]), .Z(n18571) );
  AND U27859 ( .A(n18573), .B(n18574), .Z(o[1642]) );
  AND U27860 ( .A(p_input[1642]), .B(p_input[11642]), .Z(n18574) );
  AND U27861 ( .A(p_input[31642]), .B(p_input[21642]), .Z(n18573) );
  AND U27862 ( .A(n18575), .B(n18576), .Z(o[1641]) );
  AND U27863 ( .A(p_input[1641]), .B(p_input[11641]), .Z(n18576) );
  AND U27864 ( .A(p_input[31641]), .B(p_input[21641]), .Z(n18575) );
  AND U27865 ( .A(n18577), .B(n18578), .Z(o[1640]) );
  AND U27866 ( .A(p_input[1640]), .B(p_input[11640]), .Z(n18578) );
  AND U27867 ( .A(p_input[31640]), .B(p_input[21640]), .Z(n18577) );
  AND U27868 ( .A(n18579), .B(n18580), .Z(o[163]) );
  AND U27869 ( .A(p_input[163]), .B(p_input[10163]), .Z(n18580) );
  AND U27870 ( .A(p_input[30163]), .B(p_input[20163]), .Z(n18579) );
  AND U27871 ( .A(n18581), .B(n18582), .Z(o[1639]) );
  AND U27872 ( .A(p_input[1639]), .B(p_input[11639]), .Z(n18582) );
  AND U27873 ( .A(p_input[31639]), .B(p_input[21639]), .Z(n18581) );
  AND U27874 ( .A(n18583), .B(n18584), .Z(o[1638]) );
  AND U27875 ( .A(p_input[1638]), .B(p_input[11638]), .Z(n18584) );
  AND U27876 ( .A(p_input[31638]), .B(p_input[21638]), .Z(n18583) );
  AND U27877 ( .A(n18585), .B(n18586), .Z(o[1637]) );
  AND U27878 ( .A(p_input[1637]), .B(p_input[11637]), .Z(n18586) );
  AND U27879 ( .A(p_input[31637]), .B(p_input[21637]), .Z(n18585) );
  AND U27880 ( .A(n18587), .B(n18588), .Z(o[1636]) );
  AND U27881 ( .A(p_input[1636]), .B(p_input[11636]), .Z(n18588) );
  AND U27882 ( .A(p_input[31636]), .B(p_input[21636]), .Z(n18587) );
  AND U27883 ( .A(n18589), .B(n18590), .Z(o[1635]) );
  AND U27884 ( .A(p_input[1635]), .B(p_input[11635]), .Z(n18590) );
  AND U27885 ( .A(p_input[31635]), .B(p_input[21635]), .Z(n18589) );
  AND U27886 ( .A(n18591), .B(n18592), .Z(o[1634]) );
  AND U27887 ( .A(p_input[1634]), .B(p_input[11634]), .Z(n18592) );
  AND U27888 ( .A(p_input[31634]), .B(p_input[21634]), .Z(n18591) );
  AND U27889 ( .A(n18593), .B(n18594), .Z(o[1633]) );
  AND U27890 ( .A(p_input[1633]), .B(p_input[11633]), .Z(n18594) );
  AND U27891 ( .A(p_input[31633]), .B(p_input[21633]), .Z(n18593) );
  AND U27892 ( .A(n18595), .B(n18596), .Z(o[1632]) );
  AND U27893 ( .A(p_input[1632]), .B(p_input[11632]), .Z(n18596) );
  AND U27894 ( .A(p_input[31632]), .B(p_input[21632]), .Z(n18595) );
  AND U27895 ( .A(n18597), .B(n18598), .Z(o[1631]) );
  AND U27896 ( .A(p_input[1631]), .B(p_input[11631]), .Z(n18598) );
  AND U27897 ( .A(p_input[31631]), .B(p_input[21631]), .Z(n18597) );
  AND U27898 ( .A(n18599), .B(n18600), .Z(o[1630]) );
  AND U27899 ( .A(p_input[1630]), .B(p_input[11630]), .Z(n18600) );
  AND U27900 ( .A(p_input[31630]), .B(p_input[21630]), .Z(n18599) );
  AND U27901 ( .A(n18601), .B(n18602), .Z(o[162]) );
  AND U27902 ( .A(p_input[162]), .B(p_input[10162]), .Z(n18602) );
  AND U27903 ( .A(p_input[30162]), .B(p_input[20162]), .Z(n18601) );
  AND U27904 ( .A(n18603), .B(n18604), .Z(o[1629]) );
  AND U27905 ( .A(p_input[1629]), .B(p_input[11629]), .Z(n18604) );
  AND U27906 ( .A(p_input[31629]), .B(p_input[21629]), .Z(n18603) );
  AND U27907 ( .A(n18605), .B(n18606), .Z(o[1628]) );
  AND U27908 ( .A(p_input[1628]), .B(p_input[11628]), .Z(n18606) );
  AND U27909 ( .A(p_input[31628]), .B(p_input[21628]), .Z(n18605) );
  AND U27910 ( .A(n18607), .B(n18608), .Z(o[1627]) );
  AND U27911 ( .A(p_input[1627]), .B(p_input[11627]), .Z(n18608) );
  AND U27912 ( .A(p_input[31627]), .B(p_input[21627]), .Z(n18607) );
  AND U27913 ( .A(n18609), .B(n18610), .Z(o[1626]) );
  AND U27914 ( .A(p_input[1626]), .B(p_input[11626]), .Z(n18610) );
  AND U27915 ( .A(p_input[31626]), .B(p_input[21626]), .Z(n18609) );
  AND U27916 ( .A(n18611), .B(n18612), .Z(o[1625]) );
  AND U27917 ( .A(p_input[1625]), .B(p_input[11625]), .Z(n18612) );
  AND U27918 ( .A(p_input[31625]), .B(p_input[21625]), .Z(n18611) );
  AND U27919 ( .A(n18613), .B(n18614), .Z(o[1624]) );
  AND U27920 ( .A(p_input[1624]), .B(p_input[11624]), .Z(n18614) );
  AND U27921 ( .A(p_input[31624]), .B(p_input[21624]), .Z(n18613) );
  AND U27922 ( .A(n18615), .B(n18616), .Z(o[1623]) );
  AND U27923 ( .A(p_input[1623]), .B(p_input[11623]), .Z(n18616) );
  AND U27924 ( .A(p_input[31623]), .B(p_input[21623]), .Z(n18615) );
  AND U27925 ( .A(n18617), .B(n18618), .Z(o[1622]) );
  AND U27926 ( .A(p_input[1622]), .B(p_input[11622]), .Z(n18618) );
  AND U27927 ( .A(p_input[31622]), .B(p_input[21622]), .Z(n18617) );
  AND U27928 ( .A(n18619), .B(n18620), .Z(o[1621]) );
  AND U27929 ( .A(p_input[1621]), .B(p_input[11621]), .Z(n18620) );
  AND U27930 ( .A(p_input[31621]), .B(p_input[21621]), .Z(n18619) );
  AND U27931 ( .A(n18621), .B(n18622), .Z(o[1620]) );
  AND U27932 ( .A(p_input[1620]), .B(p_input[11620]), .Z(n18622) );
  AND U27933 ( .A(p_input[31620]), .B(p_input[21620]), .Z(n18621) );
  AND U27934 ( .A(n18623), .B(n18624), .Z(o[161]) );
  AND U27935 ( .A(p_input[161]), .B(p_input[10161]), .Z(n18624) );
  AND U27936 ( .A(p_input[30161]), .B(p_input[20161]), .Z(n18623) );
  AND U27937 ( .A(n18625), .B(n18626), .Z(o[1619]) );
  AND U27938 ( .A(p_input[1619]), .B(p_input[11619]), .Z(n18626) );
  AND U27939 ( .A(p_input[31619]), .B(p_input[21619]), .Z(n18625) );
  AND U27940 ( .A(n18627), .B(n18628), .Z(o[1618]) );
  AND U27941 ( .A(p_input[1618]), .B(p_input[11618]), .Z(n18628) );
  AND U27942 ( .A(p_input[31618]), .B(p_input[21618]), .Z(n18627) );
  AND U27943 ( .A(n18629), .B(n18630), .Z(o[1617]) );
  AND U27944 ( .A(p_input[1617]), .B(p_input[11617]), .Z(n18630) );
  AND U27945 ( .A(p_input[31617]), .B(p_input[21617]), .Z(n18629) );
  AND U27946 ( .A(n18631), .B(n18632), .Z(o[1616]) );
  AND U27947 ( .A(p_input[1616]), .B(p_input[11616]), .Z(n18632) );
  AND U27948 ( .A(p_input[31616]), .B(p_input[21616]), .Z(n18631) );
  AND U27949 ( .A(n18633), .B(n18634), .Z(o[1615]) );
  AND U27950 ( .A(p_input[1615]), .B(p_input[11615]), .Z(n18634) );
  AND U27951 ( .A(p_input[31615]), .B(p_input[21615]), .Z(n18633) );
  AND U27952 ( .A(n18635), .B(n18636), .Z(o[1614]) );
  AND U27953 ( .A(p_input[1614]), .B(p_input[11614]), .Z(n18636) );
  AND U27954 ( .A(p_input[31614]), .B(p_input[21614]), .Z(n18635) );
  AND U27955 ( .A(n18637), .B(n18638), .Z(o[1613]) );
  AND U27956 ( .A(p_input[1613]), .B(p_input[11613]), .Z(n18638) );
  AND U27957 ( .A(p_input[31613]), .B(p_input[21613]), .Z(n18637) );
  AND U27958 ( .A(n18639), .B(n18640), .Z(o[1612]) );
  AND U27959 ( .A(p_input[1612]), .B(p_input[11612]), .Z(n18640) );
  AND U27960 ( .A(p_input[31612]), .B(p_input[21612]), .Z(n18639) );
  AND U27961 ( .A(n18641), .B(n18642), .Z(o[1611]) );
  AND U27962 ( .A(p_input[1611]), .B(p_input[11611]), .Z(n18642) );
  AND U27963 ( .A(p_input[31611]), .B(p_input[21611]), .Z(n18641) );
  AND U27964 ( .A(n18643), .B(n18644), .Z(o[1610]) );
  AND U27965 ( .A(p_input[1610]), .B(p_input[11610]), .Z(n18644) );
  AND U27966 ( .A(p_input[31610]), .B(p_input[21610]), .Z(n18643) );
  AND U27967 ( .A(n18645), .B(n18646), .Z(o[160]) );
  AND U27968 ( .A(p_input[160]), .B(p_input[10160]), .Z(n18646) );
  AND U27969 ( .A(p_input[30160]), .B(p_input[20160]), .Z(n18645) );
  AND U27970 ( .A(n18647), .B(n18648), .Z(o[1609]) );
  AND U27971 ( .A(p_input[1609]), .B(p_input[11609]), .Z(n18648) );
  AND U27972 ( .A(p_input[31609]), .B(p_input[21609]), .Z(n18647) );
  AND U27973 ( .A(n18649), .B(n18650), .Z(o[1608]) );
  AND U27974 ( .A(p_input[1608]), .B(p_input[11608]), .Z(n18650) );
  AND U27975 ( .A(p_input[31608]), .B(p_input[21608]), .Z(n18649) );
  AND U27976 ( .A(n18651), .B(n18652), .Z(o[1607]) );
  AND U27977 ( .A(p_input[1607]), .B(p_input[11607]), .Z(n18652) );
  AND U27978 ( .A(p_input[31607]), .B(p_input[21607]), .Z(n18651) );
  AND U27979 ( .A(n18653), .B(n18654), .Z(o[1606]) );
  AND U27980 ( .A(p_input[1606]), .B(p_input[11606]), .Z(n18654) );
  AND U27981 ( .A(p_input[31606]), .B(p_input[21606]), .Z(n18653) );
  AND U27982 ( .A(n18655), .B(n18656), .Z(o[1605]) );
  AND U27983 ( .A(p_input[1605]), .B(p_input[11605]), .Z(n18656) );
  AND U27984 ( .A(p_input[31605]), .B(p_input[21605]), .Z(n18655) );
  AND U27985 ( .A(n18657), .B(n18658), .Z(o[1604]) );
  AND U27986 ( .A(p_input[1604]), .B(p_input[11604]), .Z(n18658) );
  AND U27987 ( .A(p_input[31604]), .B(p_input[21604]), .Z(n18657) );
  AND U27988 ( .A(n18659), .B(n18660), .Z(o[1603]) );
  AND U27989 ( .A(p_input[1603]), .B(p_input[11603]), .Z(n18660) );
  AND U27990 ( .A(p_input[31603]), .B(p_input[21603]), .Z(n18659) );
  AND U27991 ( .A(n18661), .B(n18662), .Z(o[1602]) );
  AND U27992 ( .A(p_input[1602]), .B(p_input[11602]), .Z(n18662) );
  AND U27993 ( .A(p_input[31602]), .B(p_input[21602]), .Z(n18661) );
  AND U27994 ( .A(n18663), .B(n18664), .Z(o[1601]) );
  AND U27995 ( .A(p_input[1601]), .B(p_input[11601]), .Z(n18664) );
  AND U27996 ( .A(p_input[31601]), .B(p_input[21601]), .Z(n18663) );
  AND U27997 ( .A(n18665), .B(n18666), .Z(o[1600]) );
  AND U27998 ( .A(p_input[1600]), .B(p_input[11600]), .Z(n18666) );
  AND U27999 ( .A(p_input[31600]), .B(p_input[21600]), .Z(n18665) );
  AND U28000 ( .A(n18667), .B(n18668), .Z(o[15]) );
  AND U28001 ( .A(p_input[15]), .B(p_input[10015]), .Z(n18668) );
  AND U28002 ( .A(p_input[30015]), .B(p_input[20015]), .Z(n18667) );
  AND U28003 ( .A(n18669), .B(n18670), .Z(o[159]) );
  AND U28004 ( .A(p_input[159]), .B(p_input[10159]), .Z(n18670) );
  AND U28005 ( .A(p_input[30159]), .B(p_input[20159]), .Z(n18669) );
  AND U28006 ( .A(n18671), .B(n18672), .Z(o[1599]) );
  AND U28007 ( .A(p_input[1599]), .B(p_input[11599]), .Z(n18672) );
  AND U28008 ( .A(p_input[31599]), .B(p_input[21599]), .Z(n18671) );
  AND U28009 ( .A(n18673), .B(n18674), .Z(o[1598]) );
  AND U28010 ( .A(p_input[1598]), .B(p_input[11598]), .Z(n18674) );
  AND U28011 ( .A(p_input[31598]), .B(p_input[21598]), .Z(n18673) );
  AND U28012 ( .A(n18675), .B(n18676), .Z(o[1597]) );
  AND U28013 ( .A(p_input[1597]), .B(p_input[11597]), .Z(n18676) );
  AND U28014 ( .A(p_input[31597]), .B(p_input[21597]), .Z(n18675) );
  AND U28015 ( .A(n18677), .B(n18678), .Z(o[1596]) );
  AND U28016 ( .A(p_input[1596]), .B(p_input[11596]), .Z(n18678) );
  AND U28017 ( .A(p_input[31596]), .B(p_input[21596]), .Z(n18677) );
  AND U28018 ( .A(n18679), .B(n18680), .Z(o[1595]) );
  AND U28019 ( .A(p_input[1595]), .B(p_input[11595]), .Z(n18680) );
  AND U28020 ( .A(p_input[31595]), .B(p_input[21595]), .Z(n18679) );
  AND U28021 ( .A(n18681), .B(n18682), .Z(o[1594]) );
  AND U28022 ( .A(p_input[1594]), .B(p_input[11594]), .Z(n18682) );
  AND U28023 ( .A(p_input[31594]), .B(p_input[21594]), .Z(n18681) );
  AND U28024 ( .A(n18683), .B(n18684), .Z(o[1593]) );
  AND U28025 ( .A(p_input[1593]), .B(p_input[11593]), .Z(n18684) );
  AND U28026 ( .A(p_input[31593]), .B(p_input[21593]), .Z(n18683) );
  AND U28027 ( .A(n18685), .B(n18686), .Z(o[1592]) );
  AND U28028 ( .A(p_input[1592]), .B(p_input[11592]), .Z(n18686) );
  AND U28029 ( .A(p_input[31592]), .B(p_input[21592]), .Z(n18685) );
  AND U28030 ( .A(n18687), .B(n18688), .Z(o[1591]) );
  AND U28031 ( .A(p_input[1591]), .B(p_input[11591]), .Z(n18688) );
  AND U28032 ( .A(p_input[31591]), .B(p_input[21591]), .Z(n18687) );
  AND U28033 ( .A(n18689), .B(n18690), .Z(o[1590]) );
  AND U28034 ( .A(p_input[1590]), .B(p_input[11590]), .Z(n18690) );
  AND U28035 ( .A(p_input[31590]), .B(p_input[21590]), .Z(n18689) );
  AND U28036 ( .A(n18691), .B(n18692), .Z(o[158]) );
  AND U28037 ( .A(p_input[158]), .B(p_input[10158]), .Z(n18692) );
  AND U28038 ( .A(p_input[30158]), .B(p_input[20158]), .Z(n18691) );
  AND U28039 ( .A(n18693), .B(n18694), .Z(o[1589]) );
  AND U28040 ( .A(p_input[1589]), .B(p_input[11589]), .Z(n18694) );
  AND U28041 ( .A(p_input[31589]), .B(p_input[21589]), .Z(n18693) );
  AND U28042 ( .A(n18695), .B(n18696), .Z(o[1588]) );
  AND U28043 ( .A(p_input[1588]), .B(p_input[11588]), .Z(n18696) );
  AND U28044 ( .A(p_input[31588]), .B(p_input[21588]), .Z(n18695) );
  AND U28045 ( .A(n18697), .B(n18698), .Z(o[1587]) );
  AND U28046 ( .A(p_input[1587]), .B(p_input[11587]), .Z(n18698) );
  AND U28047 ( .A(p_input[31587]), .B(p_input[21587]), .Z(n18697) );
  AND U28048 ( .A(n18699), .B(n18700), .Z(o[1586]) );
  AND U28049 ( .A(p_input[1586]), .B(p_input[11586]), .Z(n18700) );
  AND U28050 ( .A(p_input[31586]), .B(p_input[21586]), .Z(n18699) );
  AND U28051 ( .A(n18701), .B(n18702), .Z(o[1585]) );
  AND U28052 ( .A(p_input[1585]), .B(p_input[11585]), .Z(n18702) );
  AND U28053 ( .A(p_input[31585]), .B(p_input[21585]), .Z(n18701) );
  AND U28054 ( .A(n18703), .B(n18704), .Z(o[1584]) );
  AND U28055 ( .A(p_input[1584]), .B(p_input[11584]), .Z(n18704) );
  AND U28056 ( .A(p_input[31584]), .B(p_input[21584]), .Z(n18703) );
  AND U28057 ( .A(n18705), .B(n18706), .Z(o[1583]) );
  AND U28058 ( .A(p_input[1583]), .B(p_input[11583]), .Z(n18706) );
  AND U28059 ( .A(p_input[31583]), .B(p_input[21583]), .Z(n18705) );
  AND U28060 ( .A(n18707), .B(n18708), .Z(o[1582]) );
  AND U28061 ( .A(p_input[1582]), .B(p_input[11582]), .Z(n18708) );
  AND U28062 ( .A(p_input[31582]), .B(p_input[21582]), .Z(n18707) );
  AND U28063 ( .A(n18709), .B(n18710), .Z(o[1581]) );
  AND U28064 ( .A(p_input[1581]), .B(p_input[11581]), .Z(n18710) );
  AND U28065 ( .A(p_input[31581]), .B(p_input[21581]), .Z(n18709) );
  AND U28066 ( .A(n18711), .B(n18712), .Z(o[1580]) );
  AND U28067 ( .A(p_input[1580]), .B(p_input[11580]), .Z(n18712) );
  AND U28068 ( .A(p_input[31580]), .B(p_input[21580]), .Z(n18711) );
  AND U28069 ( .A(n18713), .B(n18714), .Z(o[157]) );
  AND U28070 ( .A(p_input[157]), .B(p_input[10157]), .Z(n18714) );
  AND U28071 ( .A(p_input[30157]), .B(p_input[20157]), .Z(n18713) );
  AND U28072 ( .A(n18715), .B(n18716), .Z(o[1579]) );
  AND U28073 ( .A(p_input[1579]), .B(p_input[11579]), .Z(n18716) );
  AND U28074 ( .A(p_input[31579]), .B(p_input[21579]), .Z(n18715) );
  AND U28075 ( .A(n18717), .B(n18718), .Z(o[1578]) );
  AND U28076 ( .A(p_input[1578]), .B(p_input[11578]), .Z(n18718) );
  AND U28077 ( .A(p_input[31578]), .B(p_input[21578]), .Z(n18717) );
  AND U28078 ( .A(n18719), .B(n18720), .Z(o[1577]) );
  AND U28079 ( .A(p_input[1577]), .B(p_input[11577]), .Z(n18720) );
  AND U28080 ( .A(p_input[31577]), .B(p_input[21577]), .Z(n18719) );
  AND U28081 ( .A(n18721), .B(n18722), .Z(o[1576]) );
  AND U28082 ( .A(p_input[1576]), .B(p_input[11576]), .Z(n18722) );
  AND U28083 ( .A(p_input[31576]), .B(p_input[21576]), .Z(n18721) );
  AND U28084 ( .A(n18723), .B(n18724), .Z(o[1575]) );
  AND U28085 ( .A(p_input[1575]), .B(p_input[11575]), .Z(n18724) );
  AND U28086 ( .A(p_input[31575]), .B(p_input[21575]), .Z(n18723) );
  AND U28087 ( .A(n18725), .B(n18726), .Z(o[1574]) );
  AND U28088 ( .A(p_input[1574]), .B(p_input[11574]), .Z(n18726) );
  AND U28089 ( .A(p_input[31574]), .B(p_input[21574]), .Z(n18725) );
  AND U28090 ( .A(n18727), .B(n18728), .Z(o[1573]) );
  AND U28091 ( .A(p_input[1573]), .B(p_input[11573]), .Z(n18728) );
  AND U28092 ( .A(p_input[31573]), .B(p_input[21573]), .Z(n18727) );
  AND U28093 ( .A(n18729), .B(n18730), .Z(o[1572]) );
  AND U28094 ( .A(p_input[1572]), .B(p_input[11572]), .Z(n18730) );
  AND U28095 ( .A(p_input[31572]), .B(p_input[21572]), .Z(n18729) );
  AND U28096 ( .A(n18731), .B(n18732), .Z(o[1571]) );
  AND U28097 ( .A(p_input[1571]), .B(p_input[11571]), .Z(n18732) );
  AND U28098 ( .A(p_input[31571]), .B(p_input[21571]), .Z(n18731) );
  AND U28099 ( .A(n18733), .B(n18734), .Z(o[1570]) );
  AND U28100 ( .A(p_input[1570]), .B(p_input[11570]), .Z(n18734) );
  AND U28101 ( .A(p_input[31570]), .B(p_input[21570]), .Z(n18733) );
  AND U28102 ( .A(n18735), .B(n18736), .Z(o[156]) );
  AND U28103 ( .A(p_input[156]), .B(p_input[10156]), .Z(n18736) );
  AND U28104 ( .A(p_input[30156]), .B(p_input[20156]), .Z(n18735) );
  AND U28105 ( .A(n18737), .B(n18738), .Z(o[1569]) );
  AND U28106 ( .A(p_input[1569]), .B(p_input[11569]), .Z(n18738) );
  AND U28107 ( .A(p_input[31569]), .B(p_input[21569]), .Z(n18737) );
  AND U28108 ( .A(n18739), .B(n18740), .Z(o[1568]) );
  AND U28109 ( .A(p_input[1568]), .B(p_input[11568]), .Z(n18740) );
  AND U28110 ( .A(p_input[31568]), .B(p_input[21568]), .Z(n18739) );
  AND U28111 ( .A(n18741), .B(n18742), .Z(o[1567]) );
  AND U28112 ( .A(p_input[1567]), .B(p_input[11567]), .Z(n18742) );
  AND U28113 ( .A(p_input[31567]), .B(p_input[21567]), .Z(n18741) );
  AND U28114 ( .A(n18743), .B(n18744), .Z(o[1566]) );
  AND U28115 ( .A(p_input[1566]), .B(p_input[11566]), .Z(n18744) );
  AND U28116 ( .A(p_input[31566]), .B(p_input[21566]), .Z(n18743) );
  AND U28117 ( .A(n18745), .B(n18746), .Z(o[1565]) );
  AND U28118 ( .A(p_input[1565]), .B(p_input[11565]), .Z(n18746) );
  AND U28119 ( .A(p_input[31565]), .B(p_input[21565]), .Z(n18745) );
  AND U28120 ( .A(n18747), .B(n18748), .Z(o[1564]) );
  AND U28121 ( .A(p_input[1564]), .B(p_input[11564]), .Z(n18748) );
  AND U28122 ( .A(p_input[31564]), .B(p_input[21564]), .Z(n18747) );
  AND U28123 ( .A(n18749), .B(n18750), .Z(o[1563]) );
  AND U28124 ( .A(p_input[1563]), .B(p_input[11563]), .Z(n18750) );
  AND U28125 ( .A(p_input[31563]), .B(p_input[21563]), .Z(n18749) );
  AND U28126 ( .A(n18751), .B(n18752), .Z(o[1562]) );
  AND U28127 ( .A(p_input[1562]), .B(p_input[11562]), .Z(n18752) );
  AND U28128 ( .A(p_input[31562]), .B(p_input[21562]), .Z(n18751) );
  AND U28129 ( .A(n18753), .B(n18754), .Z(o[1561]) );
  AND U28130 ( .A(p_input[1561]), .B(p_input[11561]), .Z(n18754) );
  AND U28131 ( .A(p_input[31561]), .B(p_input[21561]), .Z(n18753) );
  AND U28132 ( .A(n18755), .B(n18756), .Z(o[1560]) );
  AND U28133 ( .A(p_input[1560]), .B(p_input[11560]), .Z(n18756) );
  AND U28134 ( .A(p_input[31560]), .B(p_input[21560]), .Z(n18755) );
  AND U28135 ( .A(n18757), .B(n18758), .Z(o[155]) );
  AND U28136 ( .A(p_input[155]), .B(p_input[10155]), .Z(n18758) );
  AND U28137 ( .A(p_input[30155]), .B(p_input[20155]), .Z(n18757) );
  AND U28138 ( .A(n18759), .B(n18760), .Z(o[1559]) );
  AND U28139 ( .A(p_input[1559]), .B(p_input[11559]), .Z(n18760) );
  AND U28140 ( .A(p_input[31559]), .B(p_input[21559]), .Z(n18759) );
  AND U28141 ( .A(n18761), .B(n18762), .Z(o[1558]) );
  AND U28142 ( .A(p_input[1558]), .B(p_input[11558]), .Z(n18762) );
  AND U28143 ( .A(p_input[31558]), .B(p_input[21558]), .Z(n18761) );
  AND U28144 ( .A(n18763), .B(n18764), .Z(o[1557]) );
  AND U28145 ( .A(p_input[1557]), .B(p_input[11557]), .Z(n18764) );
  AND U28146 ( .A(p_input[31557]), .B(p_input[21557]), .Z(n18763) );
  AND U28147 ( .A(n18765), .B(n18766), .Z(o[1556]) );
  AND U28148 ( .A(p_input[1556]), .B(p_input[11556]), .Z(n18766) );
  AND U28149 ( .A(p_input[31556]), .B(p_input[21556]), .Z(n18765) );
  AND U28150 ( .A(n18767), .B(n18768), .Z(o[1555]) );
  AND U28151 ( .A(p_input[1555]), .B(p_input[11555]), .Z(n18768) );
  AND U28152 ( .A(p_input[31555]), .B(p_input[21555]), .Z(n18767) );
  AND U28153 ( .A(n18769), .B(n18770), .Z(o[1554]) );
  AND U28154 ( .A(p_input[1554]), .B(p_input[11554]), .Z(n18770) );
  AND U28155 ( .A(p_input[31554]), .B(p_input[21554]), .Z(n18769) );
  AND U28156 ( .A(n18771), .B(n18772), .Z(o[1553]) );
  AND U28157 ( .A(p_input[1553]), .B(p_input[11553]), .Z(n18772) );
  AND U28158 ( .A(p_input[31553]), .B(p_input[21553]), .Z(n18771) );
  AND U28159 ( .A(n18773), .B(n18774), .Z(o[1552]) );
  AND U28160 ( .A(p_input[1552]), .B(p_input[11552]), .Z(n18774) );
  AND U28161 ( .A(p_input[31552]), .B(p_input[21552]), .Z(n18773) );
  AND U28162 ( .A(n18775), .B(n18776), .Z(o[1551]) );
  AND U28163 ( .A(p_input[1551]), .B(p_input[11551]), .Z(n18776) );
  AND U28164 ( .A(p_input[31551]), .B(p_input[21551]), .Z(n18775) );
  AND U28165 ( .A(n18777), .B(n18778), .Z(o[1550]) );
  AND U28166 ( .A(p_input[1550]), .B(p_input[11550]), .Z(n18778) );
  AND U28167 ( .A(p_input[31550]), .B(p_input[21550]), .Z(n18777) );
  AND U28168 ( .A(n18779), .B(n18780), .Z(o[154]) );
  AND U28169 ( .A(p_input[154]), .B(p_input[10154]), .Z(n18780) );
  AND U28170 ( .A(p_input[30154]), .B(p_input[20154]), .Z(n18779) );
  AND U28171 ( .A(n18781), .B(n18782), .Z(o[1549]) );
  AND U28172 ( .A(p_input[1549]), .B(p_input[11549]), .Z(n18782) );
  AND U28173 ( .A(p_input[31549]), .B(p_input[21549]), .Z(n18781) );
  AND U28174 ( .A(n18783), .B(n18784), .Z(o[1548]) );
  AND U28175 ( .A(p_input[1548]), .B(p_input[11548]), .Z(n18784) );
  AND U28176 ( .A(p_input[31548]), .B(p_input[21548]), .Z(n18783) );
  AND U28177 ( .A(n18785), .B(n18786), .Z(o[1547]) );
  AND U28178 ( .A(p_input[1547]), .B(p_input[11547]), .Z(n18786) );
  AND U28179 ( .A(p_input[31547]), .B(p_input[21547]), .Z(n18785) );
  AND U28180 ( .A(n18787), .B(n18788), .Z(o[1546]) );
  AND U28181 ( .A(p_input[1546]), .B(p_input[11546]), .Z(n18788) );
  AND U28182 ( .A(p_input[31546]), .B(p_input[21546]), .Z(n18787) );
  AND U28183 ( .A(n18789), .B(n18790), .Z(o[1545]) );
  AND U28184 ( .A(p_input[1545]), .B(p_input[11545]), .Z(n18790) );
  AND U28185 ( .A(p_input[31545]), .B(p_input[21545]), .Z(n18789) );
  AND U28186 ( .A(n18791), .B(n18792), .Z(o[1544]) );
  AND U28187 ( .A(p_input[1544]), .B(p_input[11544]), .Z(n18792) );
  AND U28188 ( .A(p_input[31544]), .B(p_input[21544]), .Z(n18791) );
  AND U28189 ( .A(n18793), .B(n18794), .Z(o[1543]) );
  AND U28190 ( .A(p_input[1543]), .B(p_input[11543]), .Z(n18794) );
  AND U28191 ( .A(p_input[31543]), .B(p_input[21543]), .Z(n18793) );
  AND U28192 ( .A(n18795), .B(n18796), .Z(o[1542]) );
  AND U28193 ( .A(p_input[1542]), .B(p_input[11542]), .Z(n18796) );
  AND U28194 ( .A(p_input[31542]), .B(p_input[21542]), .Z(n18795) );
  AND U28195 ( .A(n18797), .B(n18798), .Z(o[1541]) );
  AND U28196 ( .A(p_input[1541]), .B(p_input[11541]), .Z(n18798) );
  AND U28197 ( .A(p_input[31541]), .B(p_input[21541]), .Z(n18797) );
  AND U28198 ( .A(n18799), .B(n18800), .Z(o[1540]) );
  AND U28199 ( .A(p_input[1540]), .B(p_input[11540]), .Z(n18800) );
  AND U28200 ( .A(p_input[31540]), .B(p_input[21540]), .Z(n18799) );
  AND U28201 ( .A(n18801), .B(n18802), .Z(o[153]) );
  AND U28202 ( .A(p_input[153]), .B(p_input[10153]), .Z(n18802) );
  AND U28203 ( .A(p_input[30153]), .B(p_input[20153]), .Z(n18801) );
  AND U28204 ( .A(n18803), .B(n18804), .Z(o[1539]) );
  AND U28205 ( .A(p_input[1539]), .B(p_input[11539]), .Z(n18804) );
  AND U28206 ( .A(p_input[31539]), .B(p_input[21539]), .Z(n18803) );
  AND U28207 ( .A(n18805), .B(n18806), .Z(o[1538]) );
  AND U28208 ( .A(p_input[1538]), .B(p_input[11538]), .Z(n18806) );
  AND U28209 ( .A(p_input[31538]), .B(p_input[21538]), .Z(n18805) );
  AND U28210 ( .A(n18807), .B(n18808), .Z(o[1537]) );
  AND U28211 ( .A(p_input[1537]), .B(p_input[11537]), .Z(n18808) );
  AND U28212 ( .A(p_input[31537]), .B(p_input[21537]), .Z(n18807) );
  AND U28213 ( .A(n18809), .B(n18810), .Z(o[1536]) );
  AND U28214 ( .A(p_input[1536]), .B(p_input[11536]), .Z(n18810) );
  AND U28215 ( .A(p_input[31536]), .B(p_input[21536]), .Z(n18809) );
  AND U28216 ( .A(n18811), .B(n18812), .Z(o[1535]) );
  AND U28217 ( .A(p_input[1535]), .B(p_input[11535]), .Z(n18812) );
  AND U28218 ( .A(p_input[31535]), .B(p_input[21535]), .Z(n18811) );
  AND U28219 ( .A(n18813), .B(n18814), .Z(o[1534]) );
  AND U28220 ( .A(p_input[1534]), .B(p_input[11534]), .Z(n18814) );
  AND U28221 ( .A(p_input[31534]), .B(p_input[21534]), .Z(n18813) );
  AND U28222 ( .A(n18815), .B(n18816), .Z(o[1533]) );
  AND U28223 ( .A(p_input[1533]), .B(p_input[11533]), .Z(n18816) );
  AND U28224 ( .A(p_input[31533]), .B(p_input[21533]), .Z(n18815) );
  AND U28225 ( .A(n18817), .B(n18818), .Z(o[1532]) );
  AND U28226 ( .A(p_input[1532]), .B(p_input[11532]), .Z(n18818) );
  AND U28227 ( .A(p_input[31532]), .B(p_input[21532]), .Z(n18817) );
  AND U28228 ( .A(n18819), .B(n18820), .Z(o[1531]) );
  AND U28229 ( .A(p_input[1531]), .B(p_input[11531]), .Z(n18820) );
  AND U28230 ( .A(p_input[31531]), .B(p_input[21531]), .Z(n18819) );
  AND U28231 ( .A(n18821), .B(n18822), .Z(o[1530]) );
  AND U28232 ( .A(p_input[1530]), .B(p_input[11530]), .Z(n18822) );
  AND U28233 ( .A(p_input[31530]), .B(p_input[21530]), .Z(n18821) );
  AND U28234 ( .A(n18823), .B(n18824), .Z(o[152]) );
  AND U28235 ( .A(p_input[152]), .B(p_input[10152]), .Z(n18824) );
  AND U28236 ( .A(p_input[30152]), .B(p_input[20152]), .Z(n18823) );
  AND U28237 ( .A(n18825), .B(n18826), .Z(o[1529]) );
  AND U28238 ( .A(p_input[1529]), .B(p_input[11529]), .Z(n18826) );
  AND U28239 ( .A(p_input[31529]), .B(p_input[21529]), .Z(n18825) );
  AND U28240 ( .A(n18827), .B(n18828), .Z(o[1528]) );
  AND U28241 ( .A(p_input[1528]), .B(p_input[11528]), .Z(n18828) );
  AND U28242 ( .A(p_input[31528]), .B(p_input[21528]), .Z(n18827) );
  AND U28243 ( .A(n18829), .B(n18830), .Z(o[1527]) );
  AND U28244 ( .A(p_input[1527]), .B(p_input[11527]), .Z(n18830) );
  AND U28245 ( .A(p_input[31527]), .B(p_input[21527]), .Z(n18829) );
  AND U28246 ( .A(n18831), .B(n18832), .Z(o[1526]) );
  AND U28247 ( .A(p_input[1526]), .B(p_input[11526]), .Z(n18832) );
  AND U28248 ( .A(p_input[31526]), .B(p_input[21526]), .Z(n18831) );
  AND U28249 ( .A(n18833), .B(n18834), .Z(o[1525]) );
  AND U28250 ( .A(p_input[1525]), .B(p_input[11525]), .Z(n18834) );
  AND U28251 ( .A(p_input[31525]), .B(p_input[21525]), .Z(n18833) );
  AND U28252 ( .A(n18835), .B(n18836), .Z(o[1524]) );
  AND U28253 ( .A(p_input[1524]), .B(p_input[11524]), .Z(n18836) );
  AND U28254 ( .A(p_input[31524]), .B(p_input[21524]), .Z(n18835) );
  AND U28255 ( .A(n18837), .B(n18838), .Z(o[1523]) );
  AND U28256 ( .A(p_input[1523]), .B(p_input[11523]), .Z(n18838) );
  AND U28257 ( .A(p_input[31523]), .B(p_input[21523]), .Z(n18837) );
  AND U28258 ( .A(n18839), .B(n18840), .Z(o[1522]) );
  AND U28259 ( .A(p_input[1522]), .B(p_input[11522]), .Z(n18840) );
  AND U28260 ( .A(p_input[31522]), .B(p_input[21522]), .Z(n18839) );
  AND U28261 ( .A(n18841), .B(n18842), .Z(o[1521]) );
  AND U28262 ( .A(p_input[1521]), .B(p_input[11521]), .Z(n18842) );
  AND U28263 ( .A(p_input[31521]), .B(p_input[21521]), .Z(n18841) );
  AND U28264 ( .A(n18843), .B(n18844), .Z(o[1520]) );
  AND U28265 ( .A(p_input[1520]), .B(p_input[11520]), .Z(n18844) );
  AND U28266 ( .A(p_input[31520]), .B(p_input[21520]), .Z(n18843) );
  AND U28267 ( .A(n18845), .B(n18846), .Z(o[151]) );
  AND U28268 ( .A(p_input[151]), .B(p_input[10151]), .Z(n18846) );
  AND U28269 ( .A(p_input[30151]), .B(p_input[20151]), .Z(n18845) );
  AND U28270 ( .A(n18847), .B(n18848), .Z(o[1519]) );
  AND U28271 ( .A(p_input[1519]), .B(p_input[11519]), .Z(n18848) );
  AND U28272 ( .A(p_input[31519]), .B(p_input[21519]), .Z(n18847) );
  AND U28273 ( .A(n18849), .B(n18850), .Z(o[1518]) );
  AND U28274 ( .A(p_input[1518]), .B(p_input[11518]), .Z(n18850) );
  AND U28275 ( .A(p_input[31518]), .B(p_input[21518]), .Z(n18849) );
  AND U28276 ( .A(n18851), .B(n18852), .Z(o[1517]) );
  AND U28277 ( .A(p_input[1517]), .B(p_input[11517]), .Z(n18852) );
  AND U28278 ( .A(p_input[31517]), .B(p_input[21517]), .Z(n18851) );
  AND U28279 ( .A(n18853), .B(n18854), .Z(o[1516]) );
  AND U28280 ( .A(p_input[1516]), .B(p_input[11516]), .Z(n18854) );
  AND U28281 ( .A(p_input[31516]), .B(p_input[21516]), .Z(n18853) );
  AND U28282 ( .A(n18855), .B(n18856), .Z(o[1515]) );
  AND U28283 ( .A(p_input[1515]), .B(p_input[11515]), .Z(n18856) );
  AND U28284 ( .A(p_input[31515]), .B(p_input[21515]), .Z(n18855) );
  AND U28285 ( .A(n18857), .B(n18858), .Z(o[1514]) );
  AND U28286 ( .A(p_input[1514]), .B(p_input[11514]), .Z(n18858) );
  AND U28287 ( .A(p_input[31514]), .B(p_input[21514]), .Z(n18857) );
  AND U28288 ( .A(n18859), .B(n18860), .Z(o[1513]) );
  AND U28289 ( .A(p_input[1513]), .B(p_input[11513]), .Z(n18860) );
  AND U28290 ( .A(p_input[31513]), .B(p_input[21513]), .Z(n18859) );
  AND U28291 ( .A(n18861), .B(n18862), .Z(o[1512]) );
  AND U28292 ( .A(p_input[1512]), .B(p_input[11512]), .Z(n18862) );
  AND U28293 ( .A(p_input[31512]), .B(p_input[21512]), .Z(n18861) );
  AND U28294 ( .A(n18863), .B(n18864), .Z(o[1511]) );
  AND U28295 ( .A(p_input[1511]), .B(p_input[11511]), .Z(n18864) );
  AND U28296 ( .A(p_input[31511]), .B(p_input[21511]), .Z(n18863) );
  AND U28297 ( .A(n18865), .B(n18866), .Z(o[1510]) );
  AND U28298 ( .A(p_input[1510]), .B(p_input[11510]), .Z(n18866) );
  AND U28299 ( .A(p_input[31510]), .B(p_input[21510]), .Z(n18865) );
  AND U28300 ( .A(n18867), .B(n18868), .Z(o[150]) );
  AND U28301 ( .A(p_input[150]), .B(p_input[10150]), .Z(n18868) );
  AND U28302 ( .A(p_input[30150]), .B(p_input[20150]), .Z(n18867) );
  AND U28303 ( .A(n18869), .B(n18870), .Z(o[1509]) );
  AND U28304 ( .A(p_input[1509]), .B(p_input[11509]), .Z(n18870) );
  AND U28305 ( .A(p_input[31509]), .B(p_input[21509]), .Z(n18869) );
  AND U28306 ( .A(n18871), .B(n18872), .Z(o[1508]) );
  AND U28307 ( .A(p_input[1508]), .B(p_input[11508]), .Z(n18872) );
  AND U28308 ( .A(p_input[31508]), .B(p_input[21508]), .Z(n18871) );
  AND U28309 ( .A(n18873), .B(n18874), .Z(o[1507]) );
  AND U28310 ( .A(p_input[1507]), .B(p_input[11507]), .Z(n18874) );
  AND U28311 ( .A(p_input[31507]), .B(p_input[21507]), .Z(n18873) );
  AND U28312 ( .A(n18875), .B(n18876), .Z(o[1506]) );
  AND U28313 ( .A(p_input[1506]), .B(p_input[11506]), .Z(n18876) );
  AND U28314 ( .A(p_input[31506]), .B(p_input[21506]), .Z(n18875) );
  AND U28315 ( .A(n18877), .B(n18878), .Z(o[1505]) );
  AND U28316 ( .A(p_input[1505]), .B(p_input[11505]), .Z(n18878) );
  AND U28317 ( .A(p_input[31505]), .B(p_input[21505]), .Z(n18877) );
  AND U28318 ( .A(n18879), .B(n18880), .Z(o[1504]) );
  AND U28319 ( .A(p_input[1504]), .B(p_input[11504]), .Z(n18880) );
  AND U28320 ( .A(p_input[31504]), .B(p_input[21504]), .Z(n18879) );
  AND U28321 ( .A(n18881), .B(n18882), .Z(o[1503]) );
  AND U28322 ( .A(p_input[1503]), .B(p_input[11503]), .Z(n18882) );
  AND U28323 ( .A(p_input[31503]), .B(p_input[21503]), .Z(n18881) );
  AND U28324 ( .A(n18883), .B(n18884), .Z(o[1502]) );
  AND U28325 ( .A(p_input[1502]), .B(p_input[11502]), .Z(n18884) );
  AND U28326 ( .A(p_input[31502]), .B(p_input[21502]), .Z(n18883) );
  AND U28327 ( .A(n18885), .B(n18886), .Z(o[1501]) );
  AND U28328 ( .A(p_input[1501]), .B(p_input[11501]), .Z(n18886) );
  AND U28329 ( .A(p_input[31501]), .B(p_input[21501]), .Z(n18885) );
  AND U28330 ( .A(n18887), .B(n18888), .Z(o[1500]) );
  AND U28331 ( .A(p_input[1500]), .B(p_input[11500]), .Z(n18888) );
  AND U28332 ( .A(p_input[31500]), .B(p_input[21500]), .Z(n18887) );
  AND U28333 ( .A(n18889), .B(n18890), .Z(o[14]) );
  AND U28334 ( .A(p_input[14]), .B(p_input[10014]), .Z(n18890) );
  AND U28335 ( .A(p_input[30014]), .B(p_input[20014]), .Z(n18889) );
  AND U28336 ( .A(n18891), .B(n18892), .Z(o[149]) );
  AND U28337 ( .A(p_input[149]), .B(p_input[10149]), .Z(n18892) );
  AND U28338 ( .A(p_input[30149]), .B(p_input[20149]), .Z(n18891) );
  AND U28339 ( .A(n18893), .B(n18894), .Z(o[1499]) );
  AND U28340 ( .A(p_input[1499]), .B(p_input[11499]), .Z(n18894) );
  AND U28341 ( .A(p_input[31499]), .B(p_input[21499]), .Z(n18893) );
  AND U28342 ( .A(n18895), .B(n18896), .Z(o[1498]) );
  AND U28343 ( .A(p_input[1498]), .B(p_input[11498]), .Z(n18896) );
  AND U28344 ( .A(p_input[31498]), .B(p_input[21498]), .Z(n18895) );
  AND U28345 ( .A(n18897), .B(n18898), .Z(o[1497]) );
  AND U28346 ( .A(p_input[1497]), .B(p_input[11497]), .Z(n18898) );
  AND U28347 ( .A(p_input[31497]), .B(p_input[21497]), .Z(n18897) );
  AND U28348 ( .A(n18899), .B(n18900), .Z(o[1496]) );
  AND U28349 ( .A(p_input[1496]), .B(p_input[11496]), .Z(n18900) );
  AND U28350 ( .A(p_input[31496]), .B(p_input[21496]), .Z(n18899) );
  AND U28351 ( .A(n18901), .B(n18902), .Z(o[1495]) );
  AND U28352 ( .A(p_input[1495]), .B(p_input[11495]), .Z(n18902) );
  AND U28353 ( .A(p_input[31495]), .B(p_input[21495]), .Z(n18901) );
  AND U28354 ( .A(n18903), .B(n18904), .Z(o[1494]) );
  AND U28355 ( .A(p_input[1494]), .B(p_input[11494]), .Z(n18904) );
  AND U28356 ( .A(p_input[31494]), .B(p_input[21494]), .Z(n18903) );
  AND U28357 ( .A(n18905), .B(n18906), .Z(o[1493]) );
  AND U28358 ( .A(p_input[1493]), .B(p_input[11493]), .Z(n18906) );
  AND U28359 ( .A(p_input[31493]), .B(p_input[21493]), .Z(n18905) );
  AND U28360 ( .A(n18907), .B(n18908), .Z(o[1492]) );
  AND U28361 ( .A(p_input[1492]), .B(p_input[11492]), .Z(n18908) );
  AND U28362 ( .A(p_input[31492]), .B(p_input[21492]), .Z(n18907) );
  AND U28363 ( .A(n18909), .B(n18910), .Z(o[1491]) );
  AND U28364 ( .A(p_input[1491]), .B(p_input[11491]), .Z(n18910) );
  AND U28365 ( .A(p_input[31491]), .B(p_input[21491]), .Z(n18909) );
  AND U28366 ( .A(n18911), .B(n18912), .Z(o[1490]) );
  AND U28367 ( .A(p_input[1490]), .B(p_input[11490]), .Z(n18912) );
  AND U28368 ( .A(p_input[31490]), .B(p_input[21490]), .Z(n18911) );
  AND U28369 ( .A(n18913), .B(n18914), .Z(o[148]) );
  AND U28370 ( .A(p_input[148]), .B(p_input[10148]), .Z(n18914) );
  AND U28371 ( .A(p_input[30148]), .B(p_input[20148]), .Z(n18913) );
  AND U28372 ( .A(n18915), .B(n18916), .Z(o[1489]) );
  AND U28373 ( .A(p_input[1489]), .B(p_input[11489]), .Z(n18916) );
  AND U28374 ( .A(p_input[31489]), .B(p_input[21489]), .Z(n18915) );
  AND U28375 ( .A(n18917), .B(n18918), .Z(o[1488]) );
  AND U28376 ( .A(p_input[1488]), .B(p_input[11488]), .Z(n18918) );
  AND U28377 ( .A(p_input[31488]), .B(p_input[21488]), .Z(n18917) );
  AND U28378 ( .A(n18919), .B(n18920), .Z(o[1487]) );
  AND U28379 ( .A(p_input[1487]), .B(p_input[11487]), .Z(n18920) );
  AND U28380 ( .A(p_input[31487]), .B(p_input[21487]), .Z(n18919) );
  AND U28381 ( .A(n18921), .B(n18922), .Z(o[1486]) );
  AND U28382 ( .A(p_input[1486]), .B(p_input[11486]), .Z(n18922) );
  AND U28383 ( .A(p_input[31486]), .B(p_input[21486]), .Z(n18921) );
  AND U28384 ( .A(n18923), .B(n18924), .Z(o[1485]) );
  AND U28385 ( .A(p_input[1485]), .B(p_input[11485]), .Z(n18924) );
  AND U28386 ( .A(p_input[31485]), .B(p_input[21485]), .Z(n18923) );
  AND U28387 ( .A(n18925), .B(n18926), .Z(o[1484]) );
  AND U28388 ( .A(p_input[1484]), .B(p_input[11484]), .Z(n18926) );
  AND U28389 ( .A(p_input[31484]), .B(p_input[21484]), .Z(n18925) );
  AND U28390 ( .A(n18927), .B(n18928), .Z(o[1483]) );
  AND U28391 ( .A(p_input[1483]), .B(p_input[11483]), .Z(n18928) );
  AND U28392 ( .A(p_input[31483]), .B(p_input[21483]), .Z(n18927) );
  AND U28393 ( .A(n18929), .B(n18930), .Z(o[1482]) );
  AND U28394 ( .A(p_input[1482]), .B(p_input[11482]), .Z(n18930) );
  AND U28395 ( .A(p_input[31482]), .B(p_input[21482]), .Z(n18929) );
  AND U28396 ( .A(n18931), .B(n18932), .Z(o[1481]) );
  AND U28397 ( .A(p_input[1481]), .B(p_input[11481]), .Z(n18932) );
  AND U28398 ( .A(p_input[31481]), .B(p_input[21481]), .Z(n18931) );
  AND U28399 ( .A(n18933), .B(n18934), .Z(o[1480]) );
  AND U28400 ( .A(p_input[1480]), .B(p_input[11480]), .Z(n18934) );
  AND U28401 ( .A(p_input[31480]), .B(p_input[21480]), .Z(n18933) );
  AND U28402 ( .A(n18935), .B(n18936), .Z(o[147]) );
  AND U28403 ( .A(p_input[147]), .B(p_input[10147]), .Z(n18936) );
  AND U28404 ( .A(p_input[30147]), .B(p_input[20147]), .Z(n18935) );
  AND U28405 ( .A(n18937), .B(n18938), .Z(o[1479]) );
  AND U28406 ( .A(p_input[1479]), .B(p_input[11479]), .Z(n18938) );
  AND U28407 ( .A(p_input[31479]), .B(p_input[21479]), .Z(n18937) );
  AND U28408 ( .A(n18939), .B(n18940), .Z(o[1478]) );
  AND U28409 ( .A(p_input[1478]), .B(p_input[11478]), .Z(n18940) );
  AND U28410 ( .A(p_input[31478]), .B(p_input[21478]), .Z(n18939) );
  AND U28411 ( .A(n18941), .B(n18942), .Z(o[1477]) );
  AND U28412 ( .A(p_input[1477]), .B(p_input[11477]), .Z(n18942) );
  AND U28413 ( .A(p_input[31477]), .B(p_input[21477]), .Z(n18941) );
  AND U28414 ( .A(n18943), .B(n18944), .Z(o[1476]) );
  AND U28415 ( .A(p_input[1476]), .B(p_input[11476]), .Z(n18944) );
  AND U28416 ( .A(p_input[31476]), .B(p_input[21476]), .Z(n18943) );
  AND U28417 ( .A(n18945), .B(n18946), .Z(o[1475]) );
  AND U28418 ( .A(p_input[1475]), .B(p_input[11475]), .Z(n18946) );
  AND U28419 ( .A(p_input[31475]), .B(p_input[21475]), .Z(n18945) );
  AND U28420 ( .A(n18947), .B(n18948), .Z(o[1474]) );
  AND U28421 ( .A(p_input[1474]), .B(p_input[11474]), .Z(n18948) );
  AND U28422 ( .A(p_input[31474]), .B(p_input[21474]), .Z(n18947) );
  AND U28423 ( .A(n18949), .B(n18950), .Z(o[1473]) );
  AND U28424 ( .A(p_input[1473]), .B(p_input[11473]), .Z(n18950) );
  AND U28425 ( .A(p_input[31473]), .B(p_input[21473]), .Z(n18949) );
  AND U28426 ( .A(n18951), .B(n18952), .Z(o[1472]) );
  AND U28427 ( .A(p_input[1472]), .B(p_input[11472]), .Z(n18952) );
  AND U28428 ( .A(p_input[31472]), .B(p_input[21472]), .Z(n18951) );
  AND U28429 ( .A(n18953), .B(n18954), .Z(o[1471]) );
  AND U28430 ( .A(p_input[1471]), .B(p_input[11471]), .Z(n18954) );
  AND U28431 ( .A(p_input[31471]), .B(p_input[21471]), .Z(n18953) );
  AND U28432 ( .A(n18955), .B(n18956), .Z(o[1470]) );
  AND U28433 ( .A(p_input[1470]), .B(p_input[11470]), .Z(n18956) );
  AND U28434 ( .A(p_input[31470]), .B(p_input[21470]), .Z(n18955) );
  AND U28435 ( .A(n18957), .B(n18958), .Z(o[146]) );
  AND U28436 ( .A(p_input[146]), .B(p_input[10146]), .Z(n18958) );
  AND U28437 ( .A(p_input[30146]), .B(p_input[20146]), .Z(n18957) );
  AND U28438 ( .A(n18959), .B(n18960), .Z(o[1469]) );
  AND U28439 ( .A(p_input[1469]), .B(p_input[11469]), .Z(n18960) );
  AND U28440 ( .A(p_input[31469]), .B(p_input[21469]), .Z(n18959) );
  AND U28441 ( .A(n18961), .B(n18962), .Z(o[1468]) );
  AND U28442 ( .A(p_input[1468]), .B(p_input[11468]), .Z(n18962) );
  AND U28443 ( .A(p_input[31468]), .B(p_input[21468]), .Z(n18961) );
  AND U28444 ( .A(n18963), .B(n18964), .Z(o[1467]) );
  AND U28445 ( .A(p_input[1467]), .B(p_input[11467]), .Z(n18964) );
  AND U28446 ( .A(p_input[31467]), .B(p_input[21467]), .Z(n18963) );
  AND U28447 ( .A(n18965), .B(n18966), .Z(o[1466]) );
  AND U28448 ( .A(p_input[1466]), .B(p_input[11466]), .Z(n18966) );
  AND U28449 ( .A(p_input[31466]), .B(p_input[21466]), .Z(n18965) );
  AND U28450 ( .A(n18967), .B(n18968), .Z(o[1465]) );
  AND U28451 ( .A(p_input[1465]), .B(p_input[11465]), .Z(n18968) );
  AND U28452 ( .A(p_input[31465]), .B(p_input[21465]), .Z(n18967) );
  AND U28453 ( .A(n18969), .B(n18970), .Z(o[1464]) );
  AND U28454 ( .A(p_input[1464]), .B(p_input[11464]), .Z(n18970) );
  AND U28455 ( .A(p_input[31464]), .B(p_input[21464]), .Z(n18969) );
  AND U28456 ( .A(n18971), .B(n18972), .Z(o[1463]) );
  AND U28457 ( .A(p_input[1463]), .B(p_input[11463]), .Z(n18972) );
  AND U28458 ( .A(p_input[31463]), .B(p_input[21463]), .Z(n18971) );
  AND U28459 ( .A(n18973), .B(n18974), .Z(o[1462]) );
  AND U28460 ( .A(p_input[1462]), .B(p_input[11462]), .Z(n18974) );
  AND U28461 ( .A(p_input[31462]), .B(p_input[21462]), .Z(n18973) );
  AND U28462 ( .A(n18975), .B(n18976), .Z(o[1461]) );
  AND U28463 ( .A(p_input[1461]), .B(p_input[11461]), .Z(n18976) );
  AND U28464 ( .A(p_input[31461]), .B(p_input[21461]), .Z(n18975) );
  AND U28465 ( .A(n18977), .B(n18978), .Z(o[1460]) );
  AND U28466 ( .A(p_input[1460]), .B(p_input[11460]), .Z(n18978) );
  AND U28467 ( .A(p_input[31460]), .B(p_input[21460]), .Z(n18977) );
  AND U28468 ( .A(n18979), .B(n18980), .Z(o[145]) );
  AND U28469 ( .A(p_input[145]), .B(p_input[10145]), .Z(n18980) );
  AND U28470 ( .A(p_input[30145]), .B(p_input[20145]), .Z(n18979) );
  AND U28471 ( .A(n18981), .B(n18982), .Z(o[1459]) );
  AND U28472 ( .A(p_input[1459]), .B(p_input[11459]), .Z(n18982) );
  AND U28473 ( .A(p_input[31459]), .B(p_input[21459]), .Z(n18981) );
  AND U28474 ( .A(n18983), .B(n18984), .Z(o[1458]) );
  AND U28475 ( .A(p_input[1458]), .B(p_input[11458]), .Z(n18984) );
  AND U28476 ( .A(p_input[31458]), .B(p_input[21458]), .Z(n18983) );
  AND U28477 ( .A(n18985), .B(n18986), .Z(o[1457]) );
  AND U28478 ( .A(p_input[1457]), .B(p_input[11457]), .Z(n18986) );
  AND U28479 ( .A(p_input[31457]), .B(p_input[21457]), .Z(n18985) );
  AND U28480 ( .A(n18987), .B(n18988), .Z(o[1456]) );
  AND U28481 ( .A(p_input[1456]), .B(p_input[11456]), .Z(n18988) );
  AND U28482 ( .A(p_input[31456]), .B(p_input[21456]), .Z(n18987) );
  AND U28483 ( .A(n18989), .B(n18990), .Z(o[1455]) );
  AND U28484 ( .A(p_input[1455]), .B(p_input[11455]), .Z(n18990) );
  AND U28485 ( .A(p_input[31455]), .B(p_input[21455]), .Z(n18989) );
  AND U28486 ( .A(n18991), .B(n18992), .Z(o[1454]) );
  AND U28487 ( .A(p_input[1454]), .B(p_input[11454]), .Z(n18992) );
  AND U28488 ( .A(p_input[31454]), .B(p_input[21454]), .Z(n18991) );
  AND U28489 ( .A(n18993), .B(n18994), .Z(o[1453]) );
  AND U28490 ( .A(p_input[1453]), .B(p_input[11453]), .Z(n18994) );
  AND U28491 ( .A(p_input[31453]), .B(p_input[21453]), .Z(n18993) );
  AND U28492 ( .A(n18995), .B(n18996), .Z(o[1452]) );
  AND U28493 ( .A(p_input[1452]), .B(p_input[11452]), .Z(n18996) );
  AND U28494 ( .A(p_input[31452]), .B(p_input[21452]), .Z(n18995) );
  AND U28495 ( .A(n18997), .B(n18998), .Z(o[1451]) );
  AND U28496 ( .A(p_input[1451]), .B(p_input[11451]), .Z(n18998) );
  AND U28497 ( .A(p_input[31451]), .B(p_input[21451]), .Z(n18997) );
  AND U28498 ( .A(n18999), .B(n19000), .Z(o[1450]) );
  AND U28499 ( .A(p_input[1450]), .B(p_input[11450]), .Z(n19000) );
  AND U28500 ( .A(p_input[31450]), .B(p_input[21450]), .Z(n18999) );
  AND U28501 ( .A(n19001), .B(n19002), .Z(o[144]) );
  AND U28502 ( .A(p_input[144]), .B(p_input[10144]), .Z(n19002) );
  AND U28503 ( .A(p_input[30144]), .B(p_input[20144]), .Z(n19001) );
  AND U28504 ( .A(n19003), .B(n19004), .Z(o[1449]) );
  AND U28505 ( .A(p_input[1449]), .B(p_input[11449]), .Z(n19004) );
  AND U28506 ( .A(p_input[31449]), .B(p_input[21449]), .Z(n19003) );
  AND U28507 ( .A(n19005), .B(n19006), .Z(o[1448]) );
  AND U28508 ( .A(p_input[1448]), .B(p_input[11448]), .Z(n19006) );
  AND U28509 ( .A(p_input[31448]), .B(p_input[21448]), .Z(n19005) );
  AND U28510 ( .A(n19007), .B(n19008), .Z(o[1447]) );
  AND U28511 ( .A(p_input[1447]), .B(p_input[11447]), .Z(n19008) );
  AND U28512 ( .A(p_input[31447]), .B(p_input[21447]), .Z(n19007) );
  AND U28513 ( .A(n19009), .B(n19010), .Z(o[1446]) );
  AND U28514 ( .A(p_input[1446]), .B(p_input[11446]), .Z(n19010) );
  AND U28515 ( .A(p_input[31446]), .B(p_input[21446]), .Z(n19009) );
  AND U28516 ( .A(n19011), .B(n19012), .Z(o[1445]) );
  AND U28517 ( .A(p_input[1445]), .B(p_input[11445]), .Z(n19012) );
  AND U28518 ( .A(p_input[31445]), .B(p_input[21445]), .Z(n19011) );
  AND U28519 ( .A(n19013), .B(n19014), .Z(o[1444]) );
  AND U28520 ( .A(p_input[1444]), .B(p_input[11444]), .Z(n19014) );
  AND U28521 ( .A(p_input[31444]), .B(p_input[21444]), .Z(n19013) );
  AND U28522 ( .A(n19015), .B(n19016), .Z(o[1443]) );
  AND U28523 ( .A(p_input[1443]), .B(p_input[11443]), .Z(n19016) );
  AND U28524 ( .A(p_input[31443]), .B(p_input[21443]), .Z(n19015) );
  AND U28525 ( .A(n19017), .B(n19018), .Z(o[1442]) );
  AND U28526 ( .A(p_input[1442]), .B(p_input[11442]), .Z(n19018) );
  AND U28527 ( .A(p_input[31442]), .B(p_input[21442]), .Z(n19017) );
  AND U28528 ( .A(n19019), .B(n19020), .Z(o[1441]) );
  AND U28529 ( .A(p_input[1441]), .B(p_input[11441]), .Z(n19020) );
  AND U28530 ( .A(p_input[31441]), .B(p_input[21441]), .Z(n19019) );
  AND U28531 ( .A(n19021), .B(n19022), .Z(o[1440]) );
  AND U28532 ( .A(p_input[1440]), .B(p_input[11440]), .Z(n19022) );
  AND U28533 ( .A(p_input[31440]), .B(p_input[21440]), .Z(n19021) );
  AND U28534 ( .A(n19023), .B(n19024), .Z(o[143]) );
  AND U28535 ( .A(p_input[143]), .B(p_input[10143]), .Z(n19024) );
  AND U28536 ( .A(p_input[30143]), .B(p_input[20143]), .Z(n19023) );
  AND U28537 ( .A(n19025), .B(n19026), .Z(o[1439]) );
  AND U28538 ( .A(p_input[1439]), .B(p_input[11439]), .Z(n19026) );
  AND U28539 ( .A(p_input[31439]), .B(p_input[21439]), .Z(n19025) );
  AND U28540 ( .A(n19027), .B(n19028), .Z(o[1438]) );
  AND U28541 ( .A(p_input[1438]), .B(p_input[11438]), .Z(n19028) );
  AND U28542 ( .A(p_input[31438]), .B(p_input[21438]), .Z(n19027) );
  AND U28543 ( .A(n19029), .B(n19030), .Z(o[1437]) );
  AND U28544 ( .A(p_input[1437]), .B(p_input[11437]), .Z(n19030) );
  AND U28545 ( .A(p_input[31437]), .B(p_input[21437]), .Z(n19029) );
  AND U28546 ( .A(n19031), .B(n19032), .Z(o[1436]) );
  AND U28547 ( .A(p_input[1436]), .B(p_input[11436]), .Z(n19032) );
  AND U28548 ( .A(p_input[31436]), .B(p_input[21436]), .Z(n19031) );
  AND U28549 ( .A(n19033), .B(n19034), .Z(o[1435]) );
  AND U28550 ( .A(p_input[1435]), .B(p_input[11435]), .Z(n19034) );
  AND U28551 ( .A(p_input[31435]), .B(p_input[21435]), .Z(n19033) );
  AND U28552 ( .A(n19035), .B(n19036), .Z(o[1434]) );
  AND U28553 ( .A(p_input[1434]), .B(p_input[11434]), .Z(n19036) );
  AND U28554 ( .A(p_input[31434]), .B(p_input[21434]), .Z(n19035) );
  AND U28555 ( .A(n19037), .B(n19038), .Z(o[1433]) );
  AND U28556 ( .A(p_input[1433]), .B(p_input[11433]), .Z(n19038) );
  AND U28557 ( .A(p_input[31433]), .B(p_input[21433]), .Z(n19037) );
  AND U28558 ( .A(n19039), .B(n19040), .Z(o[1432]) );
  AND U28559 ( .A(p_input[1432]), .B(p_input[11432]), .Z(n19040) );
  AND U28560 ( .A(p_input[31432]), .B(p_input[21432]), .Z(n19039) );
  AND U28561 ( .A(n19041), .B(n19042), .Z(o[1431]) );
  AND U28562 ( .A(p_input[1431]), .B(p_input[11431]), .Z(n19042) );
  AND U28563 ( .A(p_input[31431]), .B(p_input[21431]), .Z(n19041) );
  AND U28564 ( .A(n19043), .B(n19044), .Z(o[1430]) );
  AND U28565 ( .A(p_input[1430]), .B(p_input[11430]), .Z(n19044) );
  AND U28566 ( .A(p_input[31430]), .B(p_input[21430]), .Z(n19043) );
  AND U28567 ( .A(n19045), .B(n19046), .Z(o[142]) );
  AND U28568 ( .A(p_input[142]), .B(p_input[10142]), .Z(n19046) );
  AND U28569 ( .A(p_input[30142]), .B(p_input[20142]), .Z(n19045) );
  AND U28570 ( .A(n19047), .B(n19048), .Z(o[1429]) );
  AND U28571 ( .A(p_input[1429]), .B(p_input[11429]), .Z(n19048) );
  AND U28572 ( .A(p_input[31429]), .B(p_input[21429]), .Z(n19047) );
  AND U28573 ( .A(n19049), .B(n19050), .Z(o[1428]) );
  AND U28574 ( .A(p_input[1428]), .B(p_input[11428]), .Z(n19050) );
  AND U28575 ( .A(p_input[31428]), .B(p_input[21428]), .Z(n19049) );
  AND U28576 ( .A(n19051), .B(n19052), .Z(o[1427]) );
  AND U28577 ( .A(p_input[1427]), .B(p_input[11427]), .Z(n19052) );
  AND U28578 ( .A(p_input[31427]), .B(p_input[21427]), .Z(n19051) );
  AND U28579 ( .A(n19053), .B(n19054), .Z(o[1426]) );
  AND U28580 ( .A(p_input[1426]), .B(p_input[11426]), .Z(n19054) );
  AND U28581 ( .A(p_input[31426]), .B(p_input[21426]), .Z(n19053) );
  AND U28582 ( .A(n19055), .B(n19056), .Z(o[1425]) );
  AND U28583 ( .A(p_input[1425]), .B(p_input[11425]), .Z(n19056) );
  AND U28584 ( .A(p_input[31425]), .B(p_input[21425]), .Z(n19055) );
  AND U28585 ( .A(n19057), .B(n19058), .Z(o[1424]) );
  AND U28586 ( .A(p_input[1424]), .B(p_input[11424]), .Z(n19058) );
  AND U28587 ( .A(p_input[31424]), .B(p_input[21424]), .Z(n19057) );
  AND U28588 ( .A(n19059), .B(n19060), .Z(o[1423]) );
  AND U28589 ( .A(p_input[1423]), .B(p_input[11423]), .Z(n19060) );
  AND U28590 ( .A(p_input[31423]), .B(p_input[21423]), .Z(n19059) );
  AND U28591 ( .A(n19061), .B(n19062), .Z(o[1422]) );
  AND U28592 ( .A(p_input[1422]), .B(p_input[11422]), .Z(n19062) );
  AND U28593 ( .A(p_input[31422]), .B(p_input[21422]), .Z(n19061) );
  AND U28594 ( .A(n19063), .B(n19064), .Z(o[1421]) );
  AND U28595 ( .A(p_input[1421]), .B(p_input[11421]), .Z(n19064) );
  AND U28596 ( .A(p_input[31421]), .B(p_input[21421]), .Z(n19063) );
  AND U28597 ( .A(n19065), .B(n19066), .Z(o[1420]) );
  AND U28598 ( .A(p_input[1420]), .B(p_input[11420]), .Z(n19066) );
  AND U28599 ( .A(p_input[31420]), .B(p_input[21420]), .Z(n19065) );
  AND U28600 ( .A(n19067), .B(n19068), .Z(o[141]) );
  AND U28601 ( .A(p_input[141]), .B(p_input[10141]), .Z(n19068) );
  AND U28602 ( .A(p_input[30141]), .B(p_input[20141]), .Z(n19067) );
  AND U28603 ( .A(n19069), .B(n19070), .Z(o[1419]) );
  AND U28604 ( .A(p_input[1419]), .B(p_input[11419]), .Z(n19070) );
  AND U28605 ( .A(p_input[31419]), .B(p_input[21419]), .Z(n19069) );
  AND U28606 ( .A(n19071), .B(n19072), .Z(o[1418]) );
  AND U28607 ( .A(p_input[1418]), .B(p_input[11418]), .Z(n19072) );
  AND U28608 ( .A(p_input[31418]), .B(p_input[21418]), .Z(n19071) );
  AND U28609 ( .A(n19073), .B(n19074), .Z(o[1417]) );
  AND U28610 ( .A(p_input[1417]), .B(p_input[11417]), .Z(n19074) );
  AND U28611 ( .A(p_input[31417]), .B(p_input[21417]), .Z(n19073) );
  AND U28612 ( .A(n19075), .B(n19076), .Z(o[1416]) );
  AND U28613 ( .A(p_input[1416]), .B(p_input[11416]), .Z(n19076) );
  AND U28614 ( .A(p_input[31416]), .B(p_input[21416]), .Z(n19075) );
  AND U28615 ( .A(n19077), .B(n19078), .Z(o[1415]) );
  AND U28616 ( .A(p_input[1415]), .B(p_input[11415]), .Z(n19078) );
  AND U28617 ( .A(p_input[31415]), .B(p_input[21415]), .Z(n19077) );
  AND U28618 ( .A(n19079), .B(n19080), .Z(o[1414]) );
  AND U28619 ( .A(p_input[1414]), .B(p_input[11414]), .Z(n19080) );
  AND U28620 ( .A(p_input[31414]), .B(p_input[21414]), .Z(n19079) );
  AND U28621 ( .A(n19081), .B(n19082), .Z(o[1413]) );
  AND U28622 ( .A(p_input[1413]), .B(p_input[11413]), .Z(n19082) );
  AND U28623 ( .A(p_input[31413]), .B(p_input[21413]), .Z(n19081) );
  AND U28624 ( .A(n19083), .B(n19084), .Z(o[1412]) );
  AND U28625 ( .A(p_input[1412]), .B(p_input[11412]), .Z(n19084) );
  AND U28626 ( .A(p_input[31412]), .B(p_input[21412]), .Z(n19083) );
  AND U28627 ( .A(n19085), .B(n19086), .Z(o[1411]) );
  AND U28628 ( .A(p_input[1411]), .B(p_input[11411]), .Z(n19086) );
  AND U28629 ( .A(p_input[31411]), .B(p_input[21411]), .Z(n19085) );
  AND U28630 ( .A(n19087), .B(n19088), .Z(o[1410]) );
  AND U28631 ( .A(p_input[1410]), .B(p_input[11410]), .Z(n19088) );
  AND U28632 ( .A(p_input[31410]), .B(p_input[21410]), .Z(n19087) );
  AND U28633 ( .A(n19089), .B(n19090), .Z(o[140]) );
  AND U28634 ( .A(p_input[140]), .B(p_input[10140]), .Z(n19090) );
  AND U28635 ( .A(p_input[30140]), .B(p_input[20140]), .Z(n19089) );
  AND U28636 ( .A(n19091), .B(n19092), .Z(o[1409]) );
  AND U28637 ( .A(p_input[1409]), .B(p_input[11409]), .Z(n19092) );
  AND U28638 ( .A(p_input[31409]), .B(p_input[21409]), .Z(n19091) );
  AND U28639 ( .A(n19093), .B(n19094), .Z(o[1408]) );
  AND U28640 ( .A(p_input[1408]), .B(p_input[11408]), .Z(n19094) );
  AND U28641 ( .A(p_input[31408]), .B(p_input[21408]), .Z(n19093) );
  AND U28642 ( .A(n19095), .B(n19096), .Z(o[1407]) );
  AND U28643 ( .A(p_input[1407]), .B(p_input[11407]), .Z(n19096) );
  AND U28644 ( .A(p_input[31407]), .B(p_input[21407]), .Z(n19095) );
  AND U28645 ( .A(n19097), .B(n19098), .Z(o[1406]) );
  AND U28646 ( .A(p_input[1406]), .B(p_input[11406]), .Z(n19098) );
  AND U28647 ( .A(p_input[31406]), .B(p_input[21406]), .Z(n19097) );
  AND U28648 ( .A(n19099), .B(n19100), .Z(o[1405]) );
  AND U28649 ( .A(p_input[1405]), .B(p_input[11405]), .Z(n19100) );
  AND U28650 ( .A(p_input[31405]), .B(p_input[21405]), .Z(n19099) );
  AND U28651 ( .A(n19101), .B(n19102), .Z(o[1404]) );
  AND U28652 ( .A(p_input[1404]), .B(p_input[11404]), .Z(n19102) );
  AND U28653 ( .A(p_input[31404]), .B(p_input[21404]), .Z(n19101) );
  AND U28654 ( .A(n19103), .B(n19104), .Z(o[1403]) );
  AND U28655 ( .A(p_input[1403]), .B(p_input[11403]), .Z(n19104) );
  AND U28656 ( .A(p_input[31403]), .B(p_input[21403]), .Z(n19103) );
  AND U28657 ( .A(n19105), .B(n19106), .Z(o[1402]) );
  AND U28658 ( .A(p_input[1402]), .B(p_input[11402]), .Z(n19106) );
  AND U28659 ( .A(p_input[31402]), .B(p_input[21402]), .Z(n19105) );
  AND U28660 ( .A(n19107), .B(n19108), .Z(o[1401]) );
  AND U28661 ( .A(p_input[1401]), .B(p_input[11401]), .Z(n19108) );
  AND U28662 ( .A(p_input[31401]), .B(p_input[21401]), .Z(n19107) );
  AND U28663 ( .A(n19109), .B(n19110), .Z(o[1400]) );
  AND U28664 ( .A(p_input[1400]), .B(p_input[11400]), .Z(n19110) );
  AND U28665 ( .A(p_input[31400]), .B(p_input[21400]), .Z(n19109) );
  AND U28666 ( .A(n19111), .B(n19112), .Z(o[13]) );
  AND U28667 ( .A(p_input[13]), .B(p_input[10013]), .Z(n19112) );
  AND U28668 ( .A(p_input[30013]), .B(p_input[20013]), .Z(n19111) );
  AND U28669 ( .A(n19113), .B(n19114), .Z(o[139]) );
  AND U28670 ( .A(p_input[139]), .B(p_input[10139]), .Z(n19114) );
  AND U28671 ( .A(p_input[30139]), .B(p_input[20139]), .Z(n19113) );
  AND U28672 ( .A(n19115), .B(n19116), .Z(o[1399]) );
  AND U28673 ( .A(p_input[1399]), .B(p_input[11399]), .Z(n19116) );
  AND U28674 ( .A(p_input[31399]), .B(p_input[21399]), .Z(n19115) );
  AND U28675 ( .A(n19117), .B(n19118), .Z(o[1398]) );
  AND U28676 ( .A(p_input[1398]), .B(p_input[11398]), .Z(n19118) );
  AND U28677 ( .A(p_input[31398]), .B(p_input[21398]), .Z(n19117) );
  AND U28678 ( .A(n19119), .B(n19120), .Z(o[1397]) );
  AND U28679 ( .A(p_input[1397]), .B(p_input[11397]), .Z(n19120) );
  AND U28680 ( .A(p_input[31397]), .B(p_input[21397]), .Z(n19119) );
  AND U28681 ( .A(n19121), .B(n19122), .Z(o[1396]) );
  AND U28682 ( .A(p_input[1396]), .B(p_input[11396]), .Z(n19122) );
  AND U28683 ( .A(p_input[31396]), .B(p_input[21396]), .Z(n19121) );
  AND U28684 ( .A(n19123), .B(n19124), .Z(o[1395]) );
  AND U28685 ( .A(p_input[1395]), .B(p_input[11395]), .Z(n19124) );
  AND U28686 ( .A(p_input[31395]), .B(p_input[21395]), .Z(n19123) );
  AND U28687 ( .A(n19125), .B(n19126), .Z(o[1394]) );
  AND U28688 ( .A(p_input[1394]), .B(p_input[11394]), .Z(n19126) );
  AND U28689 ( .A(p_input[31394]), .B(p_input[21394]), .Z(n19125) );
  AND U28690 ( .A(n19127), .B(n19128), .Z(o[1393]) );
  AND U28691 ( .A(p_input[1393]), .B(p_input[11393]), .Z(n19128) );
  AND U28692 ( .A(p_input[31393]), .B(p_input[21393]), .Z(n19127) );
  AND U28693 ( .A(n19129), .B(n19130), .Z(o[1392]) );
  AND U28694 ( .A(p_input[1392]), .B(p_input[11392]), .Z(n19130) );
  AND U28695 ( .A(p_input[31392]), .B(p_input[21392]), .Z(n19129) );
  AND U28696 ( .A(n19131), .B(n19132), .Z(o[1391]) );
  AND U28697 ( .A(p_input[1391]), .B(p_input[11391]), .Z(n19132) );
  AND U28698 ( .A(p_input[31391]), .B(p_input[21391]), .Z(n19131) );
  AND U28699 ( .A(n19133), .B(n19134), .Z(o[1390]) );
  AND U28700 ( .A(p_input[1390]), .B(p_input[11390]), .Z(n19134) );
  AND U28701 ( .A(p_input[31390]), .B(p_input[21390]), .Z(n19133) );
  AND U28702 ( .A(n19135), .B(n19136), .Z(o[138]) );
  AND U28703 ( .A(p_input[138]), .B(p_input[10138]), .Z(n19136) );
  AND U28704 ( .A(p_input[30138]), .B(p_input[20138]), .Z(n19135) );
  AND U28705 ( .A(n19137), .B(n19138), .Z(o[1389]) );
  AND U28706 ( .A(p_input[1389]), .B(p_input[11389]), .Z(n19138) );
  AND U28707 ( .A(p_input[31389]), .B(p_input[21389]), .Z(n19137) );
  AND U28708 ( .A(n19139), .B(n19140), .Z(o[1388]) );
  AND U28709 ( .A(p_input[1388]), .B(p_input[11388]), .Z(n19140) );
  AND U28710 ( .A(p_input[31388]), .B(p_input[21388]), .Z(n19139) );
  AND U28711 ( .A(n19141), .B(n19142), .Z(o[1387]) );
  AND U28712 ( .A(p_input[1387]), .B(p_input[11387]), .Z(n19142) );
  AND U28713 ( .A(p_input[31387]), .B(p_input[21387]), .Z(n19141) );
  AND U28714 ( .A(n19143), .B(n19144), .Z(o[1386]) );
  AND U28715 ( .A(p_input[1386]), .B(p_input[11386]), .Z(n19144) );
  AND U28716 ( .A(p_input[31386]), .B(p_input[21386]), .Z(n19143) );
  AND U28717 ( .A(n19145), .B(n19146), .Z(o[1385]) );
  AND U28718 ( .A(p_input[1385]), .B(p_input[11385]), .Z(n19146) );
  AND U28719 ( .A(p_input[31385]), .B(p_input[21385]), .Z(n19145) );
  AND U28720 ( .A(n19147), .B(n19148), .Z(o[1384]) );
  AND U28721 ( .A(p_input[1384]), .B(p_input[11384]), .Z(n19148) );
  AND U28722 ( .A(p_input[31384]), .B(p_input[21384]), .Z(n19147) );
  AND U28723 ( .A(n19149), .B(n19150), .Z(o[1383]) );
  AND U28724 ( .A(p_input[1383]), .B(p_input[11383]), .Z(n19150) );
  AND U28725 ( .A(p_input[31383]), .B(p_input[21383]), .Z(n19149) );
  AND U28726 ( .A(n19151), .B(n19152), .Z(o[1382]) );
  AND U28727 ( .A(p_input[1382]), .B(p_input[11382]), .Z(n19152) );
  AND U28728 ( .A(p_input[31382]), .B(p_input[21382]), .Z(n19151) );
  AND U28729 ( .A(n19153), .B(n19154), .Z(o[1381]) );
  AND U28730 ( .A(p_input[1381]), .B(p_input[11381]), .Z(n19154) );
  AND U28731 ( .A(p_input[31381]), .B(p_input[21381]), .Z(n19153) );
  AND U28732 ( .A(n19155), .B(n19156), .Z(o[1380]) );
  AND U28733 ( .A(p_input[1380]), .B(p_input[11380]), .Z(n19156) );
  AND U28734 ( .A(p_input[31380]), .B(p_input[21380]), .Z(n19155) );
  AND U28735 ( .A(n19157), .B(n19158), .Z(o[137]) );
  AND U28736 ( .A(p_input[137]), .B(p_input[10137]), .Z(n19158) );
  AND U28737 ( .A(p_input[30137]), .B(p_input[20137]), .Z(n19157) );
  AND U28738 ( .A(n19159), .B(n19160), .Z(o[1379]) );
  AND U28739 ( .A(p_input[1379]), .B(p_input[11379]), .Z(n19160) );
  AND U28740 ( .A(p_input[31379]), .B(p_input[21379]), .Z(n19159) );
  AND U28741 ( .A(n19161), .B(n19162), .Z(o[1378]) );
  AND U28742 ( .A(p_input[1378]), .B(p_input[11378]), .Z(n19162) );
  AND U28743 ( .A(p_input[31378]), .B(p_input[21378]), .Z(n19161) );
  AND U28744 ( .A(n19163), .B(n19164), .Z(o[1377]) );
  AND U28745 ( .A(p_input[1377]), .B(p_input[11377]), .Z(n19164) );
  AND U28746 ( .A(p_input[31377]), .B(p_input[21377]), .Z(n19163) );
  AND U28747 ( .A(n19165), .B(n19166), .Z(o[1376]) );
  AND U28748 ( .A(p_input[1376]), .B(p_input[11376]), .Z(n19166) );
  AND U28749 ( .A(p_input[31376]), .B(p_input[21376]), .Z(n19165) );
  AND U28750 ( .A(n19167), .B(n19168), .Z(o[1375]) );
  AND U28751 ( .A(p_input[1375]), .B(p_input[11375]), .Z(n19168) );
  AND U28752 ( .A(p_input[31375]), .B(p_input[21375]), .Z(n19167) );
  AND U28753 ( .A(n19169), .B(n19170), .Z(o[1374]) );
  AND U28754 ( .A(p_input[1374]), .B(p_input[11374]), .Z(n19170) );
  AND U28755 ( .A(p_input[31374]), .B(p_input[21374]), .Z(n19169) );
  AND U28756 ( .A(n19171), .B(n19172), .Z(o[1373]) );
  AND U28757 ( .A(p_input[1373]), .B(p_input[11373]), .Z(n19172) );
  AND U28758 ( .A(p_input[31373]), .B(p_input[21373]), .Z(n19171) );
  AND U28759 ( .A(n19173), .B(n19174), .Z(o[1372]) );
  AND U28760 ( .A(p_input[1372]), .B(p_input[11372]), .Z(n19174) );
  AND U28761 ( .A(p_input[31372]), .B(p_input[21372]), .Z(n19173) );
  AND U28762 ( .A(n19175), .B(n19176), .Z(o[1371]) );
  AND U28763 ( .A(p_input[1371]), .B(p_input[11371]), .Z(n19176) );
  AND U28764 ( .A(p_input[31371]), .B(p_input[21371]), .Z(n19175) );
  AND U28765 ( .A(n19177), .B(n19178), .Z(o[1370]) );
  AND U28766 ( .A(p_input[1370]), .B(p_input[11370]), .Z(n19178) );
  AND U28767 ( .A(p_input[31370]), .B(p_input[21370]), .Z(n19177) );
  AND U28768 ( .A(n19179), .B(n19180), .Z(o[136]) );
  AND U28769 ( .A(p_input[136]), .B(p_input[10136]), .Z(n19180) );
  AND U28770 ( .A(p_input[30136]), .B(p_input[20136]), .Z(n19179) );
  AND U28771 ( .A(n19181), .B(n19182), .Z(o[1369]) );
  AND U28772 ( .A(p_input[1369]), .B(p_input[11369]), .Z(n19182) );
  AND U28773 ( .A(p_input[31369]), .B(p_input[21369]), .Z(n19181) );
  AND U28774 ( .A(n19183), .B(n19184), .Z(o[1368]) );
  AND U28775 ( .A(p_input[1368]), .B(p_input[11368]), .Z(n19184) );
  AND U28776 ( .A(p_input[31368]), .B(p_input[21368]), .Z(n19183) );
  AND U28777 ( .A(n19185), .B(n19186), .Z(o[1367]) );
  AND U28778 ( .A(p_input[1367]), .B(p_input[11367]), .Z(n19186) );
  AND U28779 ( .A(p_input[31367]), .B(p_input[21367]), .Z(n19185) );
  AND U28780 ( .A(n19187), .B(n19188), .Z(o[1366]) );
  AND U28781 ( .A(p_input[1366]), .B(p_input[11366]), .Z(n19188) );
  AND U28782 ( .A(p_input[31366]), .B(p_input[21366]), .Z(n19187) );
  AND U28783 ( .A(n19189), .B(n19190), .Z(o[1365]) );
  AND U28784 ( .A(p_input[1365]), .B(p_input[11365]), .Z(n19190) );
  AND U28785 ( .A(p_input[31365]), .B(p_input[21365]), .Z(n19189) );
  AND U28786 ( .A(n19191), .B(n19192), .Z(o[1364]) );
  AND U28787 ( .A(p_input[1364]), .B(p_input[11364]), .Z(n19192) );
  AND U28788 ( .A(p_input[31364]), .B(p_input[21364]), .Z(n19191) );
  AND U28789 ( .A(n19193), .B(n19194), .Z(o[1363]) );
  AND U28790 ( .A(p_input[1363]), .B(p_input[11363]), .Z(n19194) );
  AND U28791 ( .A(p_input[31363]), .B(p_input[21363]), .Z(n19193) );
  AND U28792 ( .A(n19195), .B(n19196), .Z(o[1362]) );
  AND U28793 ( .A(p_input[1362]), .B(p_input[11362]), .Z(n19196) );
  AND U28794 ( .A(p_input[31362]), .B(p_input[21362]), .Z(n19195) );
  AND U28795 ( .A(n19197), .B(n19198), .Z(o[1361]) );
  AND U28796 ( .A(p_input[1361]), .B(p_input[11361]), .Z(n19198) );
  AND U28797 ( .A(p_input[31361]), .B(p_input[21361]), .Z(n19197) );
  AND U28798 ( .A(n19199), .B(n19200), .Z(o[1360]) );
  AND U28799 ( .A(p_input[1360]), .B(p_input[11360]), .Z(n19200) );
  AND U28800 ( .A(p_input[31360]), .B(p_input[21360]), .Z(n19199) );
  AND U28801 ( .A(n19201), .B(n19202), .Z(o[135]) );
  AND U28802 ( .A(p_input[135]), .B(p_input[10135]), .Z(n19202) );
  AND U28803 ( .A(p_input[30135]), .B(p_input[20135]), .Z(n19201) );
  AND U28804 ( .A(n19203), .B(n19204), .Z(o[1359]) );
  AND U28805 ( .A(p_input[1359]), .B(p_input[11359]), .Z(n19204) );
  AND U28806 ( .A(p_input[31359]), .B(p_input[21359]), .Z(n19203) );
  AND U28807 ( .A(n19205), .B(n19206), .Z(o[1358]) );
  AND U28808 ( .A(p_input[1358]), .B(p_input[11358]), .Z(n19206) );
  AND U28809 ( .A(p_input[31358]), .B(p_input[21358]), .Z(n19205) );
  AND U28810 ( .A(n19207), .B(n19208), .Z(o[1357]) );
  AND U28811 ( .A(p_input[1357]), .B(p_input[11357]), .Z(n19208) );
  AND U28812 ( .A(p_input[31357]), .B(p_input[21357]), .Z(n19207) );
  AND U28813 ( .A(n19209), .B(n19210), .Z(o[1356]) );
  AND U28814 ( .A(p_input[1356]), .B(p_input[11356]), .Z(n19210) );
  AND U28815 ( .A(p_input[31356]), .B(p_input[21356]), .Z(n19209) );
  AND U28816 ( .A(n19211), .B(n19212), .Z(o[1355]) );
  AND U28817 ( .A(p_input[1355]), .B(p_input[11355]), .Z(n19212) );
  AND U28818 ( .A(p_input[31355]), .B(p_input[21355]), .Z(n19211) );
  AND U28819 ( .A(n19213), .B(n19214), .Z(o[1354]) );
  AND U28820 ( .A(p_input[1354]), .B(p_input[11354]), .Z(n19214) );
  AND U28821 ( .A(p_input[31354]), .B(p_input[21354]), .Z(n19213) );
  AND U28822 ( .A(n19215), .B(n19216), .Z(o[1353]) );
  AND U28823 ( .A(p_input[1353]), .B(p_input[11353]), .Z(n19216) );
  AND U28824 ( .A(p_input[31353]), .B(p_input[21353]), .Z(n19215) );
  AND U28825 ( .A(n19217), .B(n19218), .Z(o[1352]) );
  AND U28826 ( .A(p_input[1352]), .B(p_input[11352]), .Z(n19218) );
  AND U28827 ( .A(p_input[31352]), .B(p_input[21352]), .Z(n19217) );
  AND U28828 ( .A(n19219), .B(n19220), .Z(o[1351]) );
  AND U28829 ( .A(p_input[1351]), .B(p_input[11351]), .Z(n19220) );
  AND U28830 ( .A(p_input[31351]), .B(p_input[21351]), .Z(n19219) );
  AND U28831 ( .A(n19221), .B(n19222), .Z(o[1350]) );
  AND U28832 ( .A(p_input[1350]), .B(p_input[11350]), .Z(n19222) );
  AND U28833 ( .A(p_input[31350]), .B(p_input[21350]), .Z(n19221) );
  AND U28834 ( .A(n19223), .B(n19224), .Z(o[134]) );
  AND U28835 ( .A(p_input[134]), .B(p_input[10134]), .Z(n19224) );
  AND U28836 ( .A(p_input[30134]), .B(p_input[20134]), .Z(n19223) );
  AND U28837 ( .A(n19225), .B(n19226), .Z(o[1349]) );
  AND U28838 ( .A(p_input[1349]), .B(p_input[11349]), .Z(n19226) );
  AND U28839 ( .A(p_input[31349]), .B(p_input[21349]), .Z(n19225) );
  AND U28840 ( .A(n19227), .B(n19228), .Z(o[1348]) );
  AND U28841 ( .A(p_input[1348]), .B(p_input[11348]), .Z(n19228) );
  AND U28842 ( .A(p_input[31348]), .B(p_input[21348]), .Z(n19227) );
  AND U28843 ( .A(n19229), .B(n19230), .Z(o[1347]) );
  AND U28844 ( .A(p_input[1347]), .B(p_input[11347]), .Z(n19230) );
  AND U28845 ( .A(p_input[31347]), .B(p_input[21347]), .Z(n19229) );
  AND U28846 ( .A(n19231), .B(n19232), .Z(o[1346]) );
  AND U28847 ( .A(p_input[1346]), .B(p_input[11346]), .Z(n19232) );
  AND U28848 ( .A(p_input[31346]), .B(p_input[21346]), .Z(n19231) );
  AND U28849 ( .A(n19233), .B(n19234), .Z(o[1345]) );
  AND U28850 ( .A(p_input[1345]), .B(p_input[11345]), .Z(n19234) );
  AND U28851 ( .A(p_input[31345]), .B(p_input[21345]), .Z(n19233) );
  AND U28852 ( .A(n19235), .B(n19236), .Z(o[1344]) );
  AND U28853 ( .A(p_input[1344]), .B(p_input[11344]), .Z(n19236) );
  AND U28854 ( .A(p_input[31344]), .B(p_input[21344]), .Z(n19235) );
  AND U28855 ( .A(n19237), .B(n19238), .Z(o[1343]) );
  AND U28856 ( .A(p_input[1343]), .B(p_input[11343]), .Z(n19238) );
  AND U28857 ( .A(p_input[31343]), .B(p_input[21343]), .Z(n19237) );
  AND U28858 ( .A(n19239), .B(n19240), .Z(o[1342]) );
  AND U28859 ( .A(p_input[1342]), .B(p_input[11342]), .Z(n19240) );
  AND U28860 ( .A(p_input[31342]), .B(p_input[21342]), .Z(n19239) );
  AND U28861 ( .A(n19241), .B(n19242), .Z(o[1341]) );
  AND U28862 ( .A(p_input[1341]), .B(p_input[11341]), .Z(n19242) );
  AND U28863 ( .A(p_input[31341]), .B(p_input[21341]), .Z(n19241) );
  AND U28864 ( .A(n19243), .B(n19244), .Z(o[1340]) );
  AND U28865 ( .A(p_input[1340]), .B(p_input[11340]), .Z(n19244) );
  AND U28866 ( .A(p_input[31340]), .B(p_input[21340]), .Z(n19243) );
  AND U28867 ( .A(n19245), .B(n19246), .Z(o[133]) );
  AND U28868 ( .A(p_input[133]), .B(p_input[10133]), .Z(n19246) );
  AND U28869 ( .A(p_input[30133]), .B(p_input[20133]), .Z(n19245) );
  AND U28870 ( .A(n19247), .B(n19248), .Z(o[1339]) );
  AND U28871 ( .A(p_input[1339]), .B(p_input[11339]), .Z(n19248) );
  AND U28872 ( .A(p_input[31339]), .B(p_input[21339]), .Z(n19247) );
  AND U28873 ( .A(n19249), .B(n19250), .Z(o[1338]) );
  AND U28874 ( .A(p_input[1338]), .B(p_input[11338]), .Z(n19250) );
  AND U28875 ( .A(p_input[31338]), .B(p_input[21338]), .Z(n19249) );
  AND U28876 ( .A(n19251), .B(n19252), .Z(o[1337]) );
  AND U28877 ( .A(p_input[1337]), .B(p_input[11337]), .Z(n19252) );
  AND U28878 ( .A(p_input[31337]), .B(p_input[21337]), .Z(n19251) );
  AND U28879 ( .A(n19253), .B(n19254), .Z(o[1336]) );
  AND U28880 ( .A(p_input[1336]), .B(p_input[11336]), .Z(n19254) );
  AND U28881 ( .A(p_input[31336]), .B(p_input[21336]), .Z(n19253) );
  AND U28882 ( .A(n19255), .B(n19256), .Z(o[1335]) );
  AND U28883 ( .A(p_input[1335]), .B(p_input[11335]), .Z(n19256) );
  AND U28884 ( .A(p_input[31335]), .B(p_input[21335]), .Z(n19255) );
  AND U28885 ( .A(n19257), .B(n19258), .Z(o[1334]) );
  AND U28886 ( .A(p_input[1334]), .B(p_input[11334]), .Z(n19258) );
  AND U28887 ( .A(p_input[31334]), .B(p_input[21334]), .Z(n19257) );
  AND U28888 ( .A(n19259), .B(n19260), .Z(o[1333]) );
  AND U28889 ( .A(p_input[1333]), .B(p_input[11333]), .Z(n19260) );
  AND U28890 ( .A(p_input[31333]), .B(p_input[21333]), .Z(n19259) );
  AND U28891 ( .A(n19261), .B(n19262), .Z(o[1332]) );
  AND U28892 ( .A(p_input[1332]), .B(p_input[11332]), .Z(n19262) );
  AND U28893 ( .A(p_input[31332]), .B(p_input[21332]), .Z(n19261) );
  AND U28894 ( .A(n19263), .B(n19264), .Z(o[1331]) );
  AND U28895 ( .A(p_input[1331]), .B(p_input[11331]), .Z(n19264) );
  AND U28896 ( .A(p_input[31331]), .B(p_input[21331]), .Z(n19263) );
  AND U28897 ( .A(n19265), .B(n19266), .Z(o[1330]) );
  AND U28898 ( .A(p_input[1330]), .B(p_input[11330]), .Z(n19266) );
  AND U28899 ( .A(p_input[31330]), .B(p_input[21330]), .Z(n19265) );
  AND U28900 ( .A(n19267), .B(n19268), .Z(o[132]) );
  AND U28901 ( .A(p_input[132]), .B(p_input[10132]), .Z(n19268) );
  AND U28902 ( .A(p_input[30132]), .B(p_input[20132]), .Z(n19267) );
  AND U28903 ( .A(n19269), .B(n19270), .Z(o[1329]) );
  AND U28904 ( .A(p_input[1329]), .B(p_input[11329]), .Z(n19270) );
  AND U28905 ( .A(p_input[31329]), .B(p_input[21329]), .Z(n19269) );
  AND U28906 ( .A(n19271), .B(n19272), .Z(o[1328]) );
  AND U28907 ( .A(p_input[1328]), .B(p_input[11328]), .Z(n19272) );
  AND U28908 ( .A(p_input[31328]), .B(p_input[21328]), .Z(n19271) );
  AND U28909 ( .A(n19273), .B(n19274), .Z(o[1327]) );
  AND U28910 ( .A(p_input[1327]), .B(p_input[11327]), .Z(n19274) );
  AND U28911 ( .A(p_input[31327]), .B(p_input[21327]), .Z(n19273) );
  AND U28912 ( .A(n19275), .B(n19276), .Z(o[1326]) );
  AND U28913 ( .A(p_input[1326]), .B(p_input[11326]), .Z(n19276) );
  AND U28914 ( .A(p_input[31326]), .B(p_input[21326]), .Z(n19275) );
  AND U28915 ( .A(n19277), .B(n19278), .Z(o[1325]) );
  AND U28916 ( .A(p_input[1325]), .B(p_input[11325]), .Z(n19278) );
  AND U28917 ( .A(p_input[31325]), .B(p_input[21325]), .Z(n19277) );
  AND U28918 ( .A(n19279), .B(n19280), .Z(o[1324]) );
  AND U28919 ( .A(p_input[1324]), .B(p_input[11324]), .Z(n19280) );
  AND U28920 ( .A(p_input[31324]), .B(p_input[21324]), .Z(n19279) );
  AND U28921 ( .A(n19281), .B(n19282), .Z(o[1323]) );
  AND U28922 ( .A(p_input[1323]), .B(p_input[11323]), .Z(n19282) );
  AND U28923 ( .A(p_input[31323]), .B(p_input[21323]), .Z(n19281) );
  AND U28924 ( .A(n19283), .B(n19284), .Z(o[1322]) );
  AND U28925 ( .A(p_input[1322]), .B(p_input[11322]), .Z(n19284) );
  AND U28926 ( .A(p_input[31322]), .B(p_input[21322]), .Z(n19283) );
  AND U28927 ( .A(n19285), .B(n19286), .Z(o[1321]) );
  AND U28928 ( .A(p_input[1321]), .B(p_input[11321]), .Z(n19286) );
  AND U28929 ( .A(p_input[31321]), .B(p_input[21321]), .Z(n19285) );
  AND U28930 ( .A(n19287), .B(n19288), .Z(o[1320]) );
  AND U28931 ( .A(p_input[1320]), .B(p_input[11320]), .Z(n19288) );
  AND U28932 ( .A(p_input[31320]), .B(p_input[21320]), .Z(n19287) );
  AND U28933 ( .A(n19289), .B(n19290), .Z(o[131]) );
  AND U28934 ( .A(p_input[131]), .B(p_input[10131]), .Z(n19290) );
  AND U28935 ( .A(p_input[30131]), .B(p_input[20131]), .Z(n19289) );
  AND U28936 ( .A(n19291), .B(n19292), .Z(o[1319]) );
  AND U28937 ( .A(p_input[1319]), .B(p_input[11319]), .Z(n19292) );
  AND U28938 ( .A(p_input[31319]), .B(p_input[21319]), .Z(n19291) );
  AND U28939 ( .A(n19293), .B(n19294), .Z(o[1318]) );
  AND U28940 ( .A(p_input[1318]), .B(p_input[11318]), .Z(n19294) );
  AND U28941 ( .A(p_input[31318]), .B(p_input[21318]), .Z(n19293) );
  AND U28942 ( .A(n19295), .B(n19296), .Z(o[1317]) );
  AND U28943 ( .A(p_input[1317]), .B(p_input[11317]), .Z(n19296) );
  AND U28944 ( .A(p_input[31317]), .B(p_input[21317]), .Z(n19295) );
  AND U28945 ( .A(n19297), .B(n19298), .Z(o[1316]) );
  AND U28946 ( .A(p_input[1316]), .B(p_input[11316]), .Z(n19298) );
  AND U28947 ( .A(p_input[31316]), .B(p_input[21316]), .Z(n19297) );
  AND U28948 ( .A(n19299), .B(n19300), .Z(o[1315]) );
  AND U28949 ( .A(p_input[1315]), .B(p_input[11315]), .Z(n19300) );
  AND U28950 ( .A(p_input[31315]), .B(p_input[21315]), .Z(n19299) );
  AND U28951 ( .A(n19301), .B(n19302), .Z(o[1314]) );
  AND U28952 ( .A(p_input[1314]), .B(p_input[11314]), .Z(n19302) );
  AND U28953 ( .A(p_input[31314]), .B(p_input[21314]), .Z(n19301) );
  AND U28954 ( .A(n19303), .B(n19304), .Z(o[1313]) );
  AND U28955 ( .A(p_input[1313]), .B(p_input[11313]), .Z(n19304) );
  AND U28956 ( .A(p_input[31313]), .B(p_input[21313]), .Z(n19303) );
  AND U28957 ( .A(n19305), .B(n19306), .Z(o[1312]) );
  AND U28958 ( .A(p_input[1312]), .B(p_input[11312]), .Z(n19306) );
  AND U28959 ( .A(p_input[31312]), .B(p_input[21312]), .Z(n19305) );
  AND U28960 ( .A(n19307), .B(n19308), .Z(o[1311]) );
  AND U28961 ( .A(p_input[1311]), .B(p_input[11311]), .Z(n19308) );
  AND U28962 ( .A(p_input[31311]), .B(p_input[21311]), .Z(n19307) );
  AND U28963 ( .A(n19309), .B(n19310), .Z(o[1310]) );
  AND U28964 ( .A(p_input[1310]), .B(p_input[11310]), .Z(n19310) );
  AND U28965 ( .A(p_input[31310]), .B(p_input[21310]), .Z(n19309) );
  AND U28966 ( .A(n19311), .B(n19312), .Z(o[130]) );
  AND U28967 ( .A(p_input[130]), .B(p_input[10130]), .Z(n19312) );
  AND U28968 ( .A(p_input[30130]), .B(p_input[20130]), .Z(n19311) );
  AND U28969 ( .A(n19313), .B(n19314), .Z(o[1309]) );
  AND U28970 ( .A(p_input[1309]), .B(p_input[11309]), .Z(n19314) );
  AND U28971 ( .A(p_input[31309]), .B(p_input[21309]), .Z(n19313) );
  AND U28972 ( .A(n19315), .B(n19316), .Z(o[1308]) );
  AND U28973 ( .A(p_input[1308]), .B(p_input[11308]), .Z(n19316) );
  AND U28974 ( .A(p_input[31308]), .B(p_input[21308]), .Z(n19315) );
  AND U28975 ( .A(n19317), .B(n19318), .Z(o[1307]) );
  AND U28976 ( .A(p_input[1307]), .B(p_input[11307]), .Z(n19318) );
  AND U28977 ( .A(p_input[31307]), .B(p_input[21307]), .Z(n19317) );
  AND U28978 ( .A(n19319), .B(n19320), .Z(o[1306]) );
  AND U28979 ( .A(p_input[1306]), .B(p_input[11306]), .Z(n19320) );
  AND U28980 ( .A(p_input[31306]), .B(p_input[21306]), .Z(n19319) );
  AND U28981 ( .A(n19321), .B(n19322), .Z(o[1305]) );
  AND U28982 ( .A(p_input[1305]), .B(p_input[11305]), .Z(n19322) );
  AND U28983 ( .A(p_input[31305]), .B(p_input[21305]), .Z(n19321) );
  AND U28984 ( .A(n19323), .B(n19324), .Z(o[1304]) );
  AND U28985 ( .A(p_input[1304]), .B(p_input[11304]), .Z(n19324) );
  AND U28986 ( .A(p_input[31304]), .B(p_input[21304]), .Z(n19323) );
  AND U28987 ( .A(n19325), .B(n19326), .Z(o[1303]) );
  AND U28988 ( .A(p_input[1303]), .B(p_input[11303]), .Z(n19326) );
  AND U28989 ( .A(p_input[31303]), .B(p_input[21303]), .Z(n19325) );
  AND U28990 ( .A(n19327), .B(n19328), .Z(o[1302]) );
  AND U28991 ( .A(p_input[1302]), .B(p_input[11302]), .Z(n19328) );
  AND U28992 ( .A(p_input[31302]), .B(p_input[21302]), .Z(n19327) );
  AND U28993 ( .A(n19329), .B(n19330), .Z(o[1301]) );
  AND U28994 ( .A(p_input[1301]), .B(p_input[11301]), .Z(n19330) );
  AND U28995 ( .A(p_input[31301]), .B(p_input[21301]), .Z(n19329) );
  AND U28996 ( .A(n19331), .B(n19332), .Z(o[1300]) );
  AND U28997 ( .A(p_input[1300]), .B(p_input[11300]), .Z(n19332) );
  AND U28998 ( .A(p_input[31300]), .B(p_input[21300]), .Z(n19331) );
  AND U28999 ( .A(n19333), .B(n19334), .Z(o[12]) );
  AND U29000 ( .A(p_input[12]), .B(p_input[10012]), .Z(n19334) );
  AND U29001 ( .A(p_input[30012]), .B(p_input[20012]), .Z(n19333) );
  AND U29002 ( .A(n19335), .B(n19336), .Z(o[129]) );
  AND U29003 ( .A(p_input[129]), .B(p_input[10129]), .Z(n19336) );
  AND U29004 ( .A(p_input[30129]), .B(p_input[20129]), .Z(n19335) );
  AND U29005 ( .A(n19337), .B(n19338), .Z(o[1299]) );
  AND U29006 ( .A(p_input[1299]), .B(p_input[11299]), .Z(n19338) );
  AND U29007 ( .A(p_input[31299]), .B(p_input[21299]), .Z(n19337) );
  AND U29008 ( .A(n19339), .B(n19340), .Z(o[1298]) );
  AND U29009 ( .A(p_input[1298]), .B(p_input[11298]), .Z(n19340) );
  AND U29010 ( .A(p_input[31298]), .B(p_input[21298]), .Z(n19339) );
  AND U29011 ( .A(n19341), .B(n19342), .Z(o[1297]) );
  AND U29012 ( .A(p_input[1297]), .B(p_input[11297]), .Z(n19342) );
  AND U29013 ( .A(p_input[31297]), .B(p_input[21297]), .Z(n19341) );
  AND U29014 ( .A(n19343), .B(n19344), .Z(o[1296]) );
  AND U29015 ( .A(p_input[1296]), .B(p_input[11296]), .Z(n19344) );
  AND U29016 ( .A(p_input[31296]), .B(p_input[21296]), .Z(n19343) );
  AND U29017 ( .A(n19345), .B(n19346), .Z(o[1295]) );
  AND U29018 ( .A(p_input[1295]), .B(p_input[11295]), .Z(n19346) );
  AND U29019 ( .A(p_input[31295]), .B(p_input[21295]), .Z(n19345) );
  AND U29020 ( .A(n19347), .B(n19348), .Z(o[1294]) );
  AND U29021 ( .A(p_input[1294]), .B(p_input[11294]), .Z(n19348) );
  AND U29022 ( .A(p_input[31294]), .B(p_input[21294]), .Z(n19347) );
  AND U29023 ( .A(n19349), .B(n19350), .Z(o[1293]) );
  AND U29024 ( .A(p_input[1293]), .B(p_input[11293]), .Z(n19350) );
  AND U29025 ( .A(p_input[31293]), .B(p_input[21293]), .Z(n19349) );
  AND U29026 ( .A(n19351), .B(n19352), .Z(o[1292]) );
  AND U29027 ( .A(p_input[1292]), .B(p_input[11292]), .Z(n19352) );
  AND U29028 ( .A(p_input[31292]), .B(p_input[21292]), .Z(n19351) );
  AND U29029 ( .A(n19353), .B(n19354), .Z(o[1291]) );
  AND U29030 ( .A(p_input[1291]), .B(p_input[11291]), .Z(n19354) );
  AND U29031 ( .A(p_input[31291]), .B(p_input[21291]), .Z(n19353) );
  AND U29032 ( .A(n19355), .B(n19356), .Z(o[1290]) );
  AND U29033 ( .A(p_input[1290]), .B(p_input[11290]), .Z(n19356) );
  AND U29034 ( .A(p_input[31290]), .B(p_input[21290]), .Z(n19355) );
  AND U29035 ( .A(n19357), .B(n19358), .Z(o[128]) );
  AND U29036 ( .A(p_input[128]), .B(p_input[10128]), .Z(n19358) );
  AND U29037 ( .A(p_input[30128]), .B(p_input[20128]), .Z(n19357) );
  AND U29038 ( .A(n19359), .B(n19360), .Z(o[1289]) );
  AND U29039 ( .A(p_input[1289]), .B(p_input[11289]), .Z(n19360) );
  AND U29040 ( .A(p_input[31289]), .B(p_input[21289]), .Z(n19359) );
  AND U29041 ( .A(n19361), .B(n19362), .Z(o[1288]) );
  AND U29042 ( .A(p_input[1288]), .B(p_input[11288]), .Z(n19362) );
  AND U29043 ( .A(p_input[31288]), .B(p_input[21288]), .Z(n19361) );
  AND U29044 ( .A(n19363), .B(n19364), .Z(o[1287]) );
  AND U29045 ( .A(p_input[1287]), .B(p_input[11287]), .Z(n19364) );
  AND U29046 ( .A(p_input[31287]), .B(p_input[21287]), .Z(n19363) );
  AND U29047 ( .A(n19365), .B(n19366), .Z(o[1286]) );
  AND U29048 ( .A(p_input[1286]), .B(p_input[11286]), .Z(n19366) );
  AND U29049 ( .A(p_input[31286]), .B(p_input[21286]), .Z(n19365) );
  AND U29050 ( .A(n19367), .B(n19368), .Z(o[1285]) );
  AND U29051 ( .A(p_input[1285]), .B(p_input[11285]), .Z(n19368) );
  AND U29052 ( .A(p_input[31285]), .B(p_input[21285]), .Z(n19367) );
  AND U29053 ( .A(n19369), .B(n19370), .Z(o[1284]) );
  AND U29054 ( .A(p_input[1284]), .B(p_input[11284]), .Z(n19370) );
  AND U29055 ( .A(p_input[31284]), .B(p_input[21284]), .Z(n19369) );
  AND U29056 ( .A(n19371), .B(n19372), .Z(o[1283]) );
  AND U29057 ( .A(p_input[1283]), .B(p_input[11283]), .Z(n19372) );
  AND U29058 ( .A(p_input[31283]), .B(p_input[21283]), .Z(n19371) );
  AND U29059 ( .A(n19373), .B(n19374), .Z(o[1282]) );
  AND U29060 ( .A(p_input[1282]), .B(p_input[11282]), .Z(n19374) );
  AND U29061 ( .A(p_input[31282]), .B(p_input[21282]), .Z(n19373) );
  AND U29062 ( .A(n19375), .B(n19376), .Z(o[1281]) );
  AND U29063 ( .A(p_input[1281]), .B(p_input[11281]), .Z(n19376) );
  AND U29064 ( .A(p_input[31281]), .B(p_input[21281]), .Z(n19375) );
  AND U29065 ( .A(n19377), .B(n19378), .Z(o[1280]) );
  AND U29066 ( .A(p_input[1280]), .B(p_input[11280]), .Z(n19378) );
  AND U29067 ( .A(p_input[31280]), .B(p_input[21280]), .Z(n19377) );
  AND U29068 ( .A(n19379), .B(n19380), .Z(o[127]) );
  AND U29069 ( .A(p_input[127]), .B(p_input[10127]), .Z(n19380) );
  AND U29070 ( .A(p_input[30127]), .B(p_input[20127]), .Z(n19379) );
  AND U29071 ( .A(n19381), .B(n19382), .Z(o[1279]) );
  AND U29072 ( .A(p_input[1279]), .B(p_input[11279]), .Z(n19382) );
  AND U29073 ( .A(p_input[31279]), .B(p_input[21279]), .Z(n19381) );
  AND U29074 ( .A(n19383), .B(n19384), .Z(o[1278]) );
  AND U29075 ( .A(p_input[1278]), .B(p_input[11278]), .Z(n19384) );
  AND U29076 ( .A(p_input[31278]), .B(p_input[21278]), .Z(n19383) );
  AND U29077 ( .A(n19385), .B(n19386), .Z(o[1277]) );
  AND U29078 ( .A(p_input[1277]), .B(p_input[11277]), .Z(n19386) );
  AND U29079 ( .A(p_input[31277]), .B(p_input[21277]), .Z(n19385) );
  AND U29080 ( .A(n19387), .B(n19388), .Z(o[1276]) );
  AND U29081 ( .A(p_input[1276]), .B(p_input[11276]), .Z(n19388) );
  AND U29082 ( .A(p_input[31276]), .B(p_input[21276]), .Z(n19387) );
  AND U29083 ( .A(n19389), .B(n19390), .Z(o[1275]) );
  AND U29084 ( .A(p_input[1275]), .B(p_input[11275]), .Z(n19390) );
  AND U29085 ( .A(p_input[31275]), .B(p_input[21275]), .Z(n19389) );
  AND U29086 ( .A(n19391), .B(n19392), .Z(o[1274]) );
  AND U29087 ( .A(p_input[1274]), .B(p_input[11274]), .Z(n19392) );
  AND U29088 ( .A(p_input[31274]), .B(p_input[21274]), .Z(n19391) );
  AND U29089 ( .A(n19393), .B(n19394), .Z(o[1273]) );
  AND U29090 ( .A(p_input[1273]), .B(p_input[11273]), .Z(n19394) );
  AND U29091 ( .A(p_input[31273]), .B(p_input[21273]), .Z(n19393) );
  AND U29092 ( .A(n19395), .B(n19396), .Z(o[1272]) );
  AND U29093 ( .A(p_input[1272]), .B(p_input[11272]), .Z(n19396) );
  AND U29094 ( .A(p_input[31272]), .B(p_input[21272]), .Z(n19395) );
  AND U29095 ( .A(n19397), .B(n19398), .Z(o[1271]) );
  AND U29096 ( .A(p_input[1271]), .B(p_input[11271]), .Z(n19398) );
  AND U29097 ( .A(p_input[31271]), .B(p_input[21271]), .Z(n19397) );
  AND U29098 ( .A(n19399), .B(n19400), .Z(o[1270]) );
  AND U29099 ( .A(p_input[1270]), .B(p_input[11270]), .Z(n19400) );
  AND U29100 ( .A(p_input[31270]), .B(p_input[21270]), .Z(n19399) );
  AND U29101 ( .A(n19401), .B(n19402), .Z(o[126]) );
  AND U29102 ( .A(p_input[126]), .B(p_input[10126]), .Z(n19402) );
  AND U29103 ( .A(p_input[30126]), .B(p_input[20126]), .Z(n19401) );
  AND U29104 ( .A(n19403), .B(n19404), .Z(o[1269]) );
  AND U29105 ( .A(p_input[1269]), .B(p_input[11269]), .Z(n19404) );
  AND U29106 ( .A(p_input[31269]), .B(p_input[21269]), .Z(n19403) );
  AND U29107 ( .A(n19405), .B(n19406), .Z(o[1268]) );
  AND U29108 ( .A(p_input[1268]), .B(p_input[11268]), .Z(n19406) );
  AND U29109 ( .A(p_input[31268]), .B(p_input[21268]), .Z(n19405) );
  AND U29110 ( .A(n19407), .B(n19408), .Z(o[1267]) );
  AND U29111 ( .A(p_input[1267]), .B(p_input[11267]), .Z(n19408) );
  AND U29112 ( .A(p_input[31267]), .B(p_input[21267]), .Z(n19407) );
  AND U29113 ( .A(n19409), .B(n19410), .Z(o[1266]) );
  AND U29114 ( .A(p_input[1266]), .B(p_input[11266]), .Z(n19410) );
  AND U29115 ( .A(p_input[31266]), .B(p_input[21266]), .Z(n19409) );
  AND U29116 ( .A(n19411), .B(n19412), .Z(o[1265]) );
  AND U29117 ( .A(p_input[1265]), .B(p_input[11265]), .Z(n19412) );
  AND U29118 ( .A(p_input[31265]), .B(p_input[21265]), .Z(n19411) );
  AND U29119 ( .A(n19413), .B(n19414), .Z(o[1264]) );
  AND U29120 ( .A(p_input[1264]), .B(p_input[11264]), .Z(n19414) );
  AND U29121 ( .A(p_input[31264]), .B(p_input[21264]), .Z(n19413) );
  AND U29122 ( .A(n19415), .B(n19416), .Z(o[1263]) );
  AND U29123 ( .A(p_input[1263]), .B(p_input[11263]), .Z(n19416) );
  AND U29124 ( .A(p_input[31263]), .B(p_input[21263]), .Z(n19415) );
  AND U29125 ( .A(n19417), .B(n19418), .Z(o[1262]) );
  AND U29126 ( .A(p_input[1262]), .B(p_input[11262]), .Z(n19418) );
  AND U29127 ( .A(p_input[31262]), .B(p_input[21262]), .Z(n19417) );
  AND U29128 ( .A(n19419), .B(n19420), .Z(o[1261]) );
  AND U29129 ( .A(p_input[1261]), .B(p_input[11261]), .Z(n19420) );
  AND U29130 ( .A(p_input[31261]), .B(p_input[21261]), .Z(n19419) );
  AND U29131 ( .A(n19421), .B(n19422), .Z(o[1260]) );
  AND U29132 ( .A(p_input[1260]), .B(p_input[11260]), .Z(n19422) );
  AND U29133 ( .A(p_input[31260]), .B(p_input[21260]), .Z(n19421) );
  AND U29134 ( .A(n19423), .B(n19424), .Z(o[125]) );
  AND U29135 ( .A(p_input[125]), .B(p_input[10125]), .Z(n19424) );
  AND U29136 ( .A(p_input[30125]), .B(p_input[20125]), .Z(n19423) );
  AND U29137 ( .A(n19425), .B(n19426), .Z(o[1259]) );
  AND U29138 ( .A(p_input[1259]), .B(p_input[11259]), .Z(n19426) );
  AND U29139 ( .A(p_input[31259]), .B(p_input[21259]), .Z(n19425) );
  AND U29140 ( .A(n19427), .B(n19428), .Z(o[1258]) );
  AND U29141 ( .A(p_input[1258]), .B(p_input[11258]), .Z(n19428) );
  AND U29142 ( .A(p_input[31258]), .B(p_input[21258]), .Z(n19427) );
  AND U29143 ( .A(n19429), .B(n19430), .Z(o[1257]) );
  AND U29144 ( .A(p_input[1257]), .B(p_input[11257]), .Z(n19430) );
  AND U29145 ( .A(p_input[31257]), .B(p_input[21257]), .Z(n19429) );
  AND U29146 ( .A(n19431), .B(n19432), .Z(o[1256]) );
  AND U29147 ( .A(p_input[1256]), .B(p_input[11256]), .Z(n19432) );
  AND U29148 ( .A(p_input[31256]), .B(p_input[21256]), .Z(n19431) );
  AND U29149 ( .A(n19433), .B(n19434), .Z(o[1255]) );
  AND U29150 ( .A(p_input[1255]), .B(p_input[11255]), .Z(n19434) );
  AND U29151 ( .A(p_input[31255]), .B(p_input[21255]), .Z(n19433) );
  AND U29152 ( .A(n19435), .B(n19436), .Z(o[1254]) );
  AND U29153 ( .A(p_input[1254]), .B(p_input[11254]), .Z(n19436) );
  AND U29154 ( .A(p_input[31254]), .B(p_input[21254]), .Z(n19435) );
  AND U29155 ( .A(n19437), .B(n19438), .Z(o[1253]) );
  AND U29156 ( .A(p_input[1253]), .B(p_input[11253]), .Z(n19438) );
  AND U29157 ( .A(p_input[31253]), .B(p_input[21253]), .Z(n19437) );
  AND U29158 ( .A(n19439), .B(n19440), .Z(o[1252]) );
  AND U29159 ( .A(p_input[1252]), .B(p_input[11252]), .Z(n19440) );
  AND U29160 ( .A(p_input[31252]), .B(p_input[21252]), .Z(n19439) );
  AND U29161 ( .A(n19441), .B(n19442), .Z(o[1251]) );
  AND U29162 ( .A(p_input[1251]), .B(p_input[11251]), .Z(n19442) );
  AND U29163 ( .A(p_input[31251]), .B(p_input[21251]), .Z(n19441) );
  AND U29164 ( .A(n19443), .B(n19444), .Z(o[1250]) );
  AND U29165 ( .A(p_input[1250]), .B(p_input[11250]), .Z(n19444) );
  AND U29166 ( .A(p_input[31250]), .B(p_input[21250]), .Z(n19443) );
  AND U29167 ( .A(n19445), .B(n19446), .Z(o[124]) );
  AND U29168 ( .A(p_input[124]), .B(p_input[10124]), .Z(n19446) );
  AND U29169 ( .A(p_input[30124]), .B(p_input[20124]), .Z(n19445) );
  AND U29170 ( .A(n19447), .B(n19448), .Z(o[1249]) );
  AND U29171 ( .A(p_input[1249]), .B(p_input[11249]), .Z(n19448) );
  AND U29172 ( .A(p_input[31249]), .B(p_input[21249]), .Z(n19447) );
  AND U29173 ( .A(n19449), .B(n19450), .Z(o[1248]) );
  AND U29174 ( .A(p_input[1248]), .B(p_input[11248]), .Z(n19450) );
  AND U29175 ( .A(p_input[31248]), .B(p_input[21248]), .Z(n19449) );
  AND U29176 ( .A(n19451), .B(n19452), .Z(o[1247]) );
  AND U29177 ( .A(p_input[1247]), .B(p_input[11247]), .Z(n19452) );
  AND U29178 ( .A(p_input[31247]), .B(p_input[21247]), .Z(n19451) );
  AND U29179 ( .A(n19453), .B(n19454), .Z(o[1246]) );
  AND U29180 ( .A(p_input[1246]), .B(p_input[11246]), .Z(n19454) );
  AND U29181 ( .A(p_input[31246]), .B(p_input[21246]), .Z(n19453) );
  AND U29182 ( .A(n19455), .B(n19456), .Z(o[1245]) );
  AND U29183 ( .A(p_input[1245]), .B(p_input[11245]), .Z(n19456) );
  AND U29184 ( .A(p_input[31245]), .B(p_input[21245]), .Z(n19455) );
  AND U29185 ( .A(n19457), .B(n19458), .Z(o[1244]) );
  AND U29186 ( .A(p_input[1244]), .B(p_input[11244]), .Z(n19458) );
  AND U29187 ( .A(p_input[31244]), .B(p_input[21244]), .Z(n19457) );
  AND U29188 ( .A(n19459), .B(n19460), .Z(o[1243]) );
  AND U29189 ( .A(p_input[1243]), .B(p_input[11243]), .Z(n19460) );
  AND U29190 ( .A(p_input[31243]), .B(p_input[21243]), .Z(n19459) );
  AND U29191 ( .A(n19461), .B(n19462), .Z(o[1242]) );
  AND U29192 ( .A(p_input[1242]), .B(p_input[11242]), .Z(n19462) );
  AND U29193 ( .A(p_input[31242]), .B(p_input[21242]), .Z(n19461) );
  AND U29194 ( .A(n19463), .B(n19464), .Z(o[1241]) );
  AND U29195 ( .A(p_input[1241]), .B(p_input[11241]), .Z(n19464) );
  AND U29196 ( .A(p_input[31241]), .B(p_input[21241]), .Z(n19463) );
  AND U29197 ( .A(n19465), .B(n19466), .Z(o[1240]) );
  AND U29198 ( .A(p_input[1240]), .B(p_input[11240]), .Z(n19466) );
  AND U29199 ( .A(p_input[31240]), .B(p_input[21240]), .Z(n19465) );
  AND U29200 ( .A(n19467), .B(n19468), .Z(o[123]) );
  AND U29201 ( .A(p_input[123]), .B(p_input[10123]), .Z(n19468) );
  AND U29202 ( .A(p_input[30123]), .B(p_input[20123]), .Z(n19467) );
  AND U29203 ( .A(n19469), .B(n19470), .Z(o[1239]) );
  AND U29204 ( .A(p_input[1239]), .B(p_input[11239]), .Z(n19470) );
  AND U29205 ( .A(p_input[31239]), .B(p_input[21239]), .Z(n19469) );
  AND U29206 ( .A(n19471), .B(n19472), .Z(o[1238]) );
  AND U29207 ( .A(p_input[1238]), .B(p_input[11238]), .Z(n19472) );
  AND U29208 ( .A(p_input[31238]), .B(p_input[21238]), .Z(n19471) );
  AND U29209 ( .A(n19473), .B(n19474), .Z(o[1237]) );
  AND U29210 ( .A(p_input[1237]), .B(p_input[11237]), .Z(n19474) );
  AND U29211 ( .A(p_input[31237]), .B(p_input[21237]), .Z(n19473) );
  AND U29212 ( .A(n19475), .B(n19476), .Z(o[1236]) );
  AND U29213 ( .A(p_input[1236]), .B(p_input[11236]), .Z(n19476) );
  AND U29214 ( .A(p_input[31236]), .B(p_input[21236]), .Z(n19475) );
  AND U29215 ( .A(n19477), .B(n19478), .Z(o[1235]) );
  AND U29216 ( .A(p_input[1235]), .B(p_input[11235]), .Z(n19478) );
  AND U29217 ( .A(p_input[31235]), .B(p_input[21235]), .Z(n19477) );
  AND U29218 ( .A(n19479), .B(n19480), .Z(o[1234]) );
  AND U29219 ( .A(p_input[1234]), .B(p_input[11234]), .Z(n19480) );
  AND U29220 ( .A(p_input[31234]), .B(p_input[21234]), .Z(n19479) );
  AND U29221 ( .A(n19481), .B(n19482), .Z(o[1233]) );
  AND U29222 ( .A(p_input[1233]), .B(p_input[11233]), .Z(n19482) );
  AND U29223 ( .A(p_input[31233]), .B(p_input[21233]), .Z(n19481) );
  AND U29224 ( .A(n19483), .B(n19484), .Z(o[1232]) );
  AND U29225 ( .A(p_input[1232]), .B(p_input[11232]), .Z(n19484) );
  AND U29226 ( .A(p_input[31232]), .B(p_input[21232]), .Z(n19483) );
  AND U29227 ( .A(n19485), .B(n19486), .Z(o[1231]) );
  AND U29228 ( .A(p_input[1231]), .B(p_input[11231]), .Z(n19486) );
  AND U29229 ( .A(p_input[31231]), .B(p_input[21231]), .Z(n19485) );
  AND U29230 ( .A(n19487), .B(n19488), .Z(o[1230]) );
  AND U29231 ( .A(p_input[1230]), .B(p_input[11230]), .Z(n19488) );
  AND U29232 ( .A(p_input[31230]), .B(p_input[21230]), .Z(n19487) );
  AND U29233 ( .A(n19489), .B(n19490), .Z(o[122]) );
  AND U29234 ( .A(p_input[122]), .B(p_input[10122]), .Z(n19490) );
  AND U29235 ( .A(p_input[30122]), .B(p_input[20122]), .Z(n19489) );
  AND U29236 ( .A(n19491), .B(n19492), .Z(o[1229]) );
  AND U29237 ( .A(p_input[1229]), .B(p_input[11229]), .Z(n19492) );
  AND U29238 ( .A(p_input[31229]), .B(p_input[21229]), .Z(n19491) );
  AND U29239 ( .A(n19493), .B(n19494), .Z(o[1228]) );
  AND U29240 ( .A(p_input[1228]), .B(p_input[11228]), .Z(n19494) );
  AND U29241 ( .A(p_input[31228]), .B(p_input[21228]), .Z(n19493) );
  AND U29242 ( .A(n19495), .B(n19496), .Z(o[1227]) );
  AND U29243 ( .A(p_input[1227]), .B(p_input[11227]), .Z(n19496) );
  AND U29244 ( .A(p_input[31227]), .B(p_input[21227]), .Z(n19495) );
  AND U29245 ( .A(n19497), .B(n19498), .Z(o[1226]) );
  AND U29246 ( .A(p_input[1226]), .B(p_input[11226]), .Z(n19498) );
  AND U29247 ( .A(p_input[31226]), .B(p_input[21226]), .Z(n19497) );
  AND U29248 ( .A(n19499), .B(n19500), .Z(o[1225]) );
  AND U29249 ( .A(p_input[1225]), .B(p_input[11225]), .Z(n19500) );
  AND U29250 ( .A(p_input[31225]), .B(p_input[21225]), .Z(n19499) );
  AND U29251 ( .A(n19501), .B(n19502), .Z(o[1224]) );
  AND U29252 ( .A(p_input[1224]), .B(p_input[11224]), .Z(n19502) );
  AND U29253 ( .A(p_input[31224]), .B(p_input[21224]), .Z(n19501) );
  AND U29254 ( .A(n19503), .B(n19504), .Z(o[1223]) );
  AND U29255 ( .A(p_input[1223]), .B(p_input[11223]), .Z(n19504) );
  AND U29256 ( .A(p_input[31223]), .B(p_input[21223]), .Z(n19503) );
  AND U29257 ( .A(n19505), .B(n19506), .Z(o[1222]) );
  AND U29258 ( .A(p_input[1222]), .B(p_input[11222]), .Z(n19506) );
  AND U29259 ( .A(p_input[31222]), .B(p_input[21222]), .Z(n19505) );
  AND U29260 ( .A(n19507), .B(n19508), .Z(o[1221]) );
  AND U29261 ( .A(p_input[1221]), .B(p_input[11221]), .Z(n19508) );
  AND U29262 ( .A(p_input[31221]), .B(p_input[21221]), .Z(n19507) );
  AND U29263 ( .A(n19509), .B(n19510), .Z(o[1220]) );
  AND U29264 ( .A(p_input[1220]), .B(p_input[11220]), .Z(n19510) );
  AND U29265 ( .A(p_input[31220]), .B(p_input[21220]), .Z(n19509) );
  AND U29266 ( .A(n19511), .B(n19512), .Z(o[121]) );
  AND U29267 ( .A(p_input[121]), .B(p_input[10121]), .Z(n19512) );
  AND U29268 ( .A(p_input[30121]), .B(p_input[20121]), .Z(n19511) );
  AND U29269 ( .A(n19513), .B(n19514), .Z(o[1219]) );
  AND U29270 ( .A(p_input[1219]), .B(p_input[11219]), .Z(n19514) );
  AND U29271 ( .A(p_input[31219]), .B(p_input[21219]), .Z(n19513) );
  AND U29272 ( .A(n19515), .B(n19516), .Z(o[1218]) );
  AND U29273 ( .A(p_input[1218]), .B(p_input[11218]), .Z(n19516) );
  AND U29274 ( .A(p_input[31218]), .B(p_input[21218]), .Z(n19515) );
  AND U29275 ( .A(n19517), .B(n19518), .Z(o[1217]) );
  AND U29276 ( .A(p_input[1217]), .B(p_input[11217]), .Z(n19518) );
  AND U29277 ( .A(p_input[31217]), .B(p_input[21217]), .Z(n19517) );
  AND U29278 ( .A(n19519), .B(n19520), .Z(o[1216]) );
  AND U29279 ( .A(p_input[1216]), .B(p_input[11216]), .Z(n19520) );
  AND U29280 ( .A(p_input[31216]), .B(p_input[21216]), .Z(n19519) );
  AND U29281 ( .A(n19521), .B(n19522), .Z(o[1215]) );
  AND U29282 ( .A(p_input[1215]), .B(p_input[11215]), .Z(n19522) );
  AND U29283 ( .A(p_input[31215]), .B(p_input[21215]), .Z(n19521) );
  AND U29284 ( .A(n19523), .B(n19524), .Z(o[1214]) );
  AND U29285 ( .A(p_input[1214]), .B(p_input[11214]), .Z(n19524) );
  AND U29286 ( .A(p_input[31214]), .B(p_input[21214]), .Z(n19523) );
  AND U29287 ( .A(n19525), .B(n19526), .Z(o[1213]) );
  AND U29288 ( .A(p_input[1213]), .B(p_input[11213]), .Z(n19526) );
  AND U29289 ( .A(p_input[31213]), .B(p_input[21213]), .Z(n19525) );
  AND U29290 ( .A(n19527), .B(n19528), .Z(o[1212]) );
  AND U29291 ( .A(p_input[1212]), .B(p_input[11212]), .Z(n19528) );
  AND U29292 ( .A(p_input[31212]), .B(p_input[21212]), .Z(n19527) );
  AND U29293 ( .A(n19529), .B(n19530), .Z(o[1211]) );
  AND U29294 ( .A(p_input[1211]), .B(p_input[11211]), .Z(n19530) );
  AND U29295 ( .A(p_input[31211]), .B(p_input[21211]), .Z(n19529) );
  AND U29296 ( .A(n19531), .B(n19532), .Z(o[1210]) );
  AND U29297 ( .A(p_input[1210]), .B(p_input[11210]), .Z(n19532) );
  AND U29298 ( .A(p_input[31210]), .B(p_input[21210]), .Z(n19531) );
  AND U29299 ( .A(n19533), .B(n19534), .Z(o[120]) );
  AND U29300 ( .A(p_input[120]), .B(p_input[10120]), .Z(n19534) );
  AND U29301 ( .A(p_input[30120]), .B(p_input[20120]), .Z(n19533) );
  AND U29302 ( .A(n19535), .B(n19536), .Z(o[1209]) );
  AND U29303 ( .A(p_input[1209]), .B(p_input[11209]), .Z(n19536) );
  AND U29304 ( .A(p_input[31209]), .B(p_input[21209]), .Z(n19535) );
  AND U29305 ( .A(n19537), .B(n19538), .Z(o[1208]) );
  AND U29306 ( .A(p_input[1208]), .B(p_input[11208]), .Z(n19538) );
  AND U29307 ( .A(p_input[31208]), .B(p_input[21208]), .Z(n19537) );
  AND U29308 ( .A(n19539), .B(n19540), .Z(o[1207]) );
  AND U29309 ( .A(p_input[1207]), .B(p_input[11207]), .Z(n19540) );
  AND U29310 ( .A(p_input[31207]), .B(p_input[21207]), .Z(n19539) );
  AND U29311 ( .A(n19541), .B(n19542), .Z(o[1206]) );
  AND U29312 ( .A(p_input[1206]), .B(p_input[11206]), .Z(n19542) );
  AND U29313 ( .A(p_input[31206]), .B(p_input[21206]), .Z(n19541) );
  AND U29314 ( .A(n19543), .B(n19544), .Z(o[1205]) );
  AND U29315 ( .A(p_input[1205]), .B(p_input[11205]), .Z(n19544) );
  AND U29316 ( .A(p_input[31205]), .B(p_input[21205]), .Z(n19543) );
  AND U29317 ( .A(n19545), .B(n19546), .Z(o[1204]) );
  AND U29318 ( .A(p_input[1204]), .B(p_input[11204]), .Z(n19546) );
  AND U29319 ( .A(p_input[31204]), .B(p_input[21204]), .Z(n19545) );
  AND U29320 ( .A(n19547), .B(n19548), .Z(o[1203]) );
  AND U29321 ( .A(p_input[1203]), .B(p_input[11203]), .Z(n19548) );
  AND U29322 ( .A(p_input[31203]), .B(p_input[21203]), .Z(n19547) );
  AND U29323 ( .A(n19549), .B(n19550), .Z(o[1202]) );
  AND U29324 ( .A(p_input[1202]), .B(p_input[11202]), .Z(n19550) );
  AND U29325 ( .A(p_input[31202]), .B(p_input[21202]), .Z(n19549) );
  AND U29326 ( .A(n19551), .B(n19552), .Z(o[1201]) );
  AND U29327 ( .A(p_input[1201]), .B(p_input[11201]), .Z(n19552) );
  AND U29328 ( .A(p_input[31201]), .B(p_input[21201]), .Z(n19551) );
  AND U29329 ( .A(n19553), .B(n19554), .Z(o[1200]) );
  AND U29330 ( .A(p_input[1200]), .B(p_input[11200]), .Z(n19554) );
  AND U29331 ( .A(p_input[31200]), .B(p_input[21200]), .Z(n19553) );
  AND U29332 ( .A(n19555), .B(n19556), .Z(o[11]) );
  AND U29333 ( .A(p_input[11]), .B(p_input[10011]), .Z(n19556) );
  AND U29334 ( .A(p_input[30011]), .B(p_input[20011]), .Z(n19555) );
  AND U29335 ( .A(n19557), .B(n19558), .Z(o[119]) );
  AND U29336 ( .A(p_input[119]), .B(p_input[10119]), .Z(n19558) );
  AND U29337 ( .A(p_input[30119]), .B(p_input[20119]), .Z(n19557) );
  AND U29338 ( .A(n19559), .B(n19560), .Z(o[1199]) );
  AND U29339 ( .A(p_input[1199]), .B(p_input[11199]), .Z(n19560) );
  AND U29340 ( .A(p_input[31199]), .B(p_input[21199]), .Z(n19559) );
  AND U29341 ( .A(n19561), .B(n19562), .Z(o[1198]) );
  AND U29342 ( .A(p_input[1198]), .B(p_input[11198]), .Z(n19562) );
  AND U29343 ( .A(p_input[31198]), .B(p_input[21198]), .Z(n19561) );
  AND U29344 ( .A(n19563), .B(n19564), .Z(o[1197]) );
  AND U29345 ( .A(p_input[1197]), .B(p_input[11197]), .Z(n19564) );
  AND U29346 ( .A(p_input[31197]), .B(p_input[21197]), .Z(n19563) );
  AND U29347 ( .A(n19565), .B(n19566), .Z(o[1196]) );
  AND U29348 ( .A(p_input[1196]), .B(p_input[11196]), .Z(n19566) );
  AND U29349 ( .A(p_input[31196]), .B(p_input[21196]), .Z(n19565) );
  AND U29350 ( .A(n19567), .B(n19568), .Z(o[1195]) );
  AND U29351 ( .A(p_input[1195]), .B(p_input[11195]), .Z(n19568) );
  AND U29352 ( .A(p_input[31195]), .B(p_input[21195]), .Z(n19567) );
  AND U29353 ( .A(n19569), .B(n19570), .Z(o[1194]) );
  AND U29354 ( .A(p_input[1194]), .B(p_input[11194]), .Z(n19570) );
  AND U29355 ( .A(p_input[31194]), .B(p_input[21194]), .Z(n19569) );
  AND U29356 ( .A(n19571), .B(n19572), .Z(o[1193]) );
  AND U29357 ( .A(p_input[1193]), .B(p_input[11193]), .Z(n19572) );
  AND U29358 ( .A(p_input[31193]), .B(p_input[21193]), .Z(n19571) );
  AND U29359 ( .A(n19573), .B(n19574), .Z(o[1192]) );
  AND U29360 ( .A(p_input[1192]), .B(p_input[11192]), .Z(n19574) );
  AND U29361 ( .A(p_input[31192]), .B(p_input[21192]), .Z(n19573) );
  AND U29362 ( .A(n19575), .B(n19576), .Z(o[1191]) );
  AND U29363 ( .A(p_input[1191]), .B(p_input[11191]), .Z(n19576) );
  AND U29364 ( .A(p_input[31191]), .B(p_input[21191]), .Z(n19575) );
  AND U29365 ( .A(n19577), .B(n19578), .Z(o[1190]) );
  AND U29366 ( .A(p_input[1190]), .B(p_input[11190]), .Z(n19578) );
  AND U29367 ( .A(p_input[31190]), .B(p_input[21190]), .Z(n19577) );
  AND U29368 ( .A(n19579), .B(n19580), .Z(o[118]) );
  AND U29369 ( .A(p_input[118]), .B(p_input[10118]), .Z(n19580) );
  AND U29370 ( .A(p_input[30118]), .B(p_input[20118]), .Z(n19579) );
  AND U29371 ( .A(n19581), .B(n19582), .Z(o[1189]) );
  AND U29372 ( .A(p_input[1189]), .B(p_input[11189]), .Z(n19582) );
  AND U29373 ( .A(p_input[31189]), .B(p_input[21189]), .Z(n19581) );
  AND U29374 ( .A(n19583), .B(n19584), .Z(o[1188]) );
  AND U29375 ( .A(p_input[1188]), .B(p_input[11188]), .Z(n19584) );
  AND U29376 ( .A(p_input[31188]), .B(p_input[21188]), .Z(n19583) );
  AND U29377 ( .A(n19585), .B(n19586), .Z(o[1187]) );
  AND U29378 ( .A(p_input[1187]), .B(p_input[11187]), .Z(n19586) );
  AND U29379 ( .A(p_input[31187]), .B(p_input[21187]), .Z(n19585) );
  AND U29380 ( .A(n19587), .B(n19588), .Z(o[1186]) );
  AND U29381 ( .A(p_input[1186]), .B(p_input[11186]), .Z(n19588) );
  AND U29382 ( .A(p_input[31186]), .B(p_input[21186]), .Z(n19587) );
  AND U29383 ( .A(n19589), .B(n19590), .Z(o[1185]) );
  AND U29384 ( .A(p_input[1185]), .B(p_input[11185]), .Z(n19590) );
  AND U29385 ( .A(p_input[31185]), .B(p_input[21185]), .Z(n19589) );
  AND U29386 ( .A(n19591), .B(n19592), .Z(o[1184]) );
  AND U29387 ( .A(p_input[1184]), .B(p_input[11184]), .Z(n19592) );
  AND U29388 ( .A(p_input[31184]), .B(p_input[21184]), .Z(n19591) );
  AND U29389 ( .A(n19593), .B(n19594), .Z(o[1183]) );
  AND U29390 ( .A(p_input[1183]), .B(p_input[11183]), .Z(n19594) );
  AND U29391 ( .A(p_input[31183]), .B(p_input[21183]), .Z(n19593) );
  AND U29392 ( .A(n19595), .B(n19596), .Z(o[1182]) );
  AND U29393 ( .A(p_input[1182]), .B(p_input[11182]), .Z(n19596) );
  AND U29394 ( .A(p_input[31182]), .B(p_input[21182]), .Z(n19595) );
  AND U29395 ( .A(n19597), .B(n19598), .Z(o[1181]) );
  AND U29396 ( .A(p_input[1181]), .B(p_input[11181]), .Z(n19598) );
  AND U29397 ( .A(p_input[31181]), .B(p_input[21181]), .Z(n19597) );
  AND U29398 ( .A(n19599), .B(n19600), .Z(o[1180]) );
  AND U29399 ( .A(p_input[1180]), .B(p_input[11180]), .Z(n19600) );
  AND U29400 ( .A(p_input[31180]), .B(p_input[21180]), .Z(n19599) );
  AND U29401 ( .A(n19601), .B(n19602), .Z(o[117]) );
  AND U29402 ( .A(p_input[117]), .B(p_input[10117]), .Z(n19602) );
  AND U29403 ( .A(p_input[30117]), .B(p_input[20117]), .Z(n19601) );
  AND U29404 ( .A(n19603), .B(n19604), .Z(o[1179]) );
  AND U29405 ( .A(p_input[1179]), .B(p_input[11179]), .Z(n19604) );
  AND U29406 ( .A(p_input[31179]), .B(p_input[21179]), .Z(n19603) );
  AND U29407 ( .A(n19605), .B(n19606), .Z(o[1178]) );
  AND U29408 ( .A(p_input[1178]), .B(p_input[11178]), .Z(n19606) );
  AND U29409 ( .A(p_input[31178]), .B(p_input[21178]), .Z(n19605) );
  AND U29410 ( .A(n19607), .B(n19608), .Z(o[1177]) );
  AND U29411 ( .A(p_input[1177]), .B(p_input[11177]), .Z(n19608) );
  AND U29412 ( .A(p_input[31177]), .B(p_input[21177]), .Z(n19607) );
  AND U29413 ( .A(n19609), .B(n19610), .Z(o[1176]) );
  AND U29414 ( .A(p_input[1176]), .B(p_input[11176]), .Z(n19610) );
  AND U29415 ( .A(p_input[31176]), .B(p_input[21176]), .Z(n19609) );
  AND U29416 ( .A(n19611), .B(n19612), .Z(o[1175]) );
  AND U29417 ( .A(p_input[1175]), .B(p_input[11175]), .Z(n19612) );
  AND U29418 ( .A(p_input[31175]), .B(p_input[21175]), .Z(n19611) );
  AND U29419 ( .A(n19613), .B(n19614), .Z(o[1174]) );
  AND U29420 ( .A(p_input[1174]), .B(p_input[11174]), .Z(n19614) );
  AND U29421 ( .A(p_input[31174]), .B(p_input[21174]), .Z(n19613) );
  AND U29422 ( .A(n19615), .B(n19616), .Z(o[1173]) );
  AND U29423 ( .A(p_input[1173]), .B(p_input[11173]), .Z(n19616) );
  AND U29424 ( .A(p_input[31173]), .B(p_input[21173]), .Z(n19615) );
  AND U29425 ( .A(n19617), .B(n19618), .Z(o[1172]) );
  AND U29426 ( .A(p_input[1172]), .B(p_input[11172]), .Z(n19618) );
  AND U29427 ( .A(p_input[31172]), .B(p_input[21172]), .Z(n19617) );
  AND U29428 ( .A(n19619), .B(n19620), .Z(o[1171]) );
  AND U29429 ( .A(p_input[1171]), .B(p_input[11171]), .Z(n19620) );
  AND U29430 ( .A(p_input[31171]), .B(p_input[21171]), .Z(n19619) );
  AND U29431 ( .A(n19621), .B(n19622), .Z(o[1170]) );
  AND U29432 ( .A(p_input[1170]), .B(p_input[11170]), .Z(n19622) );
  AND U29433 ( .A(p_input[31170]), .B(p_input[21170]), .Z(n19621) );
  AND U29434 ( .A(n19623), .B(n19624), .Z(o[116]) );
  AND U29435 ( .A(p_input[116]), .B(p_input[10116]), .Z(n19624) );
  AND U29436 ( .A(p_input[30116]), .B(p_input[20116]), .Z(n19623) );
  AND U29437 ( .A(n19625), .B(n19626), .Z(o[1169]) );
  AND U29438 ( .A(p_input[1169]), .B(p_input[11169]), .Z(n19626) );
  AND U29439 ( .A(p_input[31169]), .B(p_input[21169]), .Z(n19625) );
  AND U29440 ( .A(n19627), .B(n19628), .Z(o[1168]) );
  AND U29441 ( .A(p_input[1168]), .B(p_input[11168]), .Z(n19628) );
  AND U29442 ( .A(p_input[31168]), .B(p_input[21168]), .Z(n19627) );
  AND U29443 ( .A(n19629), .B(n19630), .Z(o[1167]) );
  AND U29444 ( .A(p_input[1167]), .B(p_input[11167]), .Z(n19630) );
  AND U29445 ( .A(p_input[31167]), .B(p_input[21167]), .Z(n19629) );
  AND U29446 ( .A(n19631), .B(n19632), .Z(o[1166]) );
  AND U29447 ( .A(p_input[1166]), .B(p_input[11166]), .Z(n19632) );
  AND U29448 ( .A(p_input[31166]), .B(p_input[21166]), .Z(n19631) );
  AND U29449 ( .A(n19633), .B(n19634), .Z(o[1165]) );
  AND U29450 ( .A(p_input[1165]), .B(p_input[11165]), .Z(n19634) );
  AND U29451 ( .A(p_input[31165]), .B(p_input[21165]), .Z(n19633) );
  AND U29452 ( .A(n19635), .B(n19636), .Z(o[1164]) );
  AND U29453 ( .A(p_input[1164]), .B(p_input[11164]), .Z(n19636) );
  AND U29454 ( .A(p_input[31164]), .B(p_input[21164]), .Z(n19635) );
  AND U29455 ( .A(n19637), .B(n19638), .Z(o[1163]) );
  AND U29456 ( .A(p_input[1163]), .B(p_input[11163]), .Z(n19638) );
  AND U29457 ( .A(p_input[31163]), .B(p_input[21163]), .Z(n19637) );
  AND U29458 ( .A(n19639), .B(n19640), .Z(o[1162]) );
  AND U29459 ( .A(p_input[1162]), .B(p_input[11162]), .Z(n19640) );
  AND U29460 ( .A(p_input[31162]), .B(p_input[21162]), .Z(n19639) );
  AND U29461 ( .A(n19641), .B(n19642), .Z(o[1161]) );
  AND U29462 ( .A(p_input[1161]), .B(p_input[11161]), .Z(n19642) );
  AND U29463 ( .A(p_input[31161]), .B(p_input[21161]), .Z(n19641) );
  AND U29464 ( .A(n19643), .B(n19644), .Z(o[1160]) );
  AND U29465 ( .A(p_input[1160]), .B(p_input[11160]), .Z(n19644) );
  AND U29466 ( .A(p_input[31160]), .B(p_input[21160]), .Z(n19643) );
  AND U29467 ( .A(n19645), .B(n19646), .Z(o[115]) );
  AND U29468 ( .A(p_input[115]), .B(p_input[10115]), .Z(n19646) );
  AND U29469 ( .A(p_input[30115]), .B(p_input[20115]), .Z(n19645) );
  AND U29470 ( .A(n19647), .B(n19648), .Z(o[1159]) );
  AND U29471 ( .A(p_input[1159]), .B(p_input[11159]), .Z(n19648) );
  AND U29472 ( .A(p_input[31159]), .B(p_input[21159]), .Z(n19647) );
  AND U29473 ( .A(n19649), .B(n19650), .Z(o[1158]) );
  AND U29474 ( .A(p_input[1158]), .B(p_input[11158]), .Z(n19650) );
  AND U29475 ( .A(p_input[31158]), .B(p_input[21158]), .Z(n19649) );
  AND U29476 ( .A(n19651), .B(n19652), .Z(o[1157]) );
  AND U29477 ( .A(p_input[1157]), .B(p_input[11157]), .Z(n19652) );
  AND U29478 ( .A(p_input[31157]), .B(p_input[21157]), .Z(n19651) );
  AND U29479 ( .A(n19653), .B(n19654), .Z(o[1156]) );
  AND U29480 ( .A(p_input[1156]), .B(p_input[11156]), .Z(n19654) );
  AND U29481 ( .A(p_input[31156]), .B(p_input[21156]), .Z(n19653) );
  AND U29482 ( .A(n19655), .B(n19656), .Z(o[1155]) );
  AND U29483 ( .A(p_input[1155]), .B(p_input[11155]), .Z(n19656) );
  AND U29484 ( .A(p_input[31155]), .B(p_input[21155]), .Z(n19655) );
  AND U29485 ( .A(n19657), .B(n19658), .Z(o[1154]) );
  AND U29486 ( .A(p_input[1154]), .B(p_input[11154]), .Z(n19658) );
  AND U29487 ( .A(p_input[31154]), .B(p_input[21154]), .Z(n19657) );
  AND U29488 ( .A(n19659), .B(n19660), .Z(o[1153]) );
  AND U29489 ( .A(p_input[1153]), .B(p_input[11153]), .Z(n19660) );
  AND U29490 ( .A(p_input[31153]), .B(p_input[21153]), .Z(n19659) );
  AND U29491 ( .A(n19661), .B(n19662), .Z(o[1152]) );
  AND U29492 ( .A(p_input[1152]), .B(p_input[11152]), .Z(n19662) );
  AND U29493 ( .A(p_input[31152]), .B(p_input[21152]), .Z(n19661) );
  AND U29494 ( .A(n19663), .B(n19664), .Z(o[1151]) );
  AND U29495 ( .A(p_input[1151]), .B(p_input[11151]), .Z(n19664) );
  AND U29496 ( .A(p_input[31151]), .B(p_input[21151]), .Z(n19663) );
  AND U29497 ( .A(n19665), .B(n19666), .Z(o[1150]) );
  AND U29498 ( .A(p_input[1150]), .B(p_input[11150]), .Z(n19666) );
  AND U29499 ( .A(p_input[31150]), .B(p_input[21150]), .Z(n19665) );
  AND U29500 ( .A(n19667), .B(n19668), .Z(o[114]) );
  AND U29501 ( .A(p_input[114]), .B(p_input[10114]), .Z(n19668) );
  AND U29502 ( .A(p_input[30114]), .B(p_input[20114]), .Z(n19667) );
  AND U29503 ( .A(n19669), .B(n19670), .Z(o[1149]) );
  AND U29504 ( .A(p_input[1149]), .B(p_input[11149]), .Z(n19670) );
  AND U29505 ( .A(p_input[31149]), .B(p_input[21149]), .Z(n19669) );
  AND U29506 ( .A(n19671), .B(n19672), .Z(o[1148]) );
  AND U29507 ( .A(p_input[1148]), .B(p_input[11148]), .Z(n19672) );
  AND U29508 ( .A(p_input[31148]), .B(p_input[21148]), .Z(n19671) );
  AND U29509 ( .A(n19673), .B(n19674), .Z(o[1147]) );
  AND U29510 ( .A(p_input[1147]), .B(p_input[11147]), .Z(n19674) );
  AND U29511 ( .A(p_input[31147]), .B(p_input[21147]), .Z(n19673) );
  AND U29512 ( .A(n19675), .B(n19676), .Z(o[1146]) );
  AND U29513 ( .A(p_input[1146]), .B(p_input[11146]), .Z(n19676) );
  AND U29514 ( .A(p_input[31146]), .B(p_input[21146]), .Z(n19675) );
  AND U29515 ( .A(n19677), .B(n19678), .Z(o[1145]) );
  AND U29516 ( .A(p_input[1145]), .B(p_input[11145]), .Z(n19678) );
  AND U29517 ( .A(p_input[31145]), .B(p_input[21145]), .Z(n19677) );
  AND U29518 ( .A(n19679), .B(n19680), .Z(o[1144]) );
  AND U29519 ( .A(p_input[1144]), .B(p_input[11144]), .Z(n19680) );
  AND U29520 ( .A(p_input[31144]), .B(p_input[21144]), .Z(n19679) );
  AND U29521 ( .A(n19681), .B(n19682), .Z(o[1143]) );
  AND U29522 ( .A(p_input[1143]), .B(p_input[11143]), .Z(n19682) );
  AND U29523 ( .A(p_input[31143]), .B(p_input[21143]), .Z(n19681) );
  AND U29524 ( .A(n19683), .B(n19684), .Z(o[1142]) );
  AND U29525 ( .A(p_input[1142]), .B(p_input[11142]), .Z(n19684) );
  AND U29526 ( .A(p_input[31142]), .B(p_input[21142]), .Z(n19683) );
  AND U29527 ( .A(n19685), .B(n19686), .Z(o[1141]) );
  AND U29528 ( .A(p_input[1141]), .B(p_input[11141]), .Z(n19686) );
  AND U29529 ( .A(p_input[31141]), .B(p_input[21141]), .Z(n19685) );
  AND U29530 ( .A(n19687), .B(n19688), .Z(o[1140]) );
  AND U29531 ( .A(p_input[1140]), .B(p_input[11140]), .Z(n19688) );
  AND U29532 ( .A(p_input[31140]), .B(p_input[21140]), .Z(n19687) );
  AND U29533 ( .A(n19689), .B(n19690), .Z(o[113]) );
  AND U29534 ( .A(p_input[113]), .B(p_input[10113]), .Z(n19690) );
  AND U29535 ( .A(p_input[30113]), .B(p_input[20113]), .Z(n19689) );
  AND U29536 ( .A(n19691), .B(n19692), .Z(o[1139]) );
  AND U29537 ( .A(p_input[1139]), .B(p_input[11139]), .Z(n19692) );
  AND U29538 ( .A(p_input[31139]), .B(p_input[21139]), .Z(n19691) );
  AND U29539 ( .A(n19693), .B(n19694), .Z(o[1138]) );
  AND U29540 ( .A(p_input[1138]), .B(p_input[11138]), .Z(n19694) );
  AND U29541 ( .A(p_input[31138]), .B(p_input[21138]), .Z(n19693) );
  AND U29542 ( .A(n19695), .B(n19696), .Z(o[1137]) );
  AND U29543 ( .A(p_input[1137]), .B(p_input[11137]), .Z(n19696) );
  AND U29544 ( .A(p_input[31137]), .B(p_input[21137]), .Z(n19695) );
  AND U29545 ( .A(n19697), .B(n19698), .Z(o[1136]) );
  AND U29546 ( .A(p_input[1136]), .B(p_input[11136]), .Z(n19698) );
  AND U29547 ( .A(p_input[31136]), .B(p_input[21136]), .Z(n19697) );
  AND U29548 ( .A(n19699), .B(n19700), .Z(o[1135]) );
  AND U29549 ( .A(p_input[1135]), .B(p_input[11135]), .Z(n19700) );
  AND U29550 ( .A(p_input[31135]), .B(p_input[21135]), .Z(n19699) );
  AND U29551 ( .A(n19701), .B(n19702), .Z(o[1134]) );
  AND U29552 ( .A(p_input[1134]), .B(p_input[11134]), .Z(n19702) );
  AND U29553 ( .A(p_input[31134]), .B(p_input[21134]), .Z(n19701) );
  AND U29554 ( .A(n19703), .B(n19704), .Z(o[1133]) );
  AND U29555 ( .A(p_input[1133]), .B(p_input[11133]), .Z(n19704) );
  AND U29556 ( .A(p_input[31133]), .B(p_input[21133]), .Z(n19703) );
  AND U29557 ( .A(n19705), .B(n19706), .Z(o[1132]) );
  AND U29558 ( .A(p_input[1132]), .B(p_input[11132]), .Z(n19706) );
  AND U29559 ( .A(p_input[31132]), .B(p_input[21132]), .Z(n19705) );
  AND U29560 ( .A(n19707), .B(n19708), .Z(o[1131]) );
  AND U29561 ( .A(p_input[1131]), .B(p_input[11131]), .Z(n19708) );
  AND U29562 ( .A(p_input[31131]), .B(p_input[21131]), .Z(n19707) );
  AND U29563 ( .A(n19709), .B(n19710), .Z(o[1130]) );
  AND U29564 ( .A(p_input[1130]), .B(p_input[11130]), .Z(n19710) );
  AND U29565 ( .A(p_input[31130]), .B(p_input[21130]), .Z(n19709) );
  AND U29566 ( .A(n19711), .B(n19712), .Z(o[112]) );
  AND U29567 ( .A(p_input[112]), .B(p_input[10112]), .Z(n19712) );
  AND U29568 ( .A(p_input[30112]), .B(p_input[20112]), .Z(n19711) );
  AND U29569 ( .A(n19713), .B(n19714), .Z(o[1129]) );
  AND U29570 ( .A(p_input[1129]), .B(p_input[11129]), .Z(n19714) );
  AND U29571 ( .A(p_input[31129]), .B(p_input[21129]), .Z(n19713) );
  AND U29572 ( .A(n19715), .B(n19716), .Z(o[1128]) );
  AND U29573 ( .A(p_input[1128]), .B(p_input[11128]), .Z(n19716) );
  AND U29574 ( .A(p_input[31128]), .B(p_input[21128]), .Z(n19715) );
  AND U29575 ( .A(n19717), .B(n19718), .Z(o[1127]) );
  AND U29576 ( .A(p_input[1127]), .B(p_input[11127]), .Z(n19718) );
  AND U29577 ( .A(p_input[31127]), .B(p_input[21127]), .Z(n19717) );
  AND U29578 ( .A(n19719), .B(n19720), .Z(o[1126]) );
  AND U29579 ( .A(p_input[1126]), .B(p_input[11126]), .Z(n19720) );
  AND U29580 ( .A(p_input[31126]), .B(p_input[21126]), .Z(n19719) );
  AND U29581 ( .A(n19721), .B(n19722), .Z(o[1125]) );
  AND U29582 ( .A(p_input[1125]), .B(p_input[11125]), .Z(n19722) );
  AND U29583 ( .A(p_input[31125]), .B(p_input[21125]), .Z(n19721) );
  AND U29584 ( .A(n19723), .B(n19724), .Z(o[1124]) );
  AND U29585 ( .A(p_input[1124]), .B(p_input[11124]), .Z(n19724) );
  AND U29586 ( .A(p_input[31124]), .B(p_input[21124]), .Z(n19723) );
  AND U29587 ( .A(n19725), .B(n19726), .Z(o[1123]) );
  AND U29588 ( .A(p_input[1123]), .B(p_input[11123]), .Z(n19726) );
  AND U29589 ( .A(p_input[31123]), .B(p_input[21123]), .Z(n19725) );
  AND U29590 ( .A(n19727), .B(n19728), .Z(o[1122]) );
  AND U29591 ( .A(p_input[1122]), .B(p_input[11122]), .Z(n19728) );
  AND U29592 ( .A(p_input[31122]), .B(p_input[21122]), .Z(n19727) );
  AND U29593 ( .A(n19729), .B(n19730), .Z(o[1121]) );
  AND U29594 ( .A(p_input[1121]), .B(p_input[11121]), .Z(n19730) );
  AND U29595 ( .A(p_input[31121]), .B(p_input[21121]), .Z(n19729) );
  AND U29596 ( .A(n19731), .B(n19732), .Z(o[1120]) );
  AND U29597 ( .A(p_input[1120]), .B(p_input[11120]), .Z(n19732) );
  AND U29598 ( .A(p_input[31120]), .B(p_input[21120]), .Z(n19731) );
  AND U29599 ( .A(n19733), .B(n19734), .Z(o[111]) );
  AND U29600 ( .A(p_input[111]), .B(p_input[10111]), .Z(n19734) );
  AND U29601 ( .A(p_input[30111]), .B(p_input[20111]), .Z(n19733) );
  AND U29602 ( .A(n19735), .B(n19736), .Z(o[1119]) );
  AND U29603 ( .A(p_input[1119]), .B(p_input[11119]), .Z(n19736) );
  AND U29604 ( .A(p_input[31119]), .B(p_input[21119]), .Z(n19735) );
  AND U29605 ( .A(n19737), .B(n19738), .Z(o[1118]) );
  AND U29606 ( .A(p_input[1118]), .B(p_input[11118]), .Z(n19738) );
  AND U29607 ( .A(p_input[31118]), .B(p_input[21118]), .Z(n19737) );
  AND U29608 ( .A(n19739), .B(n19740), .Z(o[1117]) );
  AND U29609 ( .A(p_input[1117]), .B(p_input[11117]), .Z(n19740) );
  AND U29610 ( .A(p_input[31117]), .B(p_input[21117]), .Z(n19739) );
  AND U29611 ( .A(n19741), .B(n19742), .Z(o[1116]) );
  AND U29612 ( .A(p_input[1116]), .B(p_input[11116]), .Z(n19742) );
  AND U29613 ( .A(p_input[31116]), .B(p_input[21116]), .Z(n19741) );
  AND U29614 ( .A(n19743), .B(n19744), .Z(o[1115]) );
  AND U29615 ( .A(p_input[1115]), .B(p_input[11115]), .Z(n19744) );
  AND U29616 ( .A(p_input[31115]), .B(p_input[21115]), .Z(n19743) );
  AND U29617 ( .A(n19745), .B(n19746), .Z(o[1114]) );
  AND U29618 ( .A(p_input[1114]), .B(p_input[11114]), .Z(n19746) );
  AND U29619 ( .A(p_input[31114]), .B(p_input[21114]), .Z(n19745) );
  AND U29620 ( .A(n19747), .B(n19748), .Z(o[1113]) );
  AND U29621 ( .A(p_input[1113]), .B(p_input[11113]), .Z(n19748) );
  AND U29622 ( .A(p_input[31113]), .B(p_input[21113]), .Z(n19747) );
  AND U29623 ( .A(n19749), .B(n19750), .Z(o[1112]) );
  AND U29624 ( .A(p_input[1112]), .B(p_input[11112]), .Z(n19750) );
  AND U29625 ( .A(p_input[31112]), .B(p_input[21112]), .Z(n19749) );
  AND U29626 ( .A(n19751), .B(n19752), .Z(o[1111]) );
  AND U29627 ( .A(p_input[1111]), .B(p_input[11111]), .Z(n19752) );
  AND U29628 ( .A(p_input[31111]), .B(p_input[21111]), .Z(n19751) );
  AND U29629 ( .A(n19753), .B(n19754), .Z(o[1110]) );
  AND U29630 ( .A(p_input[11110]), .B(p_input[1110]), .Z(n19754) );
  AND U29631 ( .A(p_input[31110]), .B(p_input[21110]), .Z(n19753) );
  AND U29632 ( .A(n19755), .B(n19756), .Z(o[110]) );
  AND U29633 ( .A(p_input[110]), .B(p_input[10110]), .Z(n19756) );
  AND U29634 ( .A(p_input[30110]), .B(p_input[20110]), .Z(n19755) );
  AND U29635 ( .A(n19757), .B(n19758), .Z(o[1109]) );
  AND U29636 ( .A(p_input[11109]), .B(p_input[1109]), .Z(n19758) );
  AND U29637 ( .A(p_input[31109]), .B(p_input[21109]), .Z(n19757) );
  AND U29638 ( .A(n19759), .B(n19760), .Z(o[1108]) );
  AND U29639 ( .A(p_input[11108]), .B(p_input[1108]), .Z(n19760) );
  AND U29640 ( .A(p_input[31108]), .B(p_input[21108]), .Z(n19759) );
  AND U29641 ( .A(n19761), .B(n19762), .Z(o[1107]) );
  AND U29642 ( .A(p_input[11107]), .B(p_input[1107]), .Z(n19762) );
  AND U29643 ( .A(p_input[31107]), .B(p_input[21107]), .Z(n19761) );
  AND U29644 ( .A(n19763), .B(n19764), .Z(o[1106]) );
  AND U29645 ( .A(p_input[11106]), .B(p_input[1106]), .Z(n19764) );
  AND U29646 ( .A(p_input[31106]), .B(p_input[21106]), .Z(n19763) );
  AND U29647 ( .A(n19765), .B(n19766), .Z(o[1105]) );
  AND U29648 ( .A(p_input[11105]), .B(p_input[1105]), .Z(n19766) );
  AND U29649 ( .A(p_input[31105]), .B(p_input[21105]), .Z(n19765) );
  AND U29650 ( .A(n19767), .B(n19768), .Z(o[1104]) );
  AND U29651 ( .A(p_input[11104]), .B(p_input[1104]), .Z(n19768) );
  AND U29652 ( .A(p_input[31104]), .B(p_input[21104]), .Z(n19767) );
  AND U29653 ( .A(n19769), .B(n19770), .Z(o[1103]) );
  AND U29654 ( .A(p_input[11103]), .B(p_input[1103]), .Z(n19770) );
  AND U29655 ( .A(p_input[31103]), .B(p_input[21103]), .Z(n19769) );
  AND U29656 ( .A(n19771), .B(n19772), .Z(o[1102]) );
  AND U29657 ( .A(p_input[11102]), .B(p_input[1102]), .Z(n19772) );
  AND U29658 ( .A(p_input[31102]), .B(p_input[21102]), .Z(n19771) );
  AND U29659 ( .A(n19773), .B(n19774), .Z(o[1101]) );
  AND U29660 ( .A(p_input[11101]), .B(p_input[1101]), .Z(n19774) );
  AND U29661 ( .A(p_input[31101]), .B(p_input[21101]), .Z(n19773) );
  AND U29662 ( .A(n19775), .B(n19776), .Z(o[1100]) );
  AND U29663 ( .A(p_input[11100]), .B(p_input[1100]), .Z(n19776) );
  AND U29664 ( .A(p_input[31100]), .B(p_input[21100]), .Z(n19775) );
  AND U29665 ( .A(n19777), .B(n19778), .Z(o[10]) );
  AND U29666 ( .A(p_input[10]), .B(p_input[10010]), .Z(n19778) );
  AND U29667 ( .A(p_input[30010]), .B(p_input[20010]), .Z(n19777) );
  AND U29668 ( .A(n19779), .B(n19780), .Z(o[109]) );
  AND U29669 ( .A(p_input[109]), .B(p_input[10109]), .Z(n19780) );
  AND U29670 ( .A(p_input[30109]), .B(p_input[20109]), .Z(n19779) );
  AND U29671 ( .A(n19781), .B(n19782), .Z(o[1099]) );
  AND U29672 ( .A(p_input[11099]), .B(p_input[1099]), .Z(n19782) );
  AND U29673 ( .A(p_input[31099]), .B(p_input[21099]), .Z(n19781) );
  AND U29674 ( .A(n19783), .B(n19784), .Z(o[1098]) );
  AND U29675 ( .A(p_input[11098]), .B(p_input[1098]), .Z(n19784) );
  AND U29676 ( .A(p_input[31098]), .B(p_input[21098]), .Z(n19783) );
  AND U29677 ( .A(n19785), .B(n19786), .Z(o[1097]) );
  AND U29678 ( .A(p_input[11097]), .B(p_input[1097]), .Z(n19786) );
  AND U29679 ( .A(p_input[31097]), .B(p_input[21097]), .Z(n19785) );
  AND U29680 ( .A(n19787), .B(n19788), .Z(o[1096]) );
  AND U29681 ( .A(p_input[11096]), .B(p_input[1096]), .Z(n19788) );
  AND U29682 ( .A(p_input[31096]), .B(p_input[21096]), .Z(n19787) );
  AND U29683 ( .A(n19789), .B(n19790), .Z(o[1095]) );
  AND U29684 ( .A(p_input[11095]), .B(p_input[1095]), .Z(n19790) );
  AND U29685 ( .A(p_input[31095]), .B(p_input[21095]), .Z(n19789) );
  AND U29686 ( .A(n19791), .B(n19792), .Z(o[1094]) );
  AND U29687 ( .A(p_input[11094]), .B(p_input[1094]), .Z(n19792) );
  AND U29688 ( .A(p_input[31094]), .B(p_input[21094]), .Z(n19791) );
  AND U29689 ( .A(n19793), .B(n19794), .Z(o[1093]) );
  AND U29690 ( .A(p_input[11093]), .B(p_input[1093]), .Z(n19794) );
  AND U29691 ( .A(p_input[31093]), .B(p_input[21093]), .Z(n19793) );
  AND U29692 ( .A(n19795), .B(n19796), .Z(o[1092]) );
  AND U29693 ( .A(p_input[11092]), .B(p_input[1092]), .Z(n19796) );
  AND U29694 ( .A(p_input[31092]), .B(p_input[21092]), .Z(n19795) );
  AND U29695 ( .A(n19797), .B(n19798), .Z(o[1091]) );
  AND U29696 ( .A(p_input[11091]), .B(p_input[1091]), .Z(n19798) );
  AND U29697 ( .A(p_input[31091]), .B(p_input[21091]), .Z(n19797) );
  AND U29698 ( .A(n19799), .B(n19800), .Z(o[1090]) );
  AND U29699 ( .A(p_input[11090]), .B(p_input[1090]), .Z(n19800) );
  AND U29700 ( .A(p_input[31090]), .B(p_input[21090]), .Z(n19799) );
  AND U29701 ( .A(n19801), .B(n19802), .Z(o[108]) );
  AND U29702 ( .A(p_input[108]), .B(p_input[10108]), .Z(n19802) );
  AND U29703 ( .A(p_input[30108]), .B(p_input[20108]), .Z(n19801) );
  AND U29704 ( .A(n19803), .B(n19804), .Z(o[1089]) );
  AND U29705 ( .A(p_input[11089]), .B(p_input[1089]), .Z(n19804) );
  AND U29706 ( .A(p_input[31089]), .B(p_input[21089]), .Z(n19803) );
  AND U29707 ( .A(n19805), .B(n19806), .Z(o[1088]) );
  AND U29708 ( .A(p_input[11088]), .B(p_input[1088]), .Z(n19806) );
  AND U29709 ( .A(p_input[31088]), .B(p_input[21088]), .Z(n19805) );
  AND U29710 ( .A(n19807), .B(n19808), .Z(o[1087]) );
  AND U29711 ( .A(p_input[11087]), .B(p_input[1087]), .Z(n19808) );
  AND U29712 ( .A(p_input[31087]), .B(p_input[21087]), .Z(n19807) );
  AND U29713 ( .A(n19809), .B(n19810), .Z(o[1086]) );
  AND U29714 ( .A(p_input[11086]), .B(p_input[1086]), .Z(n19810) );
  AND U29715 ( .A(p_input[31086]), .B(p_input[21086]), .Z(n19809) );
  AND U29716 ( .A(n19811), .B(n19812), .Z(o[1085]) );
  AND U29717 ( .A(p_input[11085]), .B(p_input[1085]), .Z(n19812) );
  AND U29718 ( .A(p_input[31085]), .B(p_input[21085]), .Z(n19811) );
  AND U29719 ( .A(n19813), .B(n19814), .Z(o[1084]) );
  AND U29720 ( .A(p_input[11084]), .B(p_input[1084]), .Z(n19814) );
  AND U29721 ( .A(p_input[31084]), .B(p_input[21084]), .Z(n19813) );
  AND U29722 ( .A(n19815), .B(n19816), .Z(o[1083]) );
  AND U29723 ( .A(p_input[11083]), .B(p_input[1083]), .Z(n19816) );
  AND U29724 ( .A(p_input[31083]), .B(p_input[21083]), .Z(n19815) );
  AND U29725 ( .A(n19817), .B(n19818), .Z(o[1082]) );
  AND U29726 ( .A(p_input[11082]), .B(p_input[1082]), .Z(n19818) );
  AND U29727 ( .A(p_input[31082]), .B(p_input[21082]), .Z(n19817) );
  AND U29728 ( .A(n19819), .B(n19820), .Z(o[1081]) );
  AND U29729 ( .A(p_input[11081]), .B(p_input[1081]), .Z(n19820) );
  AND U29730 ( .A(p_input[31081]), .B(p_input[21081]), .Z(n19819) );
  AND U29731 ( .A(n19821), .B(n19822), .Z(o[1080]) );
  AND U29732 ( .A(p_input[11080]), .B(p_input[1080]), .Z(n19822) );
  AND U29733 ( .A(p_input[31080]), .B(p_input[21080]), .Z(n19821) );
  AND U29734 ( .A(n19823), .B(n19824), .Z(o[107]) );
  AND U29735 ( .A(p_input[107]), .B(p_input[10107]), .Z(n19824) );
  AND U29736 ( .A(p_input[30107]), .B(p_input[20107]), .Z(n19823) );
  AND U29737 ( .A(n19825), .B(n19826), .Z(o[1079]) );
  AND U29738 ( .A(p_input[11079]), .B(p_input[1079]), .Z(n19826) );
  AND U29739 ( .A(p_input[31079]), .B(p_input[21079]), .Z(n19825) );
  AND U29740 ( .A(n19827), .B(n19828), .Z(o[1078]) );
  AND U29741 ( .A(p_input[11078]), .B(p_input[1078]), .Z(n19828) );
  AND U29742 ( .A(p_input[31078]), .B(p_input[21078]), .Z(n19827) );
  AND U29743 ( .A(n19829), .B(n19830), .Z(o[1077]) );
  AND U29744 ( .A(p_input[11077]), .B(p_input[1077]), .Z(n19830) );
  AND U29745 ( .A(p_input[31077]), .B(p_input[21077]), .Z(n19829) );
  AND U29746 ( .A(n19831), .B(n19832), .Z(o[1076]) );
  AND U29747 ( .A(p_input[11076]), .B(p_input[1076]), .Z(n19832) );
  AND U29748 ( .A(p_input[31076]), .B(p_input[21076]), .Z(n19831) );
  AND U29749 ( .A(n19833), .B(n19834), .Z(o[1075]) );
  AND U29750 ( .A(p_input[11075]), .B(p_input[1075]), .Z(n19834) );
  AND U29751 ( .A(p_input[31075]), .B(p_input[21075]), .Z(n19833) );
  AND U29752 ( .A(n19835), .B(n19836), .Z(o[1074]) );
  AND U29753 ( .A(p_input[11074]), .B(p_input[1074]), .Z(n19836) );
  AND U29754 ( .A(p_input[31074]), .B(p_input[21074]), .Z(n19835) );
  AND U29755 ( .A(n19837), .B(n19838), .Z(o[1073]) );
  AND U29756 ( .A(p_input[11073]), .B(p_input[1073]), .Z(n19838) );
  AND U29757 ( .A(p_input[31073]), .B(p_input[21073]), .Z(n19837) );
  AND U29758 ( .A(n19839), .B(n19840), .Z(o[1072]) );
  AND U29759 ( .A(p_input[11072]), .B(p_input[1072]), .Z(n19840) );
  AND U29760 ( .A(p_input[31072]), .B(p_input[21072]), .Z(n19839) );
  AND U29761 ( .A(n19841), .B(n19842), .Z(o[1071]) );
  AND U29762 ( .A(p_input[11071]), .B(p_input[1071]), .Z(n19842) );
  AND U29763 ( .A(p_input[31071]), .B(p_input[21071]), .Z(n19841) );
  AND U29764 ( .A(n19843), .B(n19844), .Z(o[1070]) );
  AND U29765 ( .A(p_input[11070]), .B(p_input[1070]), .Z(n19844) );
  AND U29766 ( .A(p_input[31070]), .B(p_input[21070]), .Z(n19843) );
  AND U29767 ( .A(n19845), .B(n19846), .Z(o[106]) );
  AND U29768 ( .A(p_input[106]), .B(p_input[10106]), .Z(n19846) );
  AND U29769 ( .A(p_input[30106]), .B(p_input[20106]), .Z(n19845) );
  AND U29770 ( .A(n19847), .B(n19848), .Z(o[1069]) );
  AND U29771 ( .A(p_input[11069]), .B(p_input[1069]), .Z(n19848) );
  AND U29772 ( .A(p_input[31069]), .B(p_input[21069]), .Z(n19847) );
  AND U29773 ( .A(n19849), .B(n19850), .Z(o[1068]) );
  AND U29774 ( .A(p_input[11068]), .B(p_input[1068]), .Z(n19850) );
  AND U29775 ( .A(p_input[31068]), .B(p_input[21068]), .Z(n19849) );
  AND U29776 ( .A(n19851), .B(n19852), .Z(o[1067]) );
  AND U29777 ( .A(p_input[11067]), .B(p_input[1067]), .Z(n19852) );
  AND U29778 ( .A(p_input[31067]), .B(p_input[21067]), .Z(n19851) );
  AND U29779 ( .A(n19853), .B(n19854), .Z(o[1066]) );
  AND U29780 ( .A(p_input[11066]), .B(p_input[1066]), .Z(n19854) );
  AND U29781 ( .A(p_input[31066]), .B(p_input[21066]), .Z(n19853) );
  AND U29782 ( .A(n19855), .B(n19856), .Z(o[1065]) );
  AND U29783 ( .A(p_input[11065]), .B(p_input[1065]), .Z(n19856) );
  AND U29784 ( .A(p_input[31065]), .B(p_input[21065]), .Z(n19855) );
  AND U29785 ( .A(n19857), .B(n19858), .Z(o[1064]) );
  AND U29786 ( .A(p_input[11064]), .B(p_input[1064]), .Z(n19858) );
  AND U29787 ( .A(p_input[31064]), .B(p_input[21064]), .Z(n19857) );
  AND U29788 ( .A(n19859), .B(n19860), .Z(o[1063]) );
  AND U29789 ( .A(p_input[11063]), .B(p_input[1063]), .Z(n19860) );
  AND U29790 ( .A(p_input[31063]), .B(p_input[21063]), .Z(n19859) );
  AND U29791 ( .A(n19861), .B(n19862), .Z(o[1062]) );
  AND U29792 ( .A(p_input[11062]), .B(p_input[1062]), .Z(n19862) );
  AND U29793 ( .A(p_input[31062]), .B(p_input[21062]), .Z(n19861) );
  AND U29794 ( .A(n19863), .B(n19864), .Z(o[1061]) );
  AND U29795 ( .A(p_input[11061]), .B(p_input[1061]), .Z(n19864) );
  AND U29796 ( .A(p_input[31061]), .B(p_input[21061]), .Z(n19863) );
  AND U29797 ( .A(n19865), .B(n19866), .Z(o[1060]) );
  AND U29798 ( .A(p_input[11060]), .B(p_input[1060]), .Z(n19866) );
  AND U29799 ( .A(p_input[31060]), .B(p_input[21060]), .Z(n19865) );
  AND U29800 ( .A(n19867), .B(n19868), .Z(o[105]) );
  AND U29801 ( .A(p_input[105]), .B(p_input[10105]), .Z(n19868) );
  AND U29802 ( .A(p_input[30105]), .B(p_input[20105]), .Z(n19867) );
  AND U29803 ( .A(n19869), .B(n19870), .Z(o[1059]) );
  AND U29804 ( .A(p_input[11059]), .B(p_input[1059]), .Z(n19870) );
  AND U29805 ( .A(p_input[31059]), .B(p_input[21059]), .Z(n19869) );
  AND U29806 ( .A(n19871), .B(n19872), .Z(o[1058]) );
  AND U29807 ( .A(p_input[11058]), .B(p_input[1058]), .Z(n19872) );
  AND U29808 ( .A(p_input[31058]), .B(p_input[21058]), .Z(n19871) );
  AND U29809 ( .A(n19873), .B(n19874), .Z(o[1057]) );
  AND U29810 ( .A(p_input[11057]), .B(p_input[1057]), .Z(n19874) );
  AND U29811 ( .A(p_input[31057]), .B(p_input[21057]), .Z(n19873) );
  AND U29812 ( .A(n19875), .B(n19876), .Z(o[1056]) );
  AND U29813 ( .A(p_input[11056]), .B(p_input[1056]), .Z(n19876) );
  AND U29814 ( .A(p_input[31056]), .B(p_input[21056]), .Z(n19875) );
  AND U29815 ( .A(n19877), .B(n19878), .Z(o[1055]) );
  AND U29816 ( .A(p_input[11055]), .B(p_input[1055]), .Z(n19878) );
  AND U29817 ( .A(p_input[31055]), .B(p_input[21055]), .Z(n19877) );
  AND U29818 ( .A(n19879), .B(n19880), .Z(o[1054]) );
  AND U29819 ( .A(p_input[11054]), .B(p_input[1054]), .Z(n19880) );
  AND U29820 ( .A(p_input[31054]), .B(p_input[21054]), .Z(n19879) );
  AND U29821 ( .A(n19881), .B(n19882), .Z(o[1053]) );
  AND U29822 ( .A(p_input[11053]), .B(p_input[1053]), .Z(n19882) );
  AND U29823 ( .A(p_input[31053]), .B(p_input[21053]), .Z(n19881) );
  AND U29824 ( .A(n19883), .B(n19884), .Z(o[1052]) );
  AND U29825 ( .A(p_input[11052]), .B(p_input[1052]), .Z(n19884) );
  AND U29826 ( .A(p_input[31052]), .B(p_input[21052]), .Z(n19883) );
  AND U29827 ( .A(n19885), .B(n19886), .Z(o[1051]) );
  AND U29828 ( .A(p_input[11051]), .B(p_input[1051]), .Z(n19886) );
  AND U29829 ( .A(p_input[31051]), .B(p_input[21051]), .Z(n19885) );
  AND U29830 ( .A(n19887), .B(n19888), .Z(o[1050]) );
  AND U29831 ( .A(p_input[11050]), .B(p_input[1050]), .Z(n19888) );
  AND U29832 ( .A(p_input[31050]), .B(p_input[21050]), .Z(n19887) );
  AND U29833 ( .A(n19889), .B(n19890), .Z(o[104]) );
  AND U29834 ( .A(p_input[104]), .B(p_input[10104]), .Z(n19890) );
  AND U29835 ( .A(p_input[30104]), .B(p_input[20104]), .Z(n19889) );
  AND U29836 ( .A(n19891), .B(n19892), .Z(o[1049]) );
  AND U29837 ( .A(p_input[11049]), .B(p_input[1049]), .Z(n19892) );
  AND U29838 ( .A(p_input[31049]), .B(p_input[21049]), .Z(n19891) );
  AND U29839 ( .A(n19893), .B(n19894), .Z(o[1048]) );
  AND U29840 ( .A(p_input[11048]), .B(p_input[1048]), .Z(n19894) );
  AND U29841 ( .A(p_input[31048]), .B(p_input[21048]), .Z(n19893) );
  AND U29842 ( .A(n19895), .B(n19896), .Z(o[1047]) );
  AND U29843 ( .A(p_input[11047]), .B(p_input[1047]), .Z(n19896) );
  AND U29844 ( .A(p_input[31047]), .B(p_input[21047]), .Z(n19895) );
  AND U29845 ( .A(n19897), .B(n19898), .Z(o[1046]) );
  AND U29846 ( .A(p_input[11046]), .B(p_input[1046]), .Z(n19898) );
  AND U29847 ( .A(p_input[31046]), .B(p_input[21046]), .Z(n19897) );
  AND U29848 ( .A(n19899), .B(n19900), .Z(o[1045]) );
  AND U29849 ( .A(p_input[11045]), .B(p_input[1045]), .Z(n19900) );
  AND U29850 ( .A(p_input[31045]), .B(p_input[21045]), .Z(n19899) );
  AND U29851 ( .A(n19901), .B(n19902), .Z(o[1044]) );
  AND U29852 ( .A(p_input[11044]), .B(p_input[1044]), .Z(n19902) );
  AND U29853 ( .A(p_input[31044]), .B(p_input[21044]), .Z(n19901) );
  AND U29854 ( .A(n19903), .B(n19904), .Z(o[1043]) );
  AND U29855 ( .A(p_input[11043]), .B(p_input[1043]), .Z(n19904) );
  AND U29856 ( .A(p_input[31043]), .B(p_input[21043]), .Z(n19903) );
  AND U29857 ( .A(n19905), .B(n19906), .Z(o[1042]) );
  AND U29858 ( .A(p_input[11042]), .B(p_input[1042]), .Z(n19906) );
  AND U29859 ( .A(p_input[31042]), .B(p_input[21042]), .Z(n19905) );
  AND U29860 ( .A(n19907), .B(n19908), .Z(o[1041]) );
  AND U29861 ( .A(p_input[11041]), .B(p_input[1041]), .Z(n19908) );
  AND U29862 ( .A(p_input[31041]), .B(p_input[21041]), .Z(n19907) );
  AND U29863 ( .A(n19909), .B(n19910), .Z(o[1040]) );
  AND U29864 ( .A(p_input[11040]), .B(p_input[1040]), .Z(n19910) );
  AND U29865 ( .A(p_input[31040]), .B(p_input[21040]), .Z(n19909) );
  AND U29866 ( .A(n19911), .B(n19912), .Z(o[103]) );
  AND U29867 ( .A(p_input[103]), .B(p_input[10103]), .Z(n19912) );
  AND U29868 ( .A(p_input[30103]), .B(p_input[20103]), .Z(n19911) );
  AND U29869 ( .A(n19913), .B(n19914), .Z(o[1039]) );
  AND U29870 ( .A(p_input[11039]), .B(p_input[1039]), .Z(n19914) );
  AND U29871 ( .A(p_input[31039]), .B(p_input[21039]), .Z(n19913) );
  AND U29872 ( .A(n19915), .B(n19916), .Z(o[1038]) );
  AND U29873 ( .A(p_input[11038]), .B(p_input[1038]), .Z(n19916) );
  AND U29874 ( .A(p_input[31038]), .B(p_input[21038]), .Z(n19915) );
  AND U29875 ( .A(n19917), .B(n19918), .Z(o[1037]) );
  AND U29876 ( .A(p_input[11037]), .B(p_input[1037]), .Z(n19918) );
  AND U29877 ( .A(p_input[31037]), .B(p_input[21037]), .Z(n19917) );
  AND U29878 ( .A(n19919), .B(n19920), .Z(o[1036]) );
  AND U29879 ( .A(p_input[11036]), .B(p_input[1036]), .Z(n19920) );
  AND U29880 ( .A(p_input[31036]), .B(p_input[21036]), .Z(n19919) );
  AND U29881 ( .A(n19921), .B(n19922), .Z(o[1035]) );
  AND U29882 ( .A(p_input[11035]), .B(p_input[1035]), .Z(n19922) );
  AND U29883 ( .A(p_input[31035]), .B(p_input[21035]), .Z(n19921) );
  AND U29884 ( .A(n19923), .B(n19924), .Z(o[1034]) );
  AND U29885 ( .A(p_input[11034]), .B(p_input[1034]), .Z(n19924) );
  AND U29886 ( .A(p_input[31034]), .B(p_input[21034]), .Z(n19923) );
  AND U29887 ( .A(n19925), .B(n19926), .Z(o[1033]) );
  AND U29888 ( .A(p_input[11033]), .B(p_input[1033]), .Z(n19926) );
  AND U29889 ( .A(p_input[31033]), .B(p_input[21033]), .Z(n19925) );
  AND U29890 ( .A(n19927), .B(n19928), .Z(o[1032]) );
  AND U29891 ( .A(p_input[11032]), .B(p_input[1032]), .Z(n19928) );
  AND U29892 ( .A(p_input[31032]), .B(p_input[21032]), .Z(n19927) );
  AND U29893 ( .A(n19929), .B(n19930), .Z(o[1031]) );
  AND U29894 ( .A(p_input[11031]), .B(p_input[1031]), .Z(n19930) );
  AND U29895 ( .A(p_input[31031]), .B(p_input[21031]), .Z(n19929) );
  AND U29896 ( .A(n19931), .B(n19932), .Z(o[1030]) );
  AND U29897 ( .A(p_input[11030]), .B(p_input[1030]), .Z(n19932) );
  AND U29898 ( .A(p_input[31030]), .B(p_input[21030]), .Z(n19931) );
  AND U29899 ( .A(n19933), .B(n19934), .Z(o[102]) );
  AND U29900 ( .A(p_input[102]), .B(p_input[10102]), .Z(n19934) );
  AND U29901 ( .A(p_input[30102]), .B(p_input[20102]), .Z(n19933) );
  AND U29902 ( .A(n19935), .B(n19936), .Z(o[1029]) );
  AND U29903 ( .A(p_input[11029]), .B(p_input[1029]), .Z(n19936) );
  AND U29904 ( .A(p_input[31029]), .B(p_input[21029]), .Z(n19935) );
  AND U29905 ( .A(n19937), .B(n19938), .Z(o[1028]) );
  AND U29906 ( .A(p_input[11028]), .B(p_input[1028]), .Z(n19938) );
  AND U29907 ( .A(p_input[31028]), .B(p_input[21028]), .Z(n19937) );
  AND U29908 ( .A(n19939), .B(n19940), .Z(o[1027]) );
  AND U29909 ( .A(p_input[11027]), .B(p_input[1027]), .Z(n19940) );
  AND U29910 ( .A(p_input[31027]), .B(p_input[21027]), .Z(n19939) );
  AND U29911 ( .A(n19941), .B(n19942), .Z(o[1026]) );
  AND U29912 ( .A(p_input[11026]), .B(p_input[1026]), .Z(n19942) );
  AND U29913 ( .A(p_input[31026]), .B(p_input[21026]), .Z(n19941) );
  AND U29914 ( .A(n19943), .B(n19944), .Z(o[1025]) );
  AND U29915 ( .A(p_input[11025]), .B(p_input[1025]), .Z(n19944) );
  AND U29916 ( .A(p_input[31025]), .B(p_input[21025]), .Z(n19943) );
  AND U29917 ( .A(n19945), .B(n19946), .Z(o[1024]) );
  AND U29918 ( .A(p_input[11024]), .B(p_input[1024]), .Z(n19946) );
  AND U29919 ( .A(p_input[31024]), .B(p_input[21024]), .Z(n19945) );
  AND U29920 ( .A(n19947), .B(n19948), .Z(o[1023]) );
  AND U29921 ( .A(p_input[11023]), .B(p_input[1023]), .Z(n19948) );
  AND U29922 ( .A(p_input[31023]), .B(p_input[21023]), .Z(n19947) );
  AND U29923 ( .A(n19949), .B(n19950), .Z(o[1022]) );
  AND U29924 ( .A(p_input[11022]), .B(p_input[1022]), .Z(n19950) );
  AND U29925 ( .A(p_input[31022]), .B(p_input[21022]), .Z(n19949) );
  AND U29926 ( .A(n19951), .B(n19952), .Z(o[1021]) );
  AND U29927 ( .A(p_input[11021]), .B(p_input[1021]), .Z(n19952) );
  AND U29928 ( .A(p_input[31021]), .B(p_input[21021]), .Z(n19951) );
  AND U29929 ( .A(n19953), .B(n19954), .Z(o[1020]) );
  AND U29930 ( .A(p_input[11020]), .B(p_input[1020]), .Z(n19954) );
  AND U29931 ( .A(p_input[31020]), .B(p_input[21020]), .Z(n19953) );
  AND U29932 ( .A(n19955), .B(n19956), .Z(o[101]) );
  AND U29933 ( .A(p_input[101]), .B(p_input[10101]), .Z(n19956) );
  AND U29934 ( .A(p_input[30101]), .B(p_input[20101]), .Z(n19955) );
  AND U29935 ( .A(n19957), .B(n19958), .Z(o[1019]) );
  AND U29936 ( .A(p_input[11019]), .B(p_input[1019]), .Z(n19958) );
  AND U29937 ( .A(p_input[31019]), .B(p_input[21019]), .Z(n19957) );
  AND U29938 ( .A(n19959), .B(n19960), .Z(o[1018]) );
  AND U29939 ( .A(p_input[11018]), .B(p_input[1018]), .Z(n19960) );
  AND U29940 ( .A(p_input[31018]), .B(p_input[21018]), .Z(n19959) );
  AND U29941 ( .A(n19961), .B(n19962), .Z(o[1017]) );
  AND U29942 ( .A(p_input[11017]), .B(p_input[1017]), .Z(n19962) );
  AND U29943 ( .A(p_input[31017]), .B(p_input[21017]), .Z(n19961) );
  AND U29944 ( .A(n19963), .B(n19964), .Z(o[1016]) );
  AND U29945 ( .A(p_input[11016]), .B(p_input[1016]), .Z(n19964) );
  AND U29946 ( .A(p_input[31016]), .B(p_input[21016]), .Z(n19963) );
  AND U29947 ( .A(n19965), .B(n19966), .Z(o[1015]) );
  AND U29948 ( .A(p_input[11015]), .B(p_input[1015]), .Z(n19966) );
  AND U29949 ( .A(p_input[31015]), .B(p_input[21015]), .Z(n19965) );
  AND U29950 ( .A(n19967), .B(n19968), .Z(o[1014]) );
  AND U29951 ( .A(p_input[11014]), .B(p_input[1014]), .Z(n19968) );
  AND U29952 ( .A(p_input[31014]), .B(p_input[21014]), .Z(n19967) );
  AND U29953 ( .A(n19969), .B(n19970), .Z(o[1013]) );
  AND U29954 ( .A(p_input[11013]), .B(p_input[1013]), .Z(n19970) );
  AND U29955 ( .A(p_input[31013]), .B(p_input[21013]), .Z(n19969) );
  AND U29956 ( .A(n19971), .B(n19972), .Z(o[1012]) );
  AND U29957 ( .A(p_input[11012]), .B(p_input[1012]), .Z(n19972) );
  AND U29958 ( .A(p_input[31012]), .B(p_input[21012]), .Z(n19971) );
  AND U29959 ( .A(n19973), .B(n19974), .Z(o[1011]) );
  AND U29960 ( .A(p_input[11011]), .B(p_input[1011]), .Z(n19974) );
  AND U29961 ( .A(p_input[31011]), .B(p_input[21011]), .Z(n19973) );
  AND U29962 ( .A(n19975), .B(n19976), .Z(o[1010]) );
  AND U29963 ( .A(p_input[11010]), .B(p_input[1010]), .Z(n19976) );
  AND U29964 ( .A(p_input[31010]), .B(p_input[21010]), .Z(n19975) );
  AND U29965 ( .A(n19977), .B(n19978), .Z(o[100]) );
  AND U29966 ( .A(p_input[10100]), .B(p_input[100]), .Z(n19978) );
  AND U29967 ( .A(p_input[30100]), .B(p_input[20100]), .Z(n19977) );
  AND U29968 ( .A(n19979), .B(n19980), .Z(o[1009]) );
  AND U29969 ( .A(p_input[11009]), .B(p_input[1009]), .Z(n19980) );
  AND U29970 ( .A(p_input[31009]), .B(p_input[21009]), .Z(n19979) );
  AND U29971 ( .A(n19981), .B(n19982), .Z(o[1008]) );
  AND U29972 ( .A(p_input[11008]), .B(p_input[1008]), .Z(n19982) );
  AND U29973 ( .A(p_input[31008]), .B(p_input[21008]), .Z(n19981) );
  AND U29974 ( .A(n19983), .B(n19984), .Z(o[1007]) );
  AND U29975 ( .A(p_input[11007]), .B(p_input[1007]), .Z(n19984) );
  AND U29976 ( .A(p_input[31007]), .B(p_input[21007]), .Z(n19983) );
  AND U29977 ( .A(n19985), .B(n19986), .Z(o[1006]) );
  AND U29978 ( .A(p_input[11006]), .B(p_input[1006]), .Z(n19986) );
  AND U29979 ( .A(p_input[31006]), .B(p_input[21006]), .Z(n19985) );
  AND U29980 ( .A(n19987), .B(n19988), .Z(o[1005]) );
  AND U29981 ( .A(p_input[11005]), .B(p_input[1005]), .Z(n19988) );
  AND U29982 ( .A(p_input[31005]), .B(p_input[21005]), .Z(n19987) );
  AND U29983 ( .A(n19989), .B(n19990), .Z(o[1004]) );
  AND U29984 ( .A(p_input[11004]), .B(p_input[1004]), .Z(n19990) );
  AND U29985 ( .A(p_input[31004]), .B(p_input[21004]), .Z(n19989) );
  AND U29986 ( .A(n19991), .B(n19992), .Z(o[1003]) );
  AND U29987 ( .A(p_input[11003]), .B(p_input[1003]), .Z(n19992) );
  AND U29988 ( .A(p_input[31003]), .B(p_input[21003]), .Z(n19991) );
  AND U29989 ( .A(n19993), .B(n19994), .Z(o[1002]) );
  AND U29990 ( .A(p_input[11002]), .B(p_input[1002]), .Z(n19994) );
  AND U29991 ( .A(p_input[31002]), .B(p_input[21002]), .Z(n19993) );
  AND U29992 ( .A(n19995), .B(n19996), .Z(o[1001]) );
  AND U29993 ( .A(p_input[11001]), .B(p_input[1001]), .Z(n19996) );
  AND U29994 ( .A(p_input[31001]), .B(p_input[21001]), .Z(n19995) );
  AND U29995 ( .A(n19997), .B(n19998), .Z(o[1000]) );
  AND U29996 ( .A(p_input[11000]), .B(p_input[1000]), .Z(n19998) );
  AND U29997 ( .A(p_input[31000]), .B(p_input[21000]), .Z(n19997) );
  AND U29998 ( .A(n19999), .B(n20000), .Z(o[0]) );
  AND U29999 ( .A(p_input[10000]), .B(p_input[0]), .Z(n20000) );
  AND U30000 ( .A(p_input[30000]), .B(p_input[20000]), .Z(n19999) );
endmodule

