
module auction_BMR_N7_W16 ( p_input, o );
  input [2047:0] p_input;
  output [22:0] o;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972,
         n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982,
         n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992,
         n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002,
         n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
         n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022,
         n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032,
         n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042,
         n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052,
         n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062,
         n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072,
         n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082,
         n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092,
         n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102,
         n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112,
         n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122,
         n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132,
         n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142,
         n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152,
         n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162,
         n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172,
         n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182,
         n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192,
         n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202,
         n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212,
         n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222,
         n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232,
         n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242,
         n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252,
         n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262,
         n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272,
         n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282,
         n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292,
         n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302,
         n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312,
         n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322,
         n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332,
         n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342,
         n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352,
         n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362,
         n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372,
         n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382,
         n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392,
         n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402,
         n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412,
         n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422,
         n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432,
         n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442,
         n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452,
         n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
         n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
         n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
         n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
         n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
         n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612,
         n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622,
         n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632,
         n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
         n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652,
         n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662,
         n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672,
         n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682,
         n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692,
         n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702,
         n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712,
         n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722,
         n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732,
         n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742,
         n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752,
         n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762,
         n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772,
         n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782,
         n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792,
         n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802,
         n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812,
         n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822,
         n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832,
         n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842,
         n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852,
         n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862,
         n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872,
         n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882,
         n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892,
         n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902,
         n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912,
         n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922,
         n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932,
         n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942,
         n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952,
         n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962,
         n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972,
         n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982,
         n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992,
         n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002,
         n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012,
         n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022,
         n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032,
         n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042,
         n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052,
         n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062,
         n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072,
         n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082,
         n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092,
         n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102,
         n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112,
         n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122,
         n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132,
         n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142,
         n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152,
         n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162,
         n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172,
         n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182,
         n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192,
         n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202,
         n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212,
         n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222,
         n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232,
         n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242,
         n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252,
         n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262,
         n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272,
         n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282,
         n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292,
         n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302,
         n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312,
         n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322,
         n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332,
         n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342,
         n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352,
         n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362,
         n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372,
         n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382,
         n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392,
         n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402,
         n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412,
         n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422,
         n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432,
         n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442,
         n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452,
         n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462,
         n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472,
         n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482,
         n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492,
         n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502,
         n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512,
         n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522,
         n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532,
         n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542,
         n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552,
         n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562,
         n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572,
         n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582,
         n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592,
         n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602,
         n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612,
         n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622,
         n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632,
         n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642,
         n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652,
         n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662,
         n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672,
         n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682,
         n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692,
         n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702,
         n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712,
         n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722,
         n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732,
         n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742,
         n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752,
         n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762,
         n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772,
         n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782,
         n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792,
         n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802,
         n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812,
         n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822,
         n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832,
         n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842,
         n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852,
         n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862,
         n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872,
         n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882,
         n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892,
         n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902,
         n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912,
         n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922,
         n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932,
         n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942,
         n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952,
         n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962,
         n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972,
         n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982,
         n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992,
         n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002,
         n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012,
         n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022,
         n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032,
         n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042,
         n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052,
         n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062,
         n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072,
         n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082,
         n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092,
         n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102,
         n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112,
         n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122,
         n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132,
         n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142,
         n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152,
         n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162,
         n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172,
         n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182,
         n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192,
         n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202,
         n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212,
         n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222,
         n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232,
         n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242,
         n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252,
         n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262,
         n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272,
         n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282,
         n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292,
         n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302,
         n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312,
         n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322,
         n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332,
         n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342,
         n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352,
         n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362,
         n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372,
         n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382,
         n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392,
         n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402,
         n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412,
         n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422,
         n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432,
         n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442,
         n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452,
         n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462,
         n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472,
         n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482,
         n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492,
         n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502,
         n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512,
         n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522,
         n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532,
         n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542,
         n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552,
         n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562,
         n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572,
         n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582,
         n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592,
         n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602,
         n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612,
         n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622,
         n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632,
         n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642,
         n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652,
         n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662,
         n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672,
         n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682,
         n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692,
         n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702,
         n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712,
         n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722,
         n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732,
         n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742,
         n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752,
         n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762,
         n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772,
         n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782,
         n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792,
         n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802,
         n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812,
         n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822,
         n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832,
         n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842,
         n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852,
         n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862,
         n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872,
         n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882,
         n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892,
         n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902,
         n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912,
         n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922,
         n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932,
         n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942,
         n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952,
         n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962,
         n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972,
         n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982,
         n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992,
         n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002,
         n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012,
         n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022,
         n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032,
         n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042,
         n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052,
         n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062,
         n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072,
         n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082,
         n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092,
         n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102,
         n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112,
         n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122,
         n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132,
         n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142,
         n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152,
         n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162,
         n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172,
         n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182,
         n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192,
         n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202,
         n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212,
         n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222,
         n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232,
         n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242,
         n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252,
         n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262,
         n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272,
         n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282,
         n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292,
         n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302,
         n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312,
         n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322,
         n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332,
         n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342,
         n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352,
         n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362,
         n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372,
         n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382,
         n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392,
         n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402,
         n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412,
         n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422,
         n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432,
         n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442,
         n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452,
         n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462,
         n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472,
         n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482,
         n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492,
         n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502,
         n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512,
         n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522,
         n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532,
         n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542,
         n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552,
         n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562,
         n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572,
         n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582,
         n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592,
         n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602,
         n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612,
         n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622,
         n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632,
         n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642,
         n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652,
         n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662,
         n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672,
         n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682,
         n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692,
         n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702,
         n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712,
         n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722,
         n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732,
         n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742,
         n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752,
         n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762,
         n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772,
         n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782,
         n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792,
         n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802,
         n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812,
         n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822,
         n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832,
         n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842,
         n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852,
         n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862,
         n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872,
         n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882,
         n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892,
         n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902,
         n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912,
         n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922,
         n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932,
         n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942,
         n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952,
         n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962,
         n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972,
         n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982,
         n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992,
         n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002,
         n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012,
         n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022,
         n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032,
         n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042,
         n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052,
         n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062,
         n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072,
         n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082,
         n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092,
         n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102,
         n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112,
         n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122,
         n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132,
         n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142,
         n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152,
         n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162,
         n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172,
         n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182,
         n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192,
         n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202,
         n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212,
         n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222,
         n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232,
         n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242,
         n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252,
         n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262,
         n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272,
         n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282,
         n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292,
         n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302,
         n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312,
         n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322,
         n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332,
         n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342,
         n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352,
         n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362,
         n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372,
         n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382,
         n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392,
         n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402,
         n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412,
         n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422,
         n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432,
         n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442,
         n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452,
         n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462,
         n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472,
         n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482,
         n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492,
         n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502,
         n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512,
         n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522,
         n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532,
         n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542,
         n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552,
         n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562,
         n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572,
         n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582,
         n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592,
         n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602,
         n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612,
         n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622,
         n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632,
         n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642,
         n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652,
         n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662,
         n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672,
         n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682,
         n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692,
         n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702,
         n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712,
         n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722,
         n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732,
         n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742,
         n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752,
         n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762,
         n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772,
         n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782,
         n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792,
         n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802,
         n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812,
         n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822,
         n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832,
         n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842,
         n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852,
         n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862,
         n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872,
         n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882,
         n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892,
         n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902,
         n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912,
         n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922,
         n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932,
         n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942,
         n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952,
         n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962,
         n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972,
         n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982,
         n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992,
         n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002,
         n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012,
         n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022,
         n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032,
         n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042,
         n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052,
         n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062,
         n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072,
         n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082,
         n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092,
         n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102,
         n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112,
         n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122,
         n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132,
         n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142,
         n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152,
         n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162,
         n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172,
         n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182,
         n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192,
         n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202,
         n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212,
         n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222,
         n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232,
         n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242,
         n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252,
         n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262,
         n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272,
         n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282,
         n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292,
         n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302,
         n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312,
         n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322,
         n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332,
         n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342,
         n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352,
         n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362,
         n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372,
         n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382,
         n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392,
         n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402,
         n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412,
         n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422,
         n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432,
         n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442,
         n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452,
         n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462,
         n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472,
         n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482,
         n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492,
         n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502,
         n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512,
         n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522,
         n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532,
         n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542,
         n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552,
         n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562,
         n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572,
         n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582,
         n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592,
         n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602,
         n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612,
         n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622,
         n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632,
         n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642,
         n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652,
         n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662,
         n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672,
         n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682,
         n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692,
         n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702,
         n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712,
         n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722,
         n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732,
         n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742,
         n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752,
         n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762,
         n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772,
         n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782,
         n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792,
         n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802,
         n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812,
         n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822,
         n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832,
         n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842,
         n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852,
         n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862,
         n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872,
         n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882,
         n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892,
         n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902,
         n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912,
         n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922,
         n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932,
         n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942,
         n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952,
         n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962,
         n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972,
         n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982,
         n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992,
         n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001,
         n10002, n10003, n10004, n10005, n10006, n10007, n10008, n10009,
         n10010, n10011, n10012, n10013, n10014, n10015, n10016, n10017,
         n10018, n10019, n10020, n10021, n10022, n10023, n10024, n10025,
         n10026, n10027, n10028, n10029, n10030, n10031, n10032, n10033,
         n10034, n10035, n10036, n10037, n10038, n10039, n10040, n10041,
         n10042, n10043, n10044, n10045, n10046, n10047, n10048, n10049,
         n10050, n10051, n10052, n10053, n10054, n10055, n10056, n10057,
         n10058, n10059, n10060, n10061, n10062, n10063, n10064, n10065,
         n10066, n10067, n10068, n10069, n10070, n10071, n10072, n10073,
         n10074, n10075, n10076, n10077, n10078, n10079, n10080, n10081,
         n10082, n10083, n10084, n10085, n10086, n10087, n10088, n10089,
         n10090, n10091, n10092, n10093, n10094, n10095, n10096, n10097,
         n10098, n10099, n10100, n10101, n10102, n10103, n10104, n10105,
         n10106, n10107, n10108, n10109, n10110, n10111, n10112, n10113,
         n10114, n10115, n10116, n10117, n10118, n10119, n10120, n10121,
         n10122, n10123, n10124, n10125, n10126, n10127, n10128, n10129,
         n10130, n10131, n10132, n10133, n10134, n10135, n10136, n10137,
         n10138, n10139, n10140, n10141, n10142, n10143, n10144, n10145,
         n10146, n10147, n10148, n10149, n10150, n10151, n10152, n10153,
         n10154, n10155, n10156, n10157, n10158, n10159, n10160, n10161,
         n10162, n10163, n10164, n10165, n10166, n10167, n10168, n10169,
         n10170, n10171, n10172, n10173, n10174, n10175, n10176, n10177,
         n10178, n10179, n10180, n10181, n10182, n10183, n10184, n10185,
         n10186, n10187, n10188, n10189, n10190, n10191, n10192, n10193,
         n10194, n10195, n10196, n10197, n10198, n10199, n10200, n10201,
         n10202, n10203, n10204, n10205, n10206, n10207, n10208, n10209,
         n10210, n10211, n10212, n10213, n10214, n10215, n10216, n10217,
         n10218, n10219, n10220, n10221, n10222, n10223, n10224, n10225,
         n10226, n10227, n10228, n10229, n10230, n10231, n10232, n10233,
         n10234, n10235, n10236, n10237, n10238, n10239, n10240, n10241,
         n10242, n10243, n10244, n10245, n10246, n10247, n10248, n10249,
         n10250, n10251, n10252, n10253, n10254, n10255, n10256, n10257,
         n10258, n10259, n10260, n10261, n10262, n10263, n10264, n10265,
         n10266, n10267, n10268, n10269, n10270, n10271, n10272, n10273,
         n10274, n10275, n10276, n10277, n10278, n10279, n10280, n10281,
         n10282, n10283, n10284, n10285, n10286, n10287, n10288, n10289,
         n10290, n10291, n10292, n10293, n10294, n10295, n10296, n10297,
         n10298, n10299, n10300, n10301, n10302, n10303, n10304, n10305,
         n10306, n10307, n10308, n10309, n10310, n10311, n10312, n10313,
         n10314, n10315, n10316, n10317, n10318, n10319, n10320, n10321,
         n10322, n10323, n10324, n10325, n10326, n10327, n10328, n10329,
         n10330, n10331, n10332, n10333, n10334, n10335, n10336, n10337,
         n10338, n10339, n10340, n10341, n10342, n10343, n10344, n10345,
         n10346, n10347, n10348, n10349, n10350, n10351, n10352, n10353,
         n10354, n10355, n10356, n10357, n10358, n10359, n10360, n10361,
         n10362, n10363, n10364, n10365, n10366, n10367, n10368, n10369,
         n10370, n10371, n10372, n10373, n10374, n10375, n10376, n10377,
         n10378, n10379, n10380, n10381, n10382, n10383, n10384, n10385,
         n10386, n10387, n10388, n10389, n10390, n10391, n10392, n10393,
         n10394, n10395, n10396, n10397, n10398, n10399, n10400, n10401,
         n10402, n10403, n10404, n10405, n10406, n10407, n10408, n10409,
         n10410, n10411, n10412, n10413, n10414, n10415, n10416, n10417,
         n10418, n10419, n10420, n10421, n10422, n10423, n10424, n10425,
         n10426, n10427, n10428, n10429, n10430, n10431, n10432, n10433,
         n10434, n10435, n10436, n10437, n10438, n10439, n10440, n10441,
         n10442, n10443, n10444, n10445, n10446, n10447, n10448, n10449,
         n10450, n10451, n10452, n10453, n10454, n10455, n10456, n10457,
         n10458, n10459, n10460, n10461, n10462, n10463, n10464, n10465,
         n10466, n10467, n10468, n10469, n10470, n10471, n10472, n10473,
         n10474, n10475, n10476, n10477, n10478, n10479, n10480, n10481,
         n10482, n10483, n10484, n10485, n10486, n10487, n10488, n10489,
         n10490, n10491, n10492, n10493, n10494, n10495, n10496, n10497,
         n10498, n10499, n10500, n10501, n10502, n10503, n10504, n10505,
         n10506, n10507, n10508, n10509, n10510, n10511, n10512, n10513,
         n10514, n10515, n10516, n10517, n10518, n10519, n10520, n10521,
         n10522, n10523, n10524, n10525, n10526, n10527, n10528, n10529,
         n10530, n10531, n10532, n10533, n10534, n10535, n10536, n10537,
         n10538, n10539, n10540, n10541, n10542, n10543, n10544, n10545,
         n10546, n10547, n10548, n10549, n10550, n10551, n10552, n10553,
         n10554, n10555, n10556, n10557, n10558, n10559, n10560, n10561,
         n10562, n10563, n10564, n10565, n10566, n10567, n10568, n10569,
         n10570, n10571, n10572, n10573, n10574, n10575, n10576, n10577,
         n10578, n10579, n10580, n10581, n10582, n10583, n10584, n10585,
         n10586, n10587, n10588, n10589, n10590, n10591, n10592, n10593,
         n10594, n10595, n10596, n10597, n10598, n10599, n10600, n10601,
         n10602, n10603, n10604, n10605, n10606, n10607, n10608, n10609,
         n10610, n10611, n10612, n10613, n10614, n10615, n10616, n10617,
         n10618, n10619, n10620, n10621, n10622, n10623, n10624, n10625,
         n10626, n10627, n10628, n10629, n10630, n10631, n10632, n10633,
         n10634, n10635, n10636, n10637, n10638, n10639, n10640, n10641,
         n10642, n10643, n10644, n10645, n10646, n10647, n10648, n10649,
         n10650, n10651, n10652, n10653, n10654, n10655, n10656, n10657,
         n10658, n10659, n10660, n10661, n10662, n10663, n10664, n10665,
         n10666, n10667, n10668, n10669, n10670, n10671, n10672, n10673,
         n10674, n10675, n10676, n10677, n10678, n10679, n10680, n10681,
         n10682, n10683, n10684, n10685, n10686, n10687, n10688, n10689,
         n10690, n10691, n10692, n10693, n10694, n10695, n10696, n10697,
         n10698, n10699, n10700, n10701, n10702, n10703, n10704, n10705,
         n10706, n10707, n10708, n10709, n10710, n10711, n10712, n10713,
         n10714, n10715, n10716, n10717, n10718, n10719, n10720, n10721,
         n10722, n10723, n10724, n10725, n10726, n10727, n10728, n10729,
         n10730, n10731, n10732, n10733, n10734, n10735, n10736, n10737,
         n10738, n10739, n10740, n10741, n10742, n10743, n10744, n10745,
         n10746, n10747, n10748, n10749, n10750, n10751, n10752, n10753,
         n10754, n10755, n10756, n10757, n10758, n10759, n10760, n10761,
         n10762, n10763, n10764, n10765, n10766, n10767, n10768, n10769,
         n10770, n10771, n10772, n10773, n10774, n10775, n10776, n10777,
         n10778, n10779, n10780, n10781, n10782, n10783, n10784, n10785,
         n10786, n10787, n10788, n10789, n10790, n10791, n10792, n10793,
         n10794, n10795, n10796, n10797, n10798, n10799, n10800, n10801,
         n10802, n10803, n10804, n10805, n10806, n10807, n10808, n10809,
         n10810, n10811, n10812, n10813, n10814, n10815, n10816, n10817,
         n10818, n10819, n10820, n10821, n10822, n10823, n10824, n10825,
         n10826, n10827, n10828, n10829, n10830, n10831, n10832, n10833,
         n10834, n10835, n10836, n10837, n10838, n10839, n10840, n10841,
         n10842, n10843, n10844, n10845, n10846, n10847, n10848, n10849,
         n10850, n10851, n10852, n10853, n10854, n10855, n10856, n10857,
         n10858, n10859, n10860, n10861, n10862, n10863, n10864, n10865,
         n10866, n10867, n10868, n10869, n10870, n10871, n10872, n10873,
         n10874, n10875, n10876, n10877, n10878, n10879, n10880, n10881,
         n10882, n10883, n10884, n10885, n10886, n10887, n10888, n10889,
         n10890, n10891, n10892, n10893, n10894, n10895, n10896, n10897,
         n10898, n10899, n10900, n10901, n10902, n10903, n10904, n10905,
         n10906, n10907, n10908, n10909, n10910, n10911, n10912, n10913,
         n10914, n10915, n10916, n10917, n10918, n10919, n10920, n10921,
         n10922, n10923, n10924, n10925, n10926, n10927, n10928, n10929,
         n10930, n10931, n10932, n10933, n10934, n10935, n10936, n10937,
         n10938, n10939, n10940, n10941, n10942, n10943, n10944, n10945,
         n10946, n10947, n10948, n10949, n10950, n10951, n10952, n10953,
         n10954, n10955, n10956, n10957, n10958, n10959, n10960, n10961,
         n10962, n10963, n10964, n10965, n10966, n10967, n10968, n10969,
         n10970, n10971, n10972, n10973, n10974, n10975, n10976, n10977,
         n10978, n10979, n10980, n10981, n10982, n10983, n10984, n10985,
         n10986, n10987, n10988, n10989, n10990, n10991, n10992, n10993,
         n10994, n10995, n10996, n10997, n10998, n10999, n11000, n11001,
         n11002, n11003, n11004, n11005, n11006, n11007, n11008, n11009,
         n11010, n11011, n11012, n11013, n11014, n11015, n11016, n11017,
         n11018, n11019, n11020, n11021, n11022, n11023, n11024, n11025,
         n11026, n11027, n11028, n11029, n11030, n11031, n11032, n11033,
         n11034, n11035, n11036, n11037, n11038, n11039, n11040, n11041,
         n11042, n11043, n11044, n11045, n11046, n11047, n11048, n11049,
         n11050, n11051, n11052, n11053, n11054, n11055, n11056, n11057,
         n11058, n11059, n11060, n11061, n11062, n11063, n11064, n11065,
         n11066, n11067, n11068, n11069, n11070, n11071, n11072, n11073,
         n11074, n11075, n11076, n11077, n11078, n11079, n11080, n11081,
         n11082, n11083, n11084, n11085, n11086, n11087, n11088, n11089,
         n11090, n11091, n11092, n11093, n11094, n11095, n11096, n11097,
         n11098, n11099, n11100, n11101, n11102, n11103, n11104, n11105,
         n11106, n11107, n11108, n11109, n11110, n11111, n11112, n11113,
         n11114, n11115, n11116, n11117, n11118, n11119, n11120, n11121,
         n11122, n11123, n11124, n11125, n11126, n11127, n11128, n11129,
         n11130, n11131, n11132, n11133, n11134, n11135, n11136, n11137,
         n11138, n11139, n11140, n11141, n11142, n11143, n11144, n11145,
         n11146, n11147, n11148, n11149, n11150, n11151, n11152, n11153,
         n11154, n11155, n11156, n11157, n11158, n11159, n11160, n11161,
         n11162, n11163, n11164, n11165, n11166, n11167, n11168, n11169,
         n11170, n11171, n11172, n11173, n11174, n11175, n11176, n11177,
         n11178, n11179, n11180, n11181, n11182, n11183, n11184, n11185,
         n11186, n11187, n11188, n11189, n11190, n11191, n11192, n11193,
         n11194, n11195, n11196, n11197, n11198, n11199, n11200, n11201,
         n11202, n11203, n11204, n11205, n11206, n11207, n11208, n11209,
         n11210, n11211, n11212, n11213, n11214, n11215, n11216, n11217,
         n11218, n11219, n11220, n11221, n11222, n11223, n11224, n11225,
         n11226, n11227, n11228, n11229, n11230, n11231, n11232, n11233,
         n11234, n11235, n11236, n11237, n11238, n11239, n11240, n11241,
         n11242, n11243, n11244, n11245, n11246, n11247, n11248, n11249,
         n11250, n11251, n11252, n11253, n11254, n11255, n11256, n11257,
         n11258, n11259, n11260, n11261, n11262, n11263, n11264, n11265,
         n11266, n11267, n11268, n11269, n11270, n11271, n11272, n11273,
         n11274, n11275, n11276, n11277, n11278, n11279, n11280, n11281,
         n11282, n11283, n11284, n11285, n11286, n11287, n11288, n11289,
         n11290, n11291, n11292, n11293, n11294, n11295, n11296, n11297,
         n11298, n11299, n11300, n11301, n11302, n11303, n11304, n11305,
         n11306, n11307, n11308, n11309, n11310, n11311, n11312, n11313,
         n11314, n11315, n11316, n11317, n11318, n11319, n11320, n11321,
         n11322, n11323, n11324, n11325, n11326, n11327, n11328, n11329,
         n11330, n11331, n11332, n11333, n11334, n11335, n11336, n11337,
         n11338, n11339, n11340, n11341, n11342, n11343, n11344, n11345,
         n11346, n11347, n11348, n11349, n11350, n11351, n11352, n11353,
         n11354, n11355, n11356, n11357, n11358, n11359, n11360, n11361,
         n11362, n11363, n11364, n11365, n11366, n11367, n11368, n11369,
         n11370, n11371, n11372, n11373, n11374, n11375, n11376, n11377,
         n11378, n11379, n11380, n11381, n11382, n11383, n11384, n11385,
         n11386, n11387, n11388, n11389, n11390, n11391, n11392, n11393,
         n11394, n11395, n11396, n11397, n11398, n11399, n11400, n11401,
         n11402, n11403, n11404, n11405, n11406, n11407, n11408, n11409,
         n11410, n11411, n11412, n11413, n11414, n11415, n11416, n11417,
         n11418, n11419, n11420, n11421, n11422, n11423, n11424, n11425,
         n11426, n11427, n11428, n11429, n11430, n11431, n11432, n11433,
         n11434, n11435, n11436, n11437, n11438, n11439, n11440, n11441,
         n11442, n11443, n11444, n11445, n11446, n11447, n11448, n11449,
         n11450, n11451, n11452, n11453, n11454, n11455, n11456, n11457,
         n11458, n11459, n11460, n11461, n11462, n11463, n11464, n11465,
         n11466, n11467, n11468, n11469, n11470, n11471, n11472, n11473,
         n11474, n11475, n11476, n11477, n11478, n11479, n11480, n11481,
         n11482, n11483, n11484, n11485, n11486, n11487, n11488, n11489,
         n11490, n11491, n11492, n11493, n11494, n11495, n11496, n11497,
         n11498, n11499, n11500, n11501, n11502, n11503, n11504, n11505,
         n11506, n11507, n11508, n11509, n11510, n11511, n11512, n11513,
         n11514, n11515, n11516, n11517, n11518, n11519, n11520, n11521,
         n11522, n11523, n11524, n11525, n11526, n11527, n11528, n11529,
         n11530, n11531, n11532, n11533, n11534, n11535, n11536, n11537,
         n11538, n11539, n11540, n11541, n11542, n11543, n11544, n11545,
         n11546, n11547, n11548, n11549, n11550, n11551, n11552, n11553,
         n11554, n11555, n11556, n11557, n11558, n11559, n11560, n11561,
         n11562, n11563, n11564, n11565, n11566, n11567, n11568, n11569,
         n11570, n11571, n11572, n11573, n11574, n11575, n11576, n11577,
         n11578, n11579, n11580, n11581, n11582, n11583, n11584, n11585,
         n11586, n11587, n11588, n11589, n11590, n11591, n11592, n11593,
         n11594, n11595, n11596, n11597, n11598, n11599, n11600, n11601,
         n11602, n11603, n11604, n11605, n11606, n11607, n11608, n11609,
         n11610, n11611, n11612, n11613, n11614, n11615, n11616, n11617,
         n11618, n11619, n11620, n11621, n11622, n11623, n11624, n11625,
         n11626, n11627, n11628, n11629, n11630, n11631, n11632, n11633,
         n11634, n11635, n11636, n11637, n11638, n11639, n11640, n11641,
         n11642, n11643, n11644, n11645, n11646, n11647, n11648, n11649,
         n11650, n11651, n11652, n11653, n11654, n11655, n11656, n11657,
         n11658, n11659, n11660, n11661, n11662, n11663, n11664, n11665,
         n11666, n11667, n11668, n11669, n11670, n11671, n11672, n11673,
         n11674, n11675, n11676, n11677, n11678, n11679, n11680, n11681,
         n11682, n11683, n11684, n11685, n11686, n11687, n11688, n11689,
         n11690, n11691, n11692, n11693, n11694, n11695, n11696, n11697,
         n11698, n11699, n11700, n11701, n11702, n11703, n11704, n11705,
         n11706, n11707, n11708, n11709, n11710, n11711, n11712, n11713,
         n11714, n11715, n11716, n11717, n11718, n11719, n11720, n11721,
         n11722, n11723, n11724, n11725, n11726, n11727, n11728, n11729,
         n11730, n11731, n11732, n11733, n11734, n11735, n11736, n11737,
         n11738, n11739, n11740, n11741, n11742, n11743, n11744, n11745,
         n11746, n11747, n11748, n11749, n11750, n11751, n11752, n11753,
         n11754, n11755, n11756, n11757, n11758, n11759, n11760, n11761,
         n11762, n11763, n11764, n11765, n11766, n11767, n11768, n11769,
         n11770, n11771, n11772, n11773, n11774, n11775, n11776, n11777,
         n11778, n11779, n11780, n11781, n11782, n11783, n11784, n11785,
         n11786, n11787, n11788, n11789, n11790, n11791, n11792, n11793,
         n11794, n11795, n11796, n11797, n11798, n11799, n11800, n11801,
         n11802, n11803, n11804, n11805, n11806, n11807, n11808, n11809,
         n11810, n11811, n11812, n11813, n11814, n11815, n11816, n11817,
         n11818, n11819, n11820, n11821, n11822, n11823, n11824, n11825,
         n11826, n11827, n11828, n11829, n11830, n11831, n11832, n11833,
         n11834, n11835, n11836, n11837, n11838, n11839, n11840, n11841,
         n11842, n11843, n11844, n11845, n11846, n11847, n11848, n11849,
         n11850, n11851, n11852, n11853, n11854, n11855, n11856, n11857,
         n11858, n11859, n11860, n11861, n11862, n11863, n11864, n11865,
         n11866, n11867, n11868, n11869, n11870, n11871, n11872, n11873,
         n11874, n11875, n11876, n11877, n11878, n11879, n11880, n11881,
         n11882, n11883, n11884, n11885, n11886, n11887, n11888, n11889,
         n11890, n11891, n11892, n11893, n11894, n11895, n11896, n11897,
         n11898, n11899, n11900, n11901, n11902, n11903, n11904, n11905,
         n11906, n11907, n11908, n11909, n11910, n11911, n11912, n11913,
         n11914, n11915, n11916, n11917, n11918, n11919, n11920, n11921,
         n11922, n11923, n11924, n11925, n11926, n11927, n11928, n11929,
         n11930, n11931, n11932, n11933, n11934, n11935, n11936, n11937,
         n11938, n11939, n11940, n11941, n11942, n11943, n11944, n11945,
         n11946, n11947, n11948, n11949, n11950, n11951, n11952, n11953,
         n11954, n11955, n11956, n11957, n11958, n11959, n11960, n11961,
         n11962, n11963, n11964, n11965, n11966, n11967, n11968, n11969,
         n11970, n11971, n11972, n11973, n11974, n11975, n11976, n11977,
         n11978, n11979, n11980, n11981, n11982, n11983, n11984, n11985,
         n11986, n11987, n11988, n11989, n11990, n11991, n11992, n11993,
         n11994, n11995, n11996, n11997, n11998, n11999, n12000, n12001,
         n12002, n12003, n12004, n12005, n12006, n12007, n12008, n12009,
         n12010, n12011, n12012, n12013, n12014, n12015, n12016, n12017,
         n12018, n12019, n12020, n12021, n12022, n12023, n12024, n12025,
         n12026, n12027, n12028, n12029, n12030, n12031, n12032, n12033,
         n12034, n12035, n12036, n12037, n12038, n12039, n12040, n12041,
         n12042, n12043, n12044, n12045, n12046, n12047, n12048, n12049,
         n12050, n12051, n12052, n12053, n12054, n12055, n12056, n12057,
         n12058, n12059, n12060, n12061, n12062, n12063, n12064, n12065,
         n12066, n12067, n12068, n12069, n12070, n12071, n12072, n12073,
         n12074, n12075, n12076, n12077, n12078, n12079, n12080, n12081,
         n12082, n12083, n12084, n12085, n12086, n12087, n12088, n12089,
         n12090, n12091, n12092, n12093, n12094, n12095, n12096, n12097,
         n12098, n12099, n12100, n12101, n12102, n12103, n12104, n12105,
         n12106, n12107, n12108, n12109, n12110, n12111, n12112, n12113,
         n12114, n12115, n12116, n12117, n12118, n12119, n12120, n12121,
         n12122, n12123, n12124, n12125, n12126, n12127, n12128, n12129,
         n12130, n12131, n12132, n12133, n12134, n12135, n12136, n12137,
         n12138, n12139, n12140, n12141, n12142, n12143, n12144, n12145,
         n12146, n12147, n12148, n12149, n12150, n12151, n12152, n12153,
         n12154, n12155, n12156, n12157, n12158, n12159, n12160, n12161,
         n12162, n12163, n12164, n12165, n12166, n12167, n12168, n12169,
         n12170, n12171, n12172, n12173, n12174, n12175, n12176, n12177,
         n12178, n12179, n12180, n12181, n12182, n12183, n12184, n12185,
         n12186, n12187, n12188, n12189, n12190, n12191, n12192, n12193,
         n12194, n12195, n12196, n12197, n12198, n12199, n12200, n12201,
         n12202, n12203, n12204, n12205, n12206, n12207, n12208, n12209,
         n12210, n12211, n12212, n12213, n12214, n12215, n12216, n12217,
         n12218, n12219, n12220, n12221, n12222, n12223, n12224, n12225,
         n12226, n12227, n12228, n12229, n12230, n12231, n12232, n12233,
         n12234, n12235, n12236, n12237, n12238, n12239, n12240, n12241,
         n12242, n12243, n12244, n12245, n12246, n12247, n12248, n12249,
         n12250, n12251, n12252, n12253, n12254, n12255, n12256, n12257,
         n12258, n12259, n12260, n12261, n12262, n12263, n12264, n12265,
         n12266, n12267, n12268, n12269, n12270, n12271, n12272, n12273,
         n12274, n12275, n12276, n12277, n12278, n12279, n12280, n12281,
         n12282, n12283, n12284, n12285, n12286, n12287, n12288, n12289,
         n12290, n12291, n12292, n12293, n12294, n12295, n12296, n12297,
         n12298, n12299, n12300, n12301, n12302, n12303, n12304, n12305,
         n12306, n12307, n12308, n12309, n12310, n12311, n12312, n12313,
         n12314, n12315, n12316, n12317, n12318, n12319, n12320, n12321,
         n12322, n12323, n12324, n12325, n12326, n12327, n12328, n12329,
         n12330, n12331, n12332, n12333, n12334, n12335, n12336, n12337,
         n12338, n12339, n12340, n12341, n12342, n12343, n12344, n12345,
         n12346, n12347, n12348, n12349, n12350, n12351, n12352, n12353,
         n12354, n12355, n12356, n12357, n12358, n12359, n12360, n12361,
         n12362, n12363, n12364, n12365, n12366, n12367, n12368, n12369,
         n12370, n12371, n12372, n12373, n12374, n12375, n12376, n12377,
         n12378, n12379, n12380, n12381, n12382, n12383, n12384, n12385,
         n12386, n12387, n12388, n12389, n12390, n12391, n12392, n12393,
         n12394, n12395, n12396, n12397, n12398, n12399, n12400, n12401,
         n12402, n12403, n12404, n12405, n12406, n12407, n12408, n12409,
         n12410, n12411, n12412, n12413, n12414, n12415, n12416, n12417,
         n12418, n12419, n12420, n12421, n12422, n12423, n12424, n12425,
         n12426, n12427, n12428, n12429, n12430, n12431, n12432, n12433,
         n12434, n12435, n12436, n12437, n12438, n12439, n12440, n12441,
         n12442, n12443, n12444, n12445, n12446, n12447, n12448, n12449,
         n12450, n12451, n12452, n12453, n12454, n12455, n12456, n12457,
         n12458, n12459, n12460, n12461, n12462, n12463, n12464, n12465,
         n12466, n12467, n12468, n12469, n12470, n12471, n12472, n12473,
         n12474, n12475, n12476, n12477, n12478, n12479, n12480, n12481,
         n12482, n12483, n12484, n12485, n12486, n12487, n12488, n12489,
         n12490, n12491, n12492, n12493, n12494, n12495, n12496, n12497,
         n12498, n12499, n12500, n12501, n12502, n12503, n12504, n12505,
         n12506, n12507, n12508, n12509, n12510, n12511, n12512, n12513,
         n12514, n12515, n12516, n12517, n12518, n12519, n12520, n12521,
         n12522, n12523, n12524, n12525, n12526, n12527, n12528, n12529,
         n12530, n12531, n12532, n12533, n12534, n12535, n12536, n12537,
         n12538, n12539, n12540, n12541, n12542, n12543, n12544, n12545,
         n12546, n12547, n12548, n12549, n12550, n12551, n12552, n12553,
         n12554, n12555, n12556, n12557, n12558, n12559, n12560, n12561,
         n12562, n12563, n12564, n12565, n12566, n12567, n12568, n12569,
         n12570, n12571, n12572, n12573, n12574, n12575, n12576, n12577,
         n12578, n12579, n12580, n12581, n12582, n12583, n12584, n12585,
         n12586, n12587, n12588, n12589, n12590, n12591, n12592, n12593,
         n12594, n12595, n12596, n12597, n12598, n12599, n12600, n12601,
         n12602, n12603, n12604, n12605, n12606, n12607, n12608, n12609,
         n12610, n12611, n12612, n12613, n12614, n12615, n12616, n12617,
         n12618, n12619, n12620, n12621, n12622, n12623, n12624, n12625,
         n12626, n12627, n12628, n12629, n12630, n12631, n12632, n12633,
         n12634, n12635, n12636, n12637, n12638, n12639, n12640, n12641,
         n12642, n12643, n12644, n12645, n12646, n12647, n12648, n12649,
         n12650, n12651, n12652, n12653, n12654, n12655, n12656, n12657,
         n12658, n12659, n12660, n12661, n12662, n12663, n12664, n12665,
         n12666, n12667, n12668, n12669, n12670, n12671, n12672, n12673,
         n12674, n12675, n12676, n12677, n12678, n12679, n12680, n12681,
         n12682, n12683, n12684, n12685, n12686, n12687, n12688, n12689,
         n12690, n12691, n12692, n12693, n12694, n12695, n12696, n12697,
         n12698, n12699, n12700, n12701, n12702, n12703, n12704, n12705,
         n12706, n12707, n12708, n12709, n12710, n12711, n12712, n12713,
         n12714, n12715, n12716, n12717, n12718, n12719, n12720, n12721,
         n12722, n12723, n12724, n12725, n12726, n12727, n12728, n12729,
         n12730, n12731, n12732, n12733, n12734, n12735, n12736, n12737,
         n12738, n12739, n12740, n12741, n12742, n12743, n12744, n12745,
         n12746, n12747, n12748, n12749, n12750, n12751, n12752, n12753,
         n12754, n12755, n12756, n12757, n12758, n12759, n12760, n12761,
         n12762, n12763, n12764, n12765, n12766, n12767, n12768, n12769,
         n12770, n12771, n12772, n12773, n12774, n12775, n12776, n12777,
         n12778, n12779, n12780, n12781, n12782, n12783, n12784, n12785,
         n12786, n12787, n12788, n12789, n12790, n12791, n12792, n12793,
         n12794, n12795, n12796, n12797, n12798, n12799, n12800, n12801,
         n12802, n12803, n12804, n12805, n12806, n12807, n12808, n12809,
         n12810, n12811, n12812, n12813, n12814, n12815, n12816, n12817,
         n12818, n12819, n12820, n12821, n12822, n12823, n12824, n12825,
         n12826, n12827, n12828, n12829, n12830, n12831, n12832, n12833,
         n12834, n12835, n12836, n12837, n12838, n12839, n12840, n12841,
         n12842, n12843, n12844, n12845, n12846, n12847, n12848, n12849,
         n12850, n12851, n12852, n12853, n12854, n12855, n12856, n12857,
         n12858, n12859, n12860, n12861, n12862, n12863, n12864, n12865,
         n12866, n12867, n12868, n12869, n12870, n12871, n12872, n12873,
         n12874, n12875, n12876, n12877, n12878, n12879, n12880, n12881,
         n12882, n12883, n12884, n12885, n12886, n12887, n12888, n12889,
         n12890, n12891, n12892, n12893, n12894, n12895, n12896, n12897,
         n12898, n12899, n12900, n12901, n12902, n12903, n12904, n12905,
         n12906, n12907, n12908, n12909, n12910, n12911, n12912, n12913,
         n12914, n12915, n12916, n12917, n12918, n12919, n12920, n12921,
         n12922, n12923, n12924, n12925, n12926, n12927, n12928, n12929,
         n12930, n12931, n12932, n12933, n12934, n12935, n12936, n12937,
         n12938, n12939, n12940, n12941, n12942, n12943, n12944, n12945,
         n12946, n12947, n12948, n12949, n12950, n12951, n12952, n12953,
         n12954, n12955, n12956, n12957, n12958, n12959, n12960, n12961,
         n12962, n12963, n12964, n12965, n12966, n12967, n12968, n12969,
         n12970, n12971, n12972, n12973, n12974, n12975, n12976, n12977,
         n12978, n12979, n12980, n12981, n12982, n12983, n12984, n12985,
         n12986, n12987, n12988, n12989, n12990, n12991, n12992, n12993,
         n12994, n12995, n12996, n12997, n12998, n12999, n13000, n13001,
         n13002, n13003, n13004, n13005, n13006, n13007, n13008, n13009,
         n13010, n13011, n13012, n13013, n13014, n13015, n13016, n13017,
         n13018, n13019, n13020, n13021, n13022, n13023, n13024, n13025,
         n13026, n13027, n13028, n13029, n13030, n13031, n13032, n13033,
         n13034, n13035, n13036, n13037, n13038, n13039, n13040, n13041,
         n13042, n13043, n13044, n13045, n13046, n13047, n13048, n13049,
         n13050, n13051, n13052, n13053, n13054, n13055, n13056, n13057,
         n13058, n13059, n13060, n13061, n13062, n13063, n13064, n13065,
         n13066, n13067, n13068, n13069, n13070, n13071, n13072, n13073,
         n13074, n13075, n13076, n13077, n13078, n13079, n13080, n13081,
         n13082, n13083, n13084, n13085, n13086, n13087, n13088, n13089,
         n13090, n13091, n13092, n13093, n13094, n13095, n13096, n13097,
         n13098, n13099, n13100, n13101, n13102, n13103, n13104, n13105,
         n13106, n13107, n13108, n13109, n13110, n13111, n13112, n13113,
         n13114, n13115, n13116, n13117, n13118, n13119, n13120, n13121,
         n13122, n13123, n13124, n13125, n13126, n13127, n13128, n13129,
         n13130, n13131, n13132, n13133, n13134, n13135, n13136, n13137,
         n13138, n13139, n13140, n13141, n13142, n13143, n13144, n13145,
         n13146, n13147, n13148, n13149, n13150, n13151, n13152, n13153,
         n13154, n13155, n13156, n13157, n13158, n13159, n13160, n13161,
         n13162, n13163, n13164, n13165, n13166, n13167, n13168, n13169,
         n13170, n13171, n13172, n13173, n13174, n13175, n13176, n13177,
         n13178, n13179, n13180, n13181, n13182, n13183, n13184, n13185,
         n13186, n13187, n13188, n13189, n13190, n13191, n13192, n13193,
         n13194, n13195, n13196, n13197, n13198, n13199, n13200, n13201,
         n13202, n13203, n13204, n13205, n13206, n13207, n13208, n13209,
         n13210, n13211, n13212, n13213, n13214, n13215, n13216, n13217,
         n13218, n13219, n13220, n13221, n13222, n13223, n13224, n13225,
         n13226, n13227, n13228, n13229, n13230, n13231, n13232, n13233,
         n13234, n13235, n13236, n13237, n13238, n13239, n13240, n13241,
         n13242, n13243, n13244, n13245, n13246, n13247, n13248, n13249,
         n13250, n13251, n13252, n13253, n13254, n13255, n13256, n13257,
         n13258, n13259, n13260, n13261, n13262, n13263, n13264, n13265,
         n13266, n13267, n13268, n13269, n13270, n13271, n13272, n13273,
         n13274, n13275, n13276, n13277, n13278, n13279, n13280, n13281,
         n13282, n13283, n13284, n13285, n13286, n13287, n13288, n13289,
         n13290, n13291, n13292, n13293, n13294, n13295, n13296, n13297,
         n13298, n13299, n13300, n13301, n13302, n13303, n13304, n13305,
         n13306, n13307, n13308, n13309, n13310, n13311, n13312, n13313,
         n13314, n13315, n13316, n13317, n13318, n13319, n13320, n13321,
         n13322, n13323, n13324, n13325, n13326, n13327, n13328, n13329,
         n13330, n13331, n13332, n13333, n13334, n13335, n13336, n13337,
         n13338, n13339, n13340, n13341, n13342, n13343, n13344, n13345,
         n13346, n13347, n13348, n13349, n13350, n13351, n13352, n13353,
         n13354, n13355, n13356, n13357, n13358, n13359, n13360, n13361,
         n13362, n13363, n13364, n13365, n13366, n13367, n13368, n13369,
         n13370, n13371, n13372, n13373, n13374, n13375, n13376, n13377,
         n13378, n13379, n13380, n13381, n13382, n13383, n13384, n13385,
         n13386, n13387, n13388, n13389, n13390, n13391, n13392, n13393,
         n13394, n13395, n13396, n13397, n13398, n13399, n13400, n13401,
         n13402, n13403, n13404, n13405, n13406, n13407, n13408, n13409,
         n13410, n13411, n13412, n13413, n13414, n13415, n13416, n13417,
         n13418, n13419, n13420, n13421, n13422, n13423, n13424, n13425,
         n13426, n13427, n13428, n13429, n13430, n13431, n13432, n13433,
         n13434, n13435, n13436, n13437, n13438, n13439, n13440, n13441,
         n13442, n13443, n13444, n13445, n13446, n13447, n13448, n13449,
         n13450, n13451, n13452, n13453, n13454, n13455, n13456, n13457,
         n13458, n13459, n13460, n13461, n13462, n13463, n13464, n13465,
         n13466, n13467, n13468, n13469, n13470, n13471, n13472, n13473,
         n13474, n13475, n13476, n13477, n13478, n13479, n13480, n13481,
         n13482, n13483, n13484, n13485, n13486, n13487, n13488, n13489,
         n13490, n13491, n13492, n13493, n13494, n13495, n13496, n13497,
         n13498, n13499, n13500, n13501, n13502, n13503, n13504, n13505,
         n13506, n13507, n13508, n13509, n13510, n13511, n13512, n13513,
         n13514, n13515, n13516, n13517, n13518, n13519, n13520, n13521,
         n13522, n13523, n13524, n13525, n13526, n13527, n13528, n13529,
         n13530, n13531, n13532, n13533, n13534, n13535, n13536, n13537,
         n13538, n13539, n13540, n13541, n13542, n13543, n13544, n13545,
         n13546, n13547, n13548, n13549, n13550, n13551, n13552, n13553,
         n13554, n13555, n13556, n13557, n13558, n13559, n13560, n13561,
         n13562, n13563, n13564, n13565, n13566, n13567, n13568, n13569,
         n13570, n13571, n13572, n13573, n13574, n13575, n13576, n13577,
         n13578, n13579, n13580, n13581, n13582, n13583, n13584, n13585,
         n13586, n13587, n13588, n13589, n13590, n13591, n13592, n13593,
         n13594, n13595, n13596, n13597, n13598, n13599, n13600, n13601,
         n13602, n13603, n13604, n13605, n13606, n13607, n13608, n13609,
         n13610, n13611, n13612, n13613, n13614, n13615, n13616, n13617,
         n13618, n13619, n13620, n13621, n13622, n13623, n13624, n13625,
         n13626, n13627, n13628, n13629, n13630, n13631, n13632, n13633,
         n13634, n13635, n13636, n13637, n13638, n13639, n13640, n13641,
         n13642, n13643, n13644, n13645, n13646, n13647, n13648, n13649,
         n13650, n13651, n13652, n13653, n13654, n13655, n13656, n13657,
         n13658, n13659, n13660, n13661, n13662, n13663, n13664, n13665,
         n13666, n13667, n13668, n13669, n13670, n13671, n13672, n13673,
         n13674, n13675, n13676, n13677, n13678, n13679, n13680, n13681,
         n13682, n13683, n13684, n13685, n13686, n13687, n13688, n13689,
         n13690, n13691, n13692, n13693, n13694, n13695, n13696, n13697,
         n13698, n13699, n13700, n13701, n13702, n13703, n13704, n13705,
         n13706, n13707, n13708, n13709, n13710, n13711, n13712, n13713,
         n13714, n13715, n13716, n13717, n13718, n13719, n13720, n13721,
         n13722, n13723, n13724, n13725, n13726, n13727, n13728, n13729,
         n13730, n13731, n13732, n13733, n13734, n13735, n13736, n13737,
         n13738, n13739, n13740, n13741, n13742, n13743, n13744, n13745,
         n13746, n13747, n13748, n13749, n13750, n13751, n13752, n13753,
         n13754, n13755, n13756, n13757, n13758, n13759, n13760, n13761,
         n13762, n13763, n13764, n13765, n13766, n13767, n13768, n13769,
         n13770, n13771, n13772, n13773, n13774, n13775, n13776, n13777,
         n13778, n13779, n13780, n13781, n13782, n13783, n13784, n13785,
         n13786, n13787, n13788, n13789, n13790, n13791, n13792, n13793,
         n13794, n13795, n13796, n13797, n13798, n13799, n13800, n13801,
         n13802, n13803, n13804, n13805, n13806, n13807, n13808, n13809,
         n13810, n13811, n13812, n13813, n13814, n13815, n13816, n13817,
         n13818, n13819, n13820, n13821, n13822, n13823, n13824, n13825,
         n13826, n13827, n13828, n13829, n13830, n13831, n13832, n13833,
         n13834, n13835, n13836, n13837, n13838, n13839, n13840, n13841,
         n13842, n13843, n13844, n13845, n13846, n13847, n13848, n13849,
         n13850, n13851, n13852, n13853, n13854, n13855, n13856, n13857,
         n13858, n13859, n13860, n13861, n13862, n13863, n13864, n13865,
         n13866, n13867, n13868, n13869, n13870, n13871, n13872, n13873,
         n13874, n13875, n13876, n13877, n13878, n13879, n13880, n13881,
         n13882, n13883, n13884, n13885, n13886, n13887, n13888, n13889,
         n13890, n13891, n13892, n13893, n13894, n13895, n13896, n13897,
         n13898, n13899, n13900, n13901, n13902, n13903, n13904, n13905,
         n13906, n13907, n13908, n13909, n13910, n13911, n13912, n13913,
         n13914, n13915, n13916, n13917, n13918, n13919, n13920, n13921,
         n13922, n13923, n13924, n13925, n13926, n13927, n13928, n13929,
         n13930, n13931, n13932, n13933, n13934, n13935, n13936, n13937,
         n13938, n13939, n13940, n13941, n13942, n13943, n13944, n13945,
         n13946, n13947, n13948, n13949, n13950, n13951, n13952, n13953,
         n13954, n13955, n13956, n13957, n13958, n13959, n13960, n13961,
         n13962, n13963, n13964, n13965, n13966, n13967, n13968, n13969,
         n13970, n13971, n13972, n13973, n13974, n13975, n13976, n13977,
         n13978, n13979, n13980, n13981, n13982, n13983, n13984, n13985,
         n13986, n13987, n13988, n13989, n13990, n13991, n13992, n13993,
         n13994, n13995, n13996, n13997, n13998, n13999, n14000, n14001,
         n14002, n14003, n14004, n14005, n14006, n14007, n14008, n14009,
         n14010, n14011, n14012, n14013, n14014, n14015, n14016, n14017,
         n14018, n14019, n14020, n14021, n14022, n14023, n14024, n14025,
         n14026, n14027, n14028, n14029, n14030, n14031, n14032, n14033,
         n14034, n14035, n14036, n14037, n14038, n14039, n14040, n14041,
         n14042, n14043, n14044, n14045, n14046, n14047, n14048, n14049,
         n14050, n14051, n14052, n14053, n14054, n14055, n14056, n14057,
         n14058, n14059, n14060, n14061, n14062, n14063, n14064, n14065,
         n14066, n14067, n14068, n14069, n14070, n14071, n14072, n14073,
         n14074, n14075, n14076, n14077, n14078, n14079, n14080, n14081,
         n14082, n14083, n14084, n14085, n14086, n14087, n14088, n14089,
         n14090, n14091, n14092, n14093, n14094, n14095, n14096, n14097,
         n14098, n14099, n14100, n14101, n14102, n14103, n14104, n14105,
         n14106, n14107, n14108, n14109, n14110, n14111, n14112, n14113,
         n14114, n14115, n14116, n14117, n14118, n14119, n14120, n14121,
         n14122, n14123, n14124, n14125, n14126, n14127, n14128, n14129,
         n14130, n14131, n14132, n14133, n14134, n14135, n14136, n14137,
         n14138, n14139, n14140, n14141, n14142, n14143, n14144, n14145,
         n14146, n14147, n14148, n14149, n14150, n14151, n14152, n14153,
         n14154, n14155, n14156, n14157, n14158, n14159, n14160, n14161,
         n14162, n14163, n14164, n14165, n14166, n14167, n14168, n14169,
         n14170, n14171, n14172, n14173, n14174, n14175, n14176, n14177,
         n14178, n14179, n14180, n14181, n14182, n14183, n14184, n14185,
         n14186, n14187, n14188, n14189, n14190, n14191, n14192, n14193,
         n14194, n14195, n14196, n14197, n14198, n14199, n14200, n14201,
         n14202, n14203, n14204, n14205, n14206, n14207, n14208, n14209,
         n14210, n14211, n14212, n14213, n14214, n14215, n14216, n14217,
         n14218, n14219, n14220, n14221, n14222, n14223, n14224, n14225,
         n14226, n14227, n14228, n14229, n14230, n14231, n14232, n14233,
         n14234, n14235, n14236, n14237, n14238, n14239, n14240, n14241,
         n14242, n14243, n14244, n14245, n14246, n14247, n14248, n14249,
         n14250, n14251, n14252, n14253, n14254, n14255, n14256, n14257,
         n14258, n14259, n14260, n14261, n14262, n14263, n14264, n14265,
         n14266, n14267, n14268, n14269, n14270, n14271, n14272, n14273,
         n14274, n14275, n14276, n14277, n14278, n14279, n14280, n14281,
         n14282, n14283, n14284, n14285, n14286, n14287, n14288, n14289,
         n14290, n14291, n14292, n14293, n14294, n14295, n14296, n14297,
         n14298, n14299, n14300, n14301, n14302, n14303, n14304, n14305,
         n14306, n14307, n14308, n14309, n14310, n14311, n14312, n14313,
         n14314, n14315, n14316, n14317, n14318, n14319, n14320, n14321,
         n14322, n14323, n14324, n14325, n14326, n14327, n14328, n14329,
         n14330, n14331, n14332, n14333, n14334, n14335, n14336, n14337,
         n14338, n14339, n14340, n14341, n14342, n14343, n14344, n14345,
         n14346, n14347, n14348, n14349, n14350, n14351, n14352, n14353,
         n14354, n14355, n14356, n14357, n14358, n14359, n14360, n14361,
         n14362, n14363, n14364, n14365, n14366, n14367, n14368, n14369,
         n14370, n14371, n14372, n14373, n14374, n14375, n14376, n14377,
         n14378, n14379, n14380, n14381, n14382, n14383, n14384, n14385,
         n14386, n14387, n14388, n14389, n14390, n14391, n14392, n14393,
         n14394, n14395, n14396, n14397, n14398, n14399, n14400, n14401,
         n14402, n14403, n14404, n14405, n14406, n14407, n14408, n14409,
         n14410, n14411, n14412, n14413, n14414, n14415, n14416, n14417,
         n14418, n14419, n14420, n14421, n14422, n14423, n14424, n14425,
         n14426, n14427, n14428, n14429, n14430, n14431, n14432, n14433,
         n14434, n14435, n14436, n14437, n14438, n14439, n14440, n14441,
         n14442, n14443, n14444, n14445, n14446, n14447, n14448, n14449,
         n14450, n14451, n14452, n14453, n14454, n14455, n14456, n14457,
         n14458, n14459, n14460, n14461, n14462, n14463, n14464, n14465,
         n14466, n14467, n14468, n14469, n14470, n14471, n14472, n14473,
         n14474, n14475, n14476, n14477, n14478, n14479, n14480, n14481,
         n14482, n14483, n14484, n14485, n14486, n14487, n14488, n14489,
         n14490, n14491, n14492, n14493, n14494, n14495, n14496, n14497,
         n14498, n14499, n14500, n14501, n14502, n14503, n14504, n14505,
         n14506, n14507, n14508, n14509, n14510, n14511, n14512, n14513,
         n14514, n14515, n14516, n14517, n14518, n14519, n14520, n14521,
         n14522, n14523, n14524, n14525, n14526, n14527, n14528, n14529,
         n14530, n14531, n14532, n14533, n14534, n14535, n14536, n14537,
         n14538, n14539, n14540, n14541, n14542, n14543, n14544, n14545,
         n14546, n14547, n14548, n14549, n14550, n14551, n14552;

  XNOR U1 ( .A(n1), .B(n2), .Z(o[9]) );
  AND U2 ( .A(o[6]), .B(n3), .Z(n1) );
  XOR U3 ( .A(n2), .B(n4), .Z(n3) );
  XOR U4 ( .A(n5), .B(n6), .Z(o[8]) );
  AND U5 ( .A(o[6]), .B(n7), .Z(n5) );
  XOR U6 ( .A(n8), .B(n9), .Z(n7) );
  XNOR U7 ( .A(n10), .B(n11), .Z(o[7]) );
  AND U8 ( .A(o[6]), .B(n12), .Z(n10) );
  XNOR U9 ( .A(n13), .B(n11), .Z(n12) );
  XOR U10 ( .A(n14), .B(n15), .Z(o[22]) );
  AND U11 ( .A(o[6]), .B(n16), .Z(n14) );
  XOR U12 ( .A(n17), .B(n18), .Z(n16) );
  XOR U13 ( .A(n19), .B(n20), .Z(o[21]) );
  AND U14 ( .A(o[6]), .B(n21), .Z(n19) );
  XOR U15 ( .A(n22), .B(n23), .Z(n21) );
  XOR U16 ( .A(n24), .B(n25), .Z(o[20]) );
  AND U17 ( .A(o[6]), .B(n26), .Z(n24) );
  XOR U18 ( .A(n27), .B(n28), .Z(n26) );
  XOR U19 ( .A(n29), .B(n30), .Z(o[19]) );
  AND U20 ( .A(o[6]), .B(n31), .Z(n29) );
  XOR U21 ( .A(n32), .B(n33), .Z(n31) );
  XOR U22 ( .A(n34), .B(n35), .Z(o[18]) );
  AND U23 ( .A(o[6]), .B(n36), .Z(n34) );
  XOR U24 ( .A(n37), .B(n38), .Z(n36) );
  XOR U25 ( .A(n39), .B(n40), .Z(o[17]) );
  AND U26 ( .A(o[6]), .B(n41), .Z(n39) );
  XOR U27 ( .A(n42), .B(n43), .Z(n41) );
  XOR U28 ( .A(n44), .B(n45), .Z(o[16]) );
  AND U29 ( .A(o[6]), .B(n46), .Z(n44) );
  XOR U30 ( .A(n47), .B(n48), .Z(n46) );
  XOR U31 ( .A(n49), .B(n50), .Z(o[15]) );
  AND U32 ( .A(o[6]), .B(n51), .Z(n49) );
  XOR U33 ( .A(n52), .B(n53), .Z(n51) );
  XOR U34 ( .A(n54), .B(n55), .Z(o[14]) );
  AND U35 ( .A(o[6]), .B(n56), .Z(n54) );
  XOR U36 ( .A(n57), .B(n58), .Z(n56) );
  XOR U37 ( .A(n59), .B(n60), .Z(o[13]) );
  AND U38 ( .A(o[6]), .B(n61), .Z(n59) );
  XOR U39 ( .A(n62), .B(n63), .Z(n61) );
  XOR U40 ( .A(n64), .B(n65), .Z(o[12]) );
  AND U41 ( .A(o[6]), .B(n66), .Z(n64) );
  XOR U42 ( .A(n67), .B(n68), .Z(n66) );
  XOR U43 ( .A(n69), .B(n70), .Z(o[11]) );
  AND U44 ( .A(o[6]), .B(n71), .Z(n69) );
  XOR U45 ( .A(n72), .B(n73), .Z(n71) );
  XOR U46 ( .A(n74), .B(n75), .Z(o[10]) );
  AND U47 ( .A(o[6]), .B(n76), .Z(n74) );
  XOR U48 ( .A(n77), .B(n78), .Z(n76) );
  XOR U49 ( .A(n79), .B(n80), .Z(o[0]) );
  AND U50 ( .A(o[1]), .B(n81), .Z(n80) );
  XNOR U51 ( .A(n82), .B(n83), .Z(n81) );
  XNOR U52 ( .A(n84), .B(n79), .Z(n83) );
  AND U53 ( .A(o[2]), .B(n85), .Z(n84) );
  XNOR U54 ( .A(n86), .B(n87), .Z(n85) );
  XNOR U55 ( .A(n88), .B(n82), .Z(n87) );
  AND U56 ( .A(o[3]), .B(n89), .Z(n88) );
  XNOR U57 ( .A(n90), .B(n91), .Z(n89) );
  XNOR U58 ( .A(n92), .B(n86), .Z(n91) );
  AND U59 ( .A(o[4]), .B(n93), .Z(n92) );
  XNOR U60 ( .A(n94), .B(n95), .Z(n93) );
  XNOR U61 ( .A(n96), .B(n90), .Z(n95) );
  AND U62 ( .A(o[5]), .B(n97), .Z(n96) );
  XNOR U63 ( .A(n94), .B(n98), .Z(n97) );
  XNOR U64 ( .A(n99), .B(n100), .Z(n98) );
  AND U65 ( .A(o[6]), .B(n101), .Z(n99) );
  XOR U66 ( .A(n100), .B(n102), .Z(n101) );
  XOR U67 ( .A(n103), .B(n104), .Z(n94) );
  AND U68 ( .A(o[6]), .B(n105), .Z(n104) );
  XOR U69 ( .A(n103), .B(n106), .Z(n105) );
  XOR U70 ( .A(n107), .B(n108), .Z(n90) );
  AND U71 ( .A(o[5]), .B(n109), .Z(n108) );
  XNOR U72 ( .A(n107), .B(n110), .Z(n109) );
  XNOR U73 ( .A(n111), .B(n112), .Z(n110) );
  AND U74 ( .A(o[6]), .B(n113), .Z(n111) );
  XOR U75 ( .A(n112), .B(n114), .Z(n113) );
  XOR U76 ( .A(n115), .B(n116), .Z(n107) );
  AND U77 ( .A(o[6]), .B(n117), .Z(n116) );
  XOR U78 ( .A(n115), .B(n118), .Z(n117) );
  XOR U79 ( .A(n119), .B(n120), .Z(n86) );
  AND U80 ( .A(o[4]), .B(n121), .Z(n120) );
  XNOR U81 ( .A(n122), .B(n123), .Z(n121) );
  XNOR U82 ( .A(n124), .B(n119), .Z(n123) );
  AND U83 ( .A(o[5]), .B(n125), .Z(n124) );
  XNOR U84 ( .A(n122), .B(n126), .Z(n125) );
  XNOR U85 ( .A(n127), .B(n128), .Z(n126) );
  AND U86 ( .A(o[6]), .B(n129), .Z(n127) );
  XOR U87 ( .A(n128), .B(n130), .Z(n129) );
  XOR U88 ( .A(n131), .B(n132), .Z(n122) );
  AND U89 ( .A(o[6]), .B(n133), .Z(n132) );
  XOR U90 ( .A(n131), .B(n134), .Z(n133) );
  XOR U91 ( .A(n135), .B(n136), .Z(n119) );
  AND U92 ( .A(o[5]), .B(n137), .Z(n136) );
  XNOR U93 ( .A(n135), .B(n138), .Z(n137) );
  XNOR U94 ( .A(n139), .B(n140), .Z(n138) );
  AND U95 ( .A(o[6]), .B(n141), .Z(n139) );
  XOR U96 ( .A(n140), .B(n142), .Z(n141) );
  XOR U97 ( .A(n143), .B(n144), .Z(n135) );
  AND U98 ( .A(o[6]), .B(n145), .Z(n144) );
  XOR U99 ( .A(n143), .B(n146), .Z(n145) );
  XOR U100 ( .A(n147), .B(n148), .Z(n82) );
  AND U101 ( .A(o[3]), .B(n149), .Z(n148) );
  XNOR U102 ( .A(n150), .B(n151), .Z(n149) );
  XNOR U103 ( .A(n152), .B(n147), .Z(n151) );
  AND U104 ( .A(o[4]), .B(n153), .Z(n152) );
  XNOR U105 ( .A(n154), .B(n155), .Z(n153) );
  XNOR U106 ( .A(n156), .B(n150), .Z(n155) );
  AND U107 ( .A(o[5]), .B(n157), .Z(n156) );
  XNOR U108 ( .A(n154), .B(n158), .Z(n157) );
  XNOR U109 ( .A(n159), .B(n160), .Z(n158) );
  AND U110 ( .A(o[6]), .B(n161), .Z(n159) );
  XOR U111 ( .A(n160), .B(n162), .Z(n161) );
  XOR U112 ( .A(n163), .B(n164), .Z(n154) );
  AND U113 ( .A(o[6]), .B(n165), .Z(n164) );
  XOR U114 ( .A(n163), .B(n166), .Z(n165) );
  XOR U115 ( .A(n167), .B(n168), .Z(n150) );
  AND U116 ( .A(o[5]), .B(n169), .Z(n168) );
  XNOR U117 ( .A(n167), .B(n170), .Z(n169) );
  XNOR U118 ( .A(n171), .B(n172), .Z(n170) );
  AND U119 ( .A(o[6]), .B(n173), .Z(n171) );
  XOR U120 ( .A(n172), .B(n174), .Z(n173) );
  XOR U121 ( .A(n175), .B(n176), .Z(n167) );
  AND U122 ( .A(o[6]), .B(n177), .Z(n176) );
  XOR U123 ( .A(n175), .B(n178), .Z(n177) );
  XOR U124 ( .A(n179), .B(n180), .Z(n147) );
  AND U125 ( .A(o[4]), .B(n181), .Z(n180) );
  XNOR U126 ( .A(n182), .B(n183), .Z(n181) );
  XNOR U127 ( .A(n184), .B(n179), .Z(n183) );
  AND U128 ( .A(o[5]), .B(n185), .Z(n184) );
  XNOR U129 ( .A(n182), .B(n186), .Z(n185) );
  XNOR U130 ( .A(n187), .B(n188), .Z(n186) );
  AND U131 ( .A(o[6]), .B(n189), .Z(n187) );
  XOR U132 ( .A(n188), .B(n190), .Z(n189) );
  XOR U133 ( .A(n191), .B(n192), .Z(n182) );
  AND U134 ( .A(o[6]), .B(n193), .Z(n192) );
  XOR U135 ( .A(n191), .B(n194), .Z(n193) );
  XOR U136 ( .A(n195), .B(n196), .Z(n179) );
  AND U137 ( .A(o[5]), .B(n197), .Z(n196) );
  XNOR U138 ( .A(n195), .B(n198), .Z(n197) );
  XNOR U139 ( .A(n199), .B(n200), .Z(n198) );
  AND U140 ( .A(o[6]), .B(n201), .Z(n199) );
  XOR U141 ( .A(n200), .B(n202), .Z(n201) );
  XOR U142 ( .A(n203), .B(n204), .Z(n195) );
  AND U143 ( .A(o[6]), .B(n205), .Z(n204) );
  XOR U144 ( .A(n203), .B(n206), .Z(n205) );
  XOR U145 ( .A(n207), .B(n208), .Z(o[1]) );
  AND U146 ( .A(o[2]), .B(n209), .Z(n208) );
  XNOR U147 ( .A(n210), .B(n211), .Z(n209) );
  XNOR U148 ( .A(n212), .B(n207), .Z(n211) );
  AND U149 ( .A(o[3]), .B(n213), .Z(n212) );
  XNOR U150 ( .A(n214), .B(n215), .Z(n213) );
  XNOR U151 ( .A(n216), .B(n210), .Z(n215) );
  AND U152 ( .A(o[4]), .B(n217), .Z(n216) );
  XNOR U153 ( .A(n218), .B(n219), .Z(n217) );
  XNOR U154 ( .A(n220), .B(n214), .Z(n219) );
  AND U155 ( .A(o[5]), .B(n221), .Z(n220) );
  XNOR U156 ( .A(n218), .B(n222), .Z(n221) );
  XNOR U157 ( .A(n223), .B(n224), .Z(n222) );
  AND U158 ( .A(o[6]), .B(n225), .Z(n223) );
  XOR U159 ( .A(n224), .B(n226), .Z(n225) );
  XOR U160 ( .A(n227), .B(n228), .Z(n218) );
  AND U161 ( .A(o[6]), .B(n229), .Z(n228) );
  XOR U162 ( .A(n227), .B(n230), .Z(n229) );
  XOR U163 ( .A(n231), .B(n232), .Z(n214) );
  AND U164 ( .A(o[5]), .B(n233), .Z(n232) );
  XNOR U165 ( .A(n231), .B(n234), .Z(n233) );
  XNOR U166 ( .A(n235), .B(n236), .Z(n234) );
  AND U167 ( .A(o[6]), .B(n237), .Z(n235) );
  XOR U168 ( .A(n236), .B(n238), .Z(n237) );
  XOR U169 ( .A(n239), .B(n240), .Z(n231) );
  AND U170 ( .A(o[6]), .B(n241), .Z(n240) );
  XOR U171 ( .A(n239), .B(n242), .Z(n241) );
  XOR U172 ( .A(n243), .B(n244), .Z(n210) );
  AND U173 ( .A(o[4]), .B(n245), .Z(n244) );
  XNOR U174 ( .A(n246), .B(n247), .Z(n245) );
  XNOR U175 ( .A(n248), .B(n243), .Z(n247) );
  AND U176 ( .A(o[5]), .B(n249), .Z(n248) );
  XNOR U177 ( .A(n246), .B(n250), .Z(n249) );
  XNOR U178 ( .A(n251), .B(n252), .Z(n250) );
  AND U179 ( .A(o[6]), .B(n253), .Z(n251) );
  XOR U180 ( .A(n252), .B(n254), .Z(n253) );
  XOR U181 ( .A(n255), .B(n256), .Z(n246) );
  AND U182 ( .A(o[6]), .B(n257), .Z(n256) );
  XOR U183 ( .A(n255), .B(n258), .Z(n257) );
  XOR U184 ( .A(n259), .B(n260), .Z(n243) );
  AND U185 ( .A(o[5]), .B(n261), .Z(n260) );
  XNOR U186 ( .A(n259), .B(n262), .Z(n261) );
  XNOR U187 ( .A(n263), .B(n264), .Z(n262) );
  AND U188 ( .A(o[6]), .B(n265), .Z(n263) );
  XOR U189 ( .A(n264), .B(n266), .Z(n265) );
  XOR U190 ( .A(n267), .B(n268), .Z(n259) );
  AND U191 ( .A(o[6]), .B(n269), .Z(n268) );
  XOR U192 ( .A(n267), .B(n270), .Z(n269) );
  XOR U193 ( .A(n271), .B(n272), .Z(n207) );
  AND U194 ( .A(o[3]), .B(n273), .Z(n272) );
  XNOR U195 ( .A(n274), .B(n275), .Z(n273) );
  XNOR U196 ( .A(n276), .B(n271), .Z(n275) );
  AND U197 ( .A(o[4]), .B(n277), .Z(n276) );
  XNOR U198 ( .A(n278), .B(n279), .Z(n277) );
  XNOR U199 ( .A(n280), .B(n274), .Z(n279) );
  AND U200 ( .A(o[5]), .B(n281), .Z(n280) );
  XNOR U201 ( .A(n278), .B(n282), .Z(n281) );
  XNOR U202 ( .A(n283), .B(n284), .Z(n282) );
  AND U203 ( .A(o[6]), .B(n285), .Z(n283) );
  XOR U204 ( .A(n284), .B(n286), .Z(n285) );
  XOR U205 ( .A(n287), .B(n288), .Z(n278) );
  AND U206 ( .A(o[6]), .B(n289), .Z(n288) );
  XOR U207 ( .A(n287), .B(n290), .Z(n289) );
  XOR U208 ( .A(n291), .B(n292), .Z(n274) );
  AND U209 ( .A(o[5]), .B(n293), .Z(n292) );
  XNOR U210 ( .A(n291), .B(n294), .Z(n293) );
  XNOR U211 ( .A(n295), .B(n296), .Z(n294) );
  AND U212 ( .A(o[6]), .B(n297), .Z(n295) );
  XOR U213 ( .A(n296), .B(n298), .Z(n297) );
  XOR U214 ( .A(n299), .B(n300), .Z(n291) );
  AND U215 ( .A(o[6]), .B(n301), .Z(n300) );
  XOR U216 ( .A(n299), .B(n302), .Z(n301) );
  XOR U217 ( .A(n303), .B(n304), .Z(n271) );
  AND U218 ( .A(o[4]), .B(n305), .Z(n304) );
  XNOR U219 ( .A(n306), .B(n307), .Z(n305) );
  XNOR U220 ( .A(n308), .B(n303), .Z(n307) );
  AND U221 ( .A(o[5]), .B(n309), .Z(n308) );
  XNOR U222 ( .A(n306), .B(n310), .Z(n309) );
  XNOR U223 ( .A(n311), .B(n312), .Z(n310) );
  AND U224 ( .A(o[6]), .B(n313), .Z(n311) );
  XOR U225 ( .A(n312), .B(n314), .Z(n313) );
  XOR U226 ( .A(n315), .B(n316), .Z(n306) );
  AND U227 ( .A(o[6]), .B(n317), .Z(n316) );
  XOR U228 ( .A(n315), .B(n318), .Z(n317) );
  XOR U229 ( .A(n319), .B(n320), .Z(n303) );
  AND U230 ( .A(o[5]), .B(n321), .Z(n320) );
  XNOR U231 ( .A(n319), .B(n322), .Z(n321) );
  XNOR U232 ( .A(n323), .B(n324), .Z(n322) );
  AND U233 ( .A(o[6]), .B(n325), .Z(n323) );
  XOR U234 ( .A(n324), .B(n326), .Z(n325) );
  XOR U235 ( .A(n327), .B(n328), .Z(n319) );
  AND U236 ( .A(o[6]), .B(n329), .Z(n328) );
  XOR U237 ( .A(n327), .B(n330), .Z(n329) );
  XOR U238 ( .A(n331), .B(n332), .Z(n79) );
  AND U239 ( .A(o[2]), .B(n333), .Z(n332) );
  XNOR U240 ( .A(n334), .B(n335), .Z(n333) );
  XNOR U241 ( .A(n336), .B(n331), .Z(n335) );
  AND U242 ( .A(o[3]), .B(n337), .Z(n336) );
  XNOR U243 ( .A(n338), .B(n339), .Z(n337) );
  XNOR U244 ( .A(n340), .B(n334), .Z(n339) );
  AND U245 ( .A(o[4]), .B(n341), .Z(n340) );
  XNOR U246 ( .A(n342), .B(n343), .Z(n341) );
  XNOR U247 ( .A(n344), .B(n338), .Z(n343) );
  AND U248 ( .A(o[5]), .B(n345), .Z(n344) );
  XNOR U249 ( .A(n342), .B(n346), .Z(n345) );
  XNOR U250 ( .A(n347), .B(n348), .Z(n346) );
  AND U251 ( .A(o[6]), .B(n349), .Z(n347) );
  XOR U252 ( .A(n348), .B(n350), .Z(n349) );
  XOR U253 ( .A(n351), .B(n352), .Z(n342) );
  AND U254 ( .A(o[6]), .B(n353), .Z(n352) );
  XOR U255 ( .A(n351), .B(n354), .Z(n353) );
  XOR U256 ( .A(n355), .B(n356), .Z(n338) );
  AND U257 ( .A(o[5]), .B(n357), .Z(n356) );
  XNOR U258 ( .A(n355), .B(n358), .Z(n357) );
  XNOR U259 ( .A(n359), .B(n360), .Z(n358) );
  AND U260 ( .A(o[6]), .B(n361), .Z(n359) );
  XOR U261 ( .A(n360), .B(n362), .Z(n361) );
  XOR U262 ( .A(n363), .B(n364), .Z(n355) );
  AND U263 ( .A(o[6]), .B(n365), .Z(n364) );
  XOR U264 ( .A(n363), .B(n366), .Z(n365) );
  XOR U265 ( .A(n367), .B(n368), .Z(n334) );
  AND U266 ( .A(o[4]), .B(n369), .Z(n368) );
  XNOR U267 ( .A(n370), .B(n371), .Z(n369) );
  XNOR U268 ( .A(n372), .B(n367), .Z(n371) );
  AND U269 ( .A(o[5]), .B(n373), .Z(n372) );
  XNOR U270 ( .A(n370), .B(n374), .Z(n373) );
  XNOR U271 ( .A(n375), .B(n376), .Z(n374) );
  AND U272 ( .A(o[6]), .B(n377), .Z(n375) );
  XOR U273 ( .A(n376), .B(n378), .Z(n377) );
  XOR U274 ( .A(n379), .B(n380), .Z(n370) );
  AND U275 ( .A(o[6]), .B(n381), .Z(n380) );
  XOR U276 ( .A(n379), .B(n382), .Z(n381) );
  XOR U277 ( .A(n383), .B(n384), .Z(n367) );
  AND U278 ( .A(o[5]), .B(n385), .Z(n384) );
  XNOR U279 ( .A(n383), .B(n386), .Z(n385) );
  XNOR U280 ( .A(n387), .B(n388), .Z(n386) );
  AND U281 ( .A(o[6]), .B(n389), .Z(n387) );
  XOR U282 ( .A(n388), .B(n390), .Z(n389) );
  XOR U283 ( .A(n391), .B(n392), .Z(n383) );
  AND U284 ( .A(o[6]), .B(n393), .Z(n392) );
  XOR U285 ( .A(n391), .B(n394), .Z(n393) );
  XOR U286 ( .A(n395), .B(n396), .Z(o[2]) );
  AND U287 ( .A(o[3]), .B(n397), .Z(n396) );
  XNOR U288 ( .A(n398), .B(n399), .Z(n397) );
  XNOR U289 ( .A(n400), .B(n395), .Z(n399) );
  AND U290 ( .A(o[4]), .B(n401), .Z(n400) );
  XNOR U291 ( .A(n402), .B(n403), .Z(n401) );
  XNOR U292 ( .A(n404), .B(n398), .Z(n403) );
  AND U293 ( .A(o[5]), .B(n405), .Z(n404) );
  XNOR U294 ( .A(n402), .B(n406), .Z(n405) );
  XNOR U295 ( .A(n407), .B(n408), .Z(n406) );
  AND U296 ( .A(o[6]), .B(n409), .Z(n407) );
  XOR U297 ( .A(n408), .B(n410), .Z(n409) );
  XOR U298 ( .A(n411), .B(n412), .Z(n402) );
  AND U299 ( .A(o[6]), .B(n413), .Z(n412) );
  XOR U300 ( .A(n411), .B(n414), .Z(n413) );
  XOR U301 ( .A(n415), .B(n416), .Z(n398) );
  AND U302 ( .A(o[5]), .B(n417), .Z(n416) );
  XNOR U303 ( .A(n415), .B(n418), .Z(n417) );
  XNOR U304 ( .A(n419), .B(n420), .Z(n418) );
  AND U305 ( .A(o[6]), .B(n421), .Z(n419) );
  XOR U306 ( .A(n420), .B(n422), .Z(n421) );
  XOR U307 ( .A(n423), .B(n424), .Z(n415) );
  AND U308 ( .A(o[6]), .B(n425), .Z(n424) );
  XOR U309 ( .A(n423), .B(n426), .Z(n425) );
  XOR U310 ( .A(n427), .B(n428), .Z(n395) );
  AND U311 ( .A(o[4]), .B(n429), .Z(n428) );
  XNOR U312 ( .A(n430), .B(n431), .Z(n429) );
  XNOR U313 ( .A(n432), .B(n427), .Z(n431) );
  AND U314 ( .A(o[5]), .B(n433), .Z(n432) );
  XNOR U315 ( .A(n430), .B(n434), .Z(n433) );
  XNOR U316 ( .A(n435), .B(n436), .Z(n434) );
  AND U317 ( .A(o[6]), .B(n437), .Z(n435) );
  XOR U318 ( .A(n436), .B(n438), .Z(n437) );
  XOR U319 ( .A(n439), .B(n440), .Z(n430) );
  AND U320 ( .A(o[6]), .B(n441), .Z(n440) );
  XOR U321 ( .A(n439), .B(n442), .Z(n441) );
  XOR U322 ( .A(n443), .B(n444), .Z(n427) );
  AND U323 ( .A(o[5]), .B(n445), .Z(n444) );
  XNOR U324 ( .A(n443), .B(n446), .Z(n445) );
  XNOR U325 ( .A(n447), .B(n448), .Z(n446) );
  AND U326 ( .A(o[6]), .B(n449), .Z(n447) );
  XOR U327 ( .A(n448), .B(n450), .Z(n449) );
  XOR U328 ( .A(n451), .B(n452), .Z(n443) );
  AND U329 ( .A(o[6]), .B(n453), .Z(n452) );
  XOR U330 ( .A(n451), .B(n454), .Z(n453) );
  XOR U331 ( .A(n455), .B(n456), .Z(n331) );
  AND U332 ( .A(o[3]), .B(n457), .Z(n456) );
  XNOR U333 ( .A(n458), .B(n459), .Z(n457) );
  XNOR U334 ( .A(n460), .B(n455), .Z(n459) );
  AND U335 ( .A(o[4]), .B(n461), .Z(n460) );
  XNOR U336 ( .A(n462), .B(n463), .Z(n461) );
  XNOR U337 ( .A(n464), .B(n458), .Z(n463) );
  AND U338 ( .A(o[5]), .B(n465), .Z(n464) );
  XNOR U339 ( .A(n462), .B(n466), .Z(n465) );
  XNOR U340 ( .A(n467), .B(n468), .Z(n466) );
  AND U341 ( .A(o[6]), .B(n469), .Z(n467) );
  XOR U342 ( .A(n468), .B(n470), .Z(n469) );
  XOR U343 ( .A(n471), .B(n472), .Z(n462) );
  AND U344 ( .A(o[6]), .B(n473), .Z(n472) );
  XOR U345 ( .A(n471), .B(n474), .Z(n473) );
  XOR U346 ( .A(n475), .B(n476), .Z(n458) );
  AND U347 ( .A(o[5]), .B(n477), .Z(n476) );
  XNOR U348 ( .A(n475), .B(n478), .Z(n477) );
  XNOR U349 ( .A(n479), .B(n480), .Z(n478) );
  AND U350 ( .A(o[6]), .B(n481), .Z(n479) );
  XOR U351 ( .A(n480), .B(n482), .Z(n481) );
  XOR U352 ( .A(n483), .B(n484), .Z(n475) );
  AND U353 ( .A(o[6]), .B(n485), .Z(n484) );
  XOR U354 ( .A(n483), .B(n486), .Z(n485) );
  XOR U355 ( .A(n487), .B(n488), .Z(o[3]) );
  AND U356 ( .A(o[4]), .B(n489), .Z(n488) );
  XNOR U357 ( .A(n490), .B(n491), .Z(n489) );
  XNOR U358 ( .A(n492), .B(n487), .Z(n491) );
  AND U359 ( .A(o[5]), .B(n493), .Z(n492) );
  XNOR U360 ( .A(n490), .B(n494), .Z(n493) );
  XNOR U361 ( .A(n495), .B(n496), .Z(n494) );
  AND U362 ( .A(o[6]), .B(n497), .Z(n495) );
  XOR U363 ( .A(n496), .B(n498), .Z(n497) );
  XOR U364 ( .A(n499), .B(n500), .Z(n490) );
  AND U365 ( .A(o[6]), .B(n501), .Z(n500) );
  XOR U366 ( .A(n499), .B(n502), .Z(n501) );
  XOR U367 ( .A(n503), .B(n504), .Z(n487) );
  AND U368 ( .A(o[5]), .B(n505), .Z(n504) );
  XNOR U369 ( .A(n503), .B(n506), .Z(n505) );
  XNOR U370 ( .A(n507), .B(n508), .Z(n506) );
  AND U371 ( .A(o[6]), .B(n509), .Z(n507) );
  XOR U372 ( .A(n508), .B(n510), .Z(n509) );
  XOR U373 ( .A(n511), .B(n512), .Z(n503) );
  AND U374 ( .A(o[6]), .B(n513), .Z(n512) );
  XOR U375 ( .A(n511), .B(n514), .Z(n513) );
  XOR U376 ( .A(n515), .B(n516), .Z(n455) );
  AND U377 ( .A(o[4]), .B(n517), .Z(n516) );
  XNOR U378 ( .A(n518), .B(n519), .Z(n517) );
  XNOR U379 ( .A(n520), .B(n515), .Z(n519) );
  AND U380 ( .A(o[5]), .B(n521), .Z(n520) );
  XNOR U381 ( .A(n518), .B(n522), .Z(n521) );
  XNOR U382 ( .A(n523), .B(n524), .Z(n522) );
  AND U383 ( .A(o[6]), .B(n525), .Z(n523) );
  XOR U384 ( .A(n524), .B(n526), .Z(n525) );
  XOR U385 ( .A(n527), .B(n528), .Z(n518) );
  AND U386 ( .A(o[6]), .B(n529), .Z(n528) );
  XOR U387 ( .A(n527), .B(n530), .Z(n529) );
  XOR U388 ( .A(n531), .B(n532), .Z(o[4]) );
  AND U389 ( .A(o[5]), .B(n533), .Z(n532) );
  XNOR U390 ( .A(n531), .B(n534), .Z(n533) );
  XNOR U391 ( .A(n535), .B(n536), .Z(n534) );
  AND U392 ( .A(o[6]), .B(n537), .Z(n535) );
  XOR U393 ( .A(n536), .B(n538), .Z(n537) );
  XOR U394 ( .A(n539), .B(n540), .Z(n531) );
  AND U395 ( .A(o[6]), .B(n541), .Z(n540) );
  XOR U396 ( .A(n539), .B(n542), .Z(n541) );
  XOR U397 ( .A(n543), .B(n544), .Z(n515) );
  AND U398 ( .A(o[5]), .B(n545), .Z(n544) );
  XNOR U399 ( .A(n543), .B(n546), .Z(n545) );
  XNOR U400 ( .A(n547), .B(n548), .Z(n546) );
  AND U401 ( .A(o[6]), .B(n549), .Z(n547) );
  XOR U402 ( .A(n548), .B(n550), .Z(n549) );
  XOR U403 ( .A(n551), .B(n552), .Z(o[5]) );
  AND U404 ( .A(o[6]), .B(n553), .Z(n552) );
  XOR U405 ( .A(n551), .B(n554), .Z(n553) );
  XOR U406 ( .A(n555), .B(n556), .Z(n543) );
  AND U407 ( .A(o[6]), .B(n557), .Z(n556) );
  XOR U408 ( .A(n555), .B(n558), .Z(n557) );
  XOR U409 ( .A(n559), .B(n560), .Z(o[6]) );
  AND U410 ( .A(n561), .B(n562), .Z(n560) );
  XOR U411 ( .A(n559), .B(n17), .Z(n562) );
  XOR U412 ( .A(n563), .B(n564), .Z(n17) );
  AND U413 ( .A(n554), .B(n565), .Z(n564) );
  XOR U414 ( .A(n566), .B(n563), .Z(n565) );
  XNOR U415 ( .A(n18), .B(n559), .Z(n561) );
  IV U416 ( .A(n15), .Z(n18) );
  XNOR U417 ( .A(n567), .B(n568), .Z(n15) );
  AND U418 ( .A(n551), .B(n569), .Z(n568) );
  XOR U419 ( .A(n570), .B(n567), .Z(n569) );
  XOR U420 ( .A(n571), .B(n572), .Z(n559) );
  AND U421 ( .A(n573), .B(n574), .Z(n572) );
  XOR U422 ( .A(n571), .B(n22), .Z(n574) );
  XOR U423 ( .A(n575), .B(n576), .Z(n22) );
  AND U424 ( .A(n554), .B(n577), .Z(n576) );
  XOR U425 ( .A(n578), .B(n575), .Z(n577) );
  XNOR U426 ( .A(n23), .B(n571), .Z(n573) );
  IV U427 ( .A(n20), .Z(n23) );
  XNOR U428 ( .A(n579), .B(n580), .Z(n20) );
  AND U429 ( .A(n551), .B(n581), .Z(n580) );
  XOR U430 ( .A(n582), .B(n579), .Z(n581) );
  XOR U431 ( .A(n583), .B(n584), .Z(n571) );
  AND U432 ( .A(n585), .B(n586), .Z(n584) );
  XOR U433 ( .A(n583), .B(n27), .Z(n586) );
  XOR U434 ( .A(n587), .B(n588), .Z(n27) );
  AND U435 ( .A(n554), .B(n589), .Z(n588) );
  XOR U436 ( .A(n590), .B(n587), .Z(n589) );
  XNOR U437 ( .A(n28), .B(n583), .Z(n585) );
  IV U438 ( .A(n25), .Z(n28) );
  XNOR U439 ( .A(n591), .B(n592), .Z(n25) );
  AND U440 ( .A(n551), .B(n593), .Z(n592) );
  XOR U441 ( .A(n594), .B(n591), .Z(n593) );
  XOR U442 ( .A(n595), .B(n596), .Z(n583) );
  AND U443 ( .A(n597), .B(n598), .Z(n596) );
  XOR U444 ( .A(n595), .B(n32), .Z(n598) );
  XOR U445 ( .A(n599), .B(n600), .Z(n32) );
  AND U446 ( .A(n554), .B(n601), .Z(n600) );
  XOR U447 ( .A(n602), .B(n599), .Z(n601) );
  XNOR U448 ( .A(n33), .B(n595), .Z(n597) );
  IV U449 ( .A(n30), .Z(n33) );
  XNOR U450 ( .A(n603), .B(n604), .Z(n30) );
  AND U451 ( .A(n551), .B(n605), .Z(n604) );
  XOR U452 ( .A(n606), .B(n603), .Z(n605) );
  XOR U453 ( .A(n607), .B(n608), .Z(n595) );
  AND U454 ( .A(n609), .B(n610), .Z(n608) );
  XOR U455 ( .A(n607), .B(n37), .Z(n610) );
  XOR U456 ( .A(n611), .B(n612), .Z(n37) );
  AND U457 ( .A(n554), .B(n613), .Z(n612) );
  XOR U458 ( .A(n614), .B(n611), .Z(n613) );
  XNOR U459 ( .A(n38), .B(n607), .Z(n609) );
  IV U460 ( .A(n35), .Z(n38) );
  XNOR U461 ( .A(n615), .B(n616), .Z(n35) );
  AND U462 ( .A(n551), .B(n617), .Z(n616) );
  XOR U463 ( .A(n618), .B(n615), .Z(n617) );
  XOR U464 ( .A(n619), .B(n620), .Z(n607) );
  AND U465 ( .A(n621), .B(n622), .Z(n620) );
  XOR U466 ( .A(n619), .B(n42), .Z(n622) );
  XOR U467 ( .A(n623), .B(n624), .Z(n42) );
  AND U468 ( .A(n554), .B(n625), .Z(n624) );
  XOR U469 ( .A(n626), .B(n623), .Z(n625) );
  XNOR U470 ( .A(n43), .B(n619), .Z(n621) );
  IV U471 ( .A(n40), .Z(n43) );
  XNOR U472 ( .A(n627), .B(n628), .Z(n40) );
  AND U473 ( .A(n551), .B(n629), .Z(n628) );
  XOR U474 ( .A(n630), .B(n627), .Z(n629) );
  XOR U475 ( .A(n631), .B(n632), .Z(n619) );
  AND U476 ( .A(n633), .B(n634), .Z(n632) );
  XOR U477 ( .A(n631), .B(n47), .Z(n634) );
  XOR U478 ( .A(n635), .B(n636), .Z(n47) );
  AND U479 ( .A(n554), .B(n637), .Z(n636) );
  XOR U480 ( .A(n638), .B(n635), .Z(n637) );
  XNOR U481 ( .A(n48), .B(n631), .Z(n633) );
  IV U482 ( .A(n45), .Z(n48) );
  XNOR U483 ( .A(n639), .B(n640), .Z(n45) );
  AND U484 ( .A(n551), .B(n641), .Z(n640) );
  XOR U485 ( .A(n642), .B(n639), .Z(n641) );
  XOR U486 ( .A(n643), .B(n644), .Z(n631) );
  AND U487 ( .A(n645), .B(n646), .Z(n644) );
  XOR U488 ( .A(n643), .B(n52), .Z(n646) );
  XOR U489 ( .A(n647), .B(n648), .Z(n52) );
  AND U490 ( .A(n554), .B(n649), .Z(n648) );
  XOR U491 ( .A(n650), .B(n647), .Z(n649) );
  XNOR U492 ( .A(n53), .B(n643), .Z(n645) );
  IV U493 ( .A(n50), .Z(n53) );
  XNOR U494 ( .A(n651), .B(n652), .Z(n50) );
  AND U495 ( .A(n551), .B(n653), .Z(n652) );
  XOR U496 ( .A(n654), .B(n651), .Z(n653) );
  XOR U497 ( .A(n655), .B(n656), .Z(n643) );
  AND U498 ( .A(n657), .B(n658), .Z(n656) );
  XOR U499 ( .A(n655), .B(n57), .Z(n658) );
  XOR U500 ( .A(n659), .B(n660), .Z(n57) );
  AND U501 ( .A(n554), .B(n661), .Z(n660) );
  XOR U502 ( .A(n662), .B(n659), .Z(n661) );
  XNOR U503 ( .A(n58), .B(n655), .Z(n657) );
  IV U504 ( .A(n55), .Z(n58) );
  XNOR U505 ( .A(n663), .B(n664), .Z(n55) );
  AND U506 ( .A(n551), .B(n665), .Z(n664) );
  XOR U507 ( .A(n666), .B(n663), .Z(n665) );
  XOR U508 ( .A(n667), .B(n668), .Z(n655) );
  AND U509 ( .A(n669), .B(n670), .Z(n668) );
  XOR U510 ( .A(n667), .B(n62), .Z(n670) );
  XOR U511 ( .A(n671), .B(n672), .Z(n62) );
  AND U512 ( .A(n554), .B(n673), .Z(n672) );
  XOR U513 ( .A(n674), .B(n671), .Z(n673) );
  XNOR U514 ( .A(n63), .B(n667), .Z(n669) );
  IV U515 ( .A(n60), .Z(n63) );
  XNOR U516 ( .A(n675), .B(n676), .Z(n60) );
  AND U517 ( .A(n551), .B(n677), .Z(n676) );
  XOR U518 ( .A(n678), .B(n675), .Z(n677) );
  XOR U519 ( .A(n679), .B(n680), .Z(n667) );
  AND U520 ( .A(n681), .B(n682), .Z(n680) );
  XOR U521 ( .A(n679), .B(n67), .Z(n682) );
  XOR U522 ( .A(n683), .B(n684), .Z(n67) );
  AND U523 ( .A(n554), .B(n685), .Z(n684) );
  XOR U524 ( .A(n686), .B(n683), .Z(n685) );
  XNOR U525 ( .A(n68), .B(n679), .Z(n681) );
  IV U526 ( .A(n65), .Z(n68) );
  XNOR U527 ( .A(n687), .B(n688), .Z(n65) );
  AND U528 ( .A(n551), .B(n689), .Z(n688) );
  XOR U529 ( .A(n690), .B(n687), .Z(n689) );
  XOR U530 ( .A(n691), .B(n692), .Z(n679) );
  AND U531 ( .A(n693), .B(n694), .Z(n692) );
  XOR U532 ( .A(n691), .B(n72), .Z(n694) );
  XOR U533 ( .A(n695), .B(n696), .Z(n72) );
  AND U534 ( .A(n554), .B(n697), .Z(n696) );
  XOR U535 ( .A(n698), .B(n695), .Z(n697) );
  XNOR U536 ( .A(n73), .B(n691), .Z(n693) );
  IV U537 ( .A(n70), .Z(n73) );
  XNOR U538 ( .A(n699), .B(n700), .Z(n70) );
  AND U539 ( .A(n551), .B(n701), .Z(n700) );
  XOR U540 ( .A(n702), .B(n699), .Z(n701) );
  XOR U541 ( .A(n703), .B(n704), .Z(n691) );
  AND U542 ( .A(n705), .B(n706), .Z(n704) );
  XOR U543 ( .A(n703), .B(n77), .Z(n706) );
  XOR U544 ( .A(n707), .B(n708), .Z(n77) );
  AND U545 ( .A(n554), .B(n709), .Z(n708) );
  XOR U546 ( .A(n710), .B(n707), .Z(n709) );
  XNOR U547 ( .A(n78), .B(n703), .Z(n705) );
  IV U548 ( .A(n75), .Z(n78) );
  XNOR U549 ( .A(n711), .B(n712), .Z(n75) );
  AND U550 ( .A(n551), .B(n713), .Z(n712) );
  XOR U551 ( .A(n714), .B(n711), .Z(n713) );
  XOR U552 ( .A(n715), .B(n716), .Z(n703) );
  AND U553 ( .A(n717), .B(n718), .Z(n716) );
  XOR U554 ( .A(n4), .B(n715), .Z(n718) );
  XOR U555 ( .A(n719), .B(n720), .Z(n4) );
  AND U556 ( .A(n554), .B(n721), .Z(n720) );
  XOR U557 ( .A(n719), .B(n722), .Z(n721) );
  XNOR U558 ( .A(n715), .B(n2), .Z(n717) );
  XOR U559 ( .A(n723), .B(n724), .Z(n2) );
  AND U560 ( .A(n551), .B(n725), .Z(n724) );
  XOR U561 ( .A(n723), .B(n726), .Z(n725) );
  XNOR U562 ( .A(n727), .B(n728), .Z(n715) );
  AND U563 ( .A(n729), .B(n730), .Z(n728) );
  XNOR U564 ( .A(n727), .B(n8), .Z(n730) );
  XOR U565 ( .A(n731), .B(n732), .Z(n8) );
  AND U566 ( .A(n554), .B(n733), .Z(n732) );
  XOR U567 ( .A(n734), .B(n731), .Z(n733) );
  XOR U568 ( .A(n9), .B(n727), .Z(n729) );
  IV U569 ( .A(n6), .Z(n9) );
  XNOR U570 ( .A(n735), .B(n736), .Z(n6) );
  AND U571 ( .A(n551), .B(n737), .Z(n736) );
  XOR U572 ( .A(n738), .B(n735), .Z(n737) );
  AND U573 ( .A(n11), .B(n13), .Z(n727) );
  XNOR U574 ( .A(n739), .B(n740), .Z(n13) );
  AND U575 ( .A(n554), .B(n741), .Z(n740) );
  XNOR U576 ( .A(n742), .B(n739), .Z(n741) );
  XOR U577 ( .A(n743), .B(n744), .Z(n554) );
  AND U578 ( .A(n745), .B(n746), .Z(n744) );
  XOR U579 ( .A(n743), .B(n566), .Z(n746) );
  XOR U580 ( .A(n747), .B(n748), .Z(n566) );
  AND U581 ( .A(n538), .B(n749), .Z(n748) );
  XOR U582 ( .A(n750), .B(n747), .Z(n749) );
  XNOR U583 ( .A(n563), .B(n743), .Z(n745) );
  XOR U584 ( .A(n751), .B(n752), .Z(n563) );
  AND U585 ( .A(n536), .B(n753), .Z(n752) );
  XOR U586 ( .A(n754), .B(n751), .Z(n753) );
  XOR U587 ( .A(n755), .B(n756), .Z(n743) );
  AND U588 ( .A(n757), .B(n758), .Z(n756) );
  XOR U589 ( .A(n755), .B(n578), .Z(n758) );
  XOR U590 ( .A(n759), .B(n760), .Z(n578) );
  AND U591 ( .A(n538), .B(n761), .Z(n760) );
  XOR U592 ( .A(n762), .B(n759), .Z(n761) );
  XNOR U593 ( .A(n575), .B(n755), .Z(n757) );
  XOR U594 ( .A(n763), .B(n764), .Z(n575) );
  AND U595 ( .A(n536), .B(n765), .Z(n764) );
  XOR U596 ( .A(n766), .B(n763), .Z(n765) );
  XOR U597 ( .A(n767), .B(n768), .Z(n755) );
  AND U598 ( .A(n769), .B(n770), .Z(n768) );
  XOR U599 ( .A(n767), .B(n590), .Z(n770) );
  XOR U600 ( .A(n771), .B(n772), .Z(n590) );
  AND U601 ( .A(n538), .B(n773), .Z(n772) );
  XOR U602 ( .A(n774), .B(n771), .Z(n773) );
  XNOR U603 ( .A(n587), .B(n767), .Z(n769) );
  XOR U604 ( .A(n775), .B(n776), .Z(n587) );
  AND U605 ( .A(n536), .B(n777), .Z(n776) );
  XOR U606 ( .A(n778), .B(n775), .Z(n777) );
  XOR U607 ( .A(n779), .B(n780), .Z(n767) );
  AND U608 ( .A(n781), .B(n782), .Z(n780) );
  XOR U609 ( .A(n779), .B(n602), .Z(n782) );
  XOR U610 ( .A(n783), .B(n784), .Z(n602) );
  AND U611 ( .A(n538), .B(n785), .Z(n784) );
  XOR U612 ( .A(n786), .B(n783), .Z(n785) );
  XNOR U613 ( .A(n599), .B(n779), .Z(n781) );
  XOR U614 ( .A(n787), .B(n788), .Z(n599) );
  AND U615 ( .A(n536), .B(n789), .Z(n788) );
  XOR U616 ( .A(n790), .B(n787), .Z(n789) );
  XOR U617 ( .A(n791), .B(n792), .Z(n779) );
  AND U618 ( .A(n793), .B(n794), .Z(n792) );
  XOR U619 ( .A(n791), .B(n614), .Z(n794) );
  XOR U620 ( .A(n795), .B(n796), .Z(n614) );
  AND U621 ( .A(n538), .B(n797), .Z(n796) );
  XOR U622 ( .A(n798), .B(n795), .Z(n797) );
  XNOR U623 ( .A(n611), .B(n791), .Z(n793) );
  XOR U624 ( .A(n799), .B(n800), .Z(n611) );
  AND U625 ( .A(n536), .B(n801), .Z(n800) );
  XOR U626 ( .A(n802), .B(n799), .Z(n801) );
  XOR U627 ( .A(n803), .B(n804), .Z(n791) );
  AND U628 ( .A(n805), .B(n806), .Z(n804) );
  XOR U629 ( .A(n803), .B(n626), .Z(n806) );
  XOR U630 ( .A(n807), .B(n808), .Z(n626) );
  AND U631 ( .A(n538), .B(n809), .Z(n808) );
  XOR U632 ( .A(n810), .B(n807), .Z(n809) );
  XNOR U633 ( .A(n623), .B(n803), .Z(n805) );
  XOR U634 ( .A(n811), .B(n812), .Z(n623) );
  AND U635 ( .A(n536), .B(n813), .Z(n812) );
  XOR U636 ( .A(n814), .B(n811), .Z(n813) );
  XOR U637 ( .A(n815), .B(n816), .Z(n803) );
  AND U638 ( .A(n817), .B(n818), .Z(n816) );
  XOR U639 ( .A(n815), .B(n638), .Z(n818) );
  XOR U640 ( .A(n819), .B(n820), .Z(n638) );
  AND U641 ( .A(n538), .B(n821), .Z(n820) );
  XOR U642 ( .A(n822), .B(n819), .Z(n821) );
  XNOR U643 ( .A(n635), .B(n815), .Z(n817) );
  XOR U644 ( .A(n823), .B(n824), .Z(n635) );
  AND U645 ( .A(n536), .B(n825), .Z(n824) );
  XOR U646 ( .A(n826), .B(n823), .Z(n825) );
  XOR U647 ( .A(n827), .B(n828), .Z(n815) );
  AND U648 ( .A(n829), .B(n830), .Z(n828) );
  XOR U649 ( .A(n827), .B(n650), .Z(n830) );
  XOR U650 ( .A(n831), .B(n832), .Z(n650) );
  AND U651 ( .A(n538), .B(n833), .Z(n832) );
  XOR U652 ( .A(n834), .B(n831), .Z(n833) );
  XNOR U653 ( .A(n647), .B(n827), .Z(n829) );
  XOR U654 ( .A(n835), .B(n836), .Z(n647) );
  AND U655 ( .A(n536), .B(n837), .Z(n836) );
  XOR U656 ( .A(n838), .B(n835), .Z(n837) );
  XOR U657 ( .A(n839), .B(n840), .Z(n827) );
  AND U658 ( .A(n841), .B(n842), .Z(n840) );
  XOR U659 ( .A(n839), .B(n662), .Z(n842) );
  XOR U660 ( .A(n843), .B(n844), .Z(n662) );
  AND U661 ( .A(n538), .B(n845), .Z(n844) );
  XOR U662 ( .A(n846), .B(n843), .Z(n845) );
  XNOR U663 ( .A(n659), .B(n839), .Z(n841) );
  XOR U664 ( .A(n847), .B(n848), .Z(n659) );
  AND U665 ( .A(n536), .B(n849), .Z(n848) );
  XOR U666 ( .A(n850), .B(n847), .Z(n849) );
  XOR U667 ( .A(n851), .B(n852), .Z(n839) );
  AND U668 ( .A(n853), .B(n854), .Z(n852) );
  XOR U669 ( .A(n851), .B(n674), .Z(n854) );
  XOR U670 ( .A(n855), .B(n856), .Z(n674) );
  AND U671 ( .A(n538), .B(n857), .Z(n856) );
  XOR U672 ( .A(n858), .B(n855), .Z(n857) );
  XNOR U673 ( .A(n671), .B(n851), .Z(n853) );
  XOR U674 ( .A(n859), .B(n860), .Z(n671) );
  AND U675 ( .A(n536), .B(n861), .Z(n860) );
  XOR U676 ( .A(n862), .B(n859), .Z(n861) );
  XOR U677 ( .A(n863), .B(n864), .Z(n851) );
  AND U678 ( .A(n865), .B(n866), .Z(n864) );
  XOR U679 ( .A(n863), .B(n686), .Z(n866) );
  XOR U680 ( .A(n867), .B(n868), .Z(n686) );
  AND U681 ( .A(n538), .B(n869), .Z(n868) );
  XOR U682 ( .A(n870), .B(n867), .Z(n869) );
  XNOR U683 ( .A(n683), .B(n863), .Z(n865) );
  XOR U684 ( .A(n871), .B(n872), .Z(n683) );
  AND U685 ( .A(n536), .B(n873), .Z(n872) );
  XOR U686 ( .A(n874), .B(n871), .Z(n873) );
  XOR U687 ( .A(n875), .B(n876), .Z(n863) );
  AND U688 ( .A(n877), .B(n878), .Z(n876) );
  XOR U689 ( .A(n875), .B(n698), .Z(n878) );
  XOR U690 ( .A(n879), .B(n880), .Z(n698) );
  AND U691 ( .A(n538), .B(n881), .Z(n880) );
  XOR U692 ( .A(n882), .B(n879), .Z(n881) );
  XNOR U693 ( .A(n695), .B(n875), .Z(n877) );
  XOR U694 ( .A(n883), .B(n884), .Z(n695) );
  AND U695 ( .A(n536), .B(n885), .Z(n884) );
  XOR U696 ( .A(n886), .B(n883), .Z(n885) );
  XOR U697 ( .A(n887), .B(n888), .Z(n875) );
  AND U698 ( .A(n889), .B(n890), .Z(n888) );
  XOR U699 ( .A(n887), .B(n710), .Z(n890) );
  XOR U700 ( .A(n891), .B(n892), .Z(n710) );
  AND U701 ( .A(n538), .B(n893), .Z(n892) );
  XOR U702 ( .A(n894), .B(n891), .Z(n893) );
  XNOR U703 ( .A(n707), .B(n887), .Z(n889) );
  XOR U704 ( .A(n895), .B(n896), .Z(n707) );
  AND U705 ( .A(n536), .B(n897), .Z(n896) );
  XOR U706 ( .A(n898), .B(n895), .Z(n897) );
  XOR U707 ( .A(n899), .B(n900), .Z(n887) );
  AND U708 ( .A(n901), .B(n902), .Z(n900) );
  XOR U709 ( .A(n722), .B(n899), .Z(n902) );
  XOR U710 ( .A(n903), .B(n904), .Z(n722) );
  AND U711 ( .A(n538), .B(n905), .Z(n904) );
  XOR U712 ( .A(n903), .B(n906), .Z(n905) );
  XNOR U713 ( .A(n899), .B(n719), .Z(n901) );
  XOR U714 ( .A(n907), .B(n908), .Z(n719) );
  AND U715 ( .A(n536), .B(n909), .Z(n908) );
  XOR U716 ( .A(n907), .B(n910), .Z(n909) );
  XOR U717 ( .A(n911), .B(n912), .Z(n899) );
  AND U718 ( .A(n913), .B(n914), .Z(n912) );
  XNOR U719 ( .A(n915), .B(n734), .Z(n914) );
  XOR U720 ( .A(n916), .B(n917), .Z(n734) );
  AND U721 ( .A(n538), .B(n918), .Z(n917) );
  XOR U722 ( .A(n919), .B(n916), .Z(n918) );
  XNOR U723 ( .A(n731), .B(n911), .Z(n913) );
  XOR U724 ( .A(n920), .B(n921), .Z(n731) );
  AND U725 ( .A(n536), .B(n922), .Z(n921) );
  XOR U726 ( .A(n923), .B(n920), .Z(n922) );
  IV U727 ( .A(n915), .Z(n911) );
  AND U728 ( .A(n739), .B(n742), .Z(n915) );
  XNOR U729 ( .A(n924), .B(n925), .Z(n742) );
  AND U730 ( .A(n538), .B(n926), .Z(n925) );
  XNOR U731 ( .A(n927), .B(n924), .Z(n926) );
  XOR U732 ( .A(n928), .B(n929), .Z(n538) );
  AND U733 ( .A(n930), .B(n931), .Z(n929) );
  XOR U734 ( .A(n928), .B(n750), .Z(n931) );
  XNOR U735 ( .A(n932), .B(n933), .Z(n750) );
  AND U736 ( .A(n934), .B(n498), .Z(n933) );
  AND U737 ( .A(n932), .B(n935), .Z(n934) );
  XNOR U738 ( .A(n747), .B(n928), .Z(n930) );
  XOR U739 ( .A(n936), .B(n937), .Z(n747) );
  AND U740 ( .A(n938), .B(n496), .Z(n937) );
  NOR U741 ( .A(n936), .B(n939), .Z(n938) );
  XOR U742 ( .A(n940), .B(n941), .Z(n928) );
  AND U743 ( .A(n942), .B(n943), .Z(n941) );
  XOR U744 ( .A(n940), .B(n762), .Z(n943) );
  XOR U745 ( .A(n944), .B(n945), .Z(n762) );
  AND U746 ( .A(n498), .B(n946), .Z(n945) );
  XOR U747 ( .A(n947), .B(n944), .Z(n946) );
  XNOR U748 ( .A(n759), .B(n940), .Z(n942) );
  XOR U749 ( .A(n948), .B(n949), .Z(n759) );
  AND U750 ( .A(n496), .B(n950), .Z(n949) );
  XOR U751 ( .A(n951), .B(n948), .Z(n950) );
  XOR U752 ( .A(n952), .B(n953), .Z(n940) );
  AND U753 ( .A(n954), .B(n955), .Z(n953) );
  XOR U754 ( .A(n952), .B(n774), .Z(n955) );
  XOR U755 ( .A(n956), .B(n957), .Z(n774) );
  AND U756 ( .A(n498), .B(n958), .Z(n957) );
  XOR U757 ( .A(n959), .B(n956), .Z(n958) );
  XNOR U758 ( .A(n771), .B(n952), .Z(n954) );
  XOR U759 ( .A(n960), .B(n961), .Z(n771) );
  AND U760 ( .A(n496), .B(n962), .Z(n961) );
  XOR U761 ( .A(n963), .B(n960), .Z(n962) );
  XOR U762 ( .A(n964), .B(n965), .Z(n952) );
  AND U763 ( .A(n966), .B(n967), .Z(n965) );
  XOR U764 ( .A(n964), .B(n786), .Z(n967) );
  XOR U765 ( .A(n968), .B(n969), .Z(n786) );
  AND U766 ( .A(n498), .B(n970), .Z(n969) );
  XOR U767 ( .A(n971), .B(n968), .Z(n970) );
  XNOR U768 ( .A(n783), .B(n964), .Z(n966) );
  XOR U769 ( .A(n972), .B(n973), .Z(n783) );
  AND U770 ( .A(n496), .B(n974), .Z(n973) );
  XOR U771 ( .A(n975), .B(n972), .Z(n974) );
  XOR U772 ( .A(n976), .B(n977), .Z(n964) );
  AND U773 ( .A(n978), .B(n979), .Z(n977) );
  XOR U774 ( .A(n976), .B(n798), .Z(n979) );
  XOR U775 ( .A(n980), .B(n981), .Z(n798) );
  AND U776 ( .A(n498), .B(n982), .Z(n981) );
  XOR U777 ( .A(n983), .B(n980), .Z(n982) );
  XNOR U778 ( .A(n795), .B(n976), .Z(n978) );
  XOR U779 ( .A(n984), .B(n985), .Z(n795) );
  AND U780 ( .A(n496), .B(n986), .Z(n985) );
  XOR U781 ( .A(n987), .B(n984), .Z(n986) );
  XOR U782 ( .A(n988), .B(n989), .Z(n976) );
  AND U783 ( .A(n990), .B(n991), .Z(n989) );
  XOR U784 ( .A(n988), .B(n810), .Z(n991) );
  XOR U785 ( .A(n992), .B(n993), .Z(n810) );
  AND U786 ( .A(n498), .B(n994), .Z(n993) );
  XOR U787 ( .A(n995), .B(n992), .Z(n994) );
  XNOR U788 ( .A(n807), .B(n988), .Z(n990) );
  XOR U789 ( .A(n996), .B(n997), .Z(n807) );
  AND U790 ( .A(n496), .B(n998), .Z(n997) );
  XOR U791 ( .A(n999), .B(n996), .Z(n998) );
  XOR U792 ( .A(n1000), .B(n1001), .Z(n988) );
  AND U793 ( .A(n1002), .B(n1003), .Z(n1001) );
  XOR U794 ( .A(n1000), .B(n822), .Z(n1003) );
  XOR U795 ( .A(n1004), .B(n1005), .Z(n822) );
  AND U796 ( .A(n498), .B(n1006), .Z(n1005) );
  XOR U797 ( .A(n1007), .B(n1004), .Z(n1006) );
  XNOR U798 ( .A(n819), .B(n1000), .Z(n1002) );
  XOR U799 ( .A(n1008), .B(n1009), .Z(n819) );
  AND U800 ( .A(n496), .B(n1010), .Z(n1009) );
  XOR U801 ( .A(n1011), .B(n1008), .Z(n1010) );
  XOR U802 ( .A(n1012), .B(n1013), .Z(n1000) );
  AND U803 ( .A(n1014), .B(n1015), .Z(n1013) );
  XOR U804 ( .A(n1012), .B(n834), .Z(n1015) );
  XOR U805 ( .A(n1016), .B(n1017), .Z(n834) );
  AND U806 ( .A(n498), .B(n1018), .Z(n1017) );
  XOR U807 ( .A(n1019), .B(n1016), .Z(n1018) );
  XNOR U808 ( .A(n831), .B(n1012), .Z(n1014) );
  XOR U809 ( .A(n1020), .B(n1021), .Z(n831) );
  AND U810 ( .A(n496), .B(n1022), .Z(n1021) );
  XOR U811 ( .A(n1023), .B(n1020), .Z(n1022) );
  XOR U812 ( .A(n1024), .B(n1025), .Z(n1012) );
  AND U813 ( .A(n1026), .B(n1027), .Z(n1025) );
  XOR U814 ( .A(n1024), .B(n846), .Z(n1027) );
  XOR U815 ( .A(n1028), .B(n1029), .Z(n846) );
  AND U816 ( .A(n498), .B(n1030), .Z(n1029) );
  XOR U817 ( .A(n1031), .B(n1028), .Z(n1030) );
  XNOR U818 ( .A(n843), .B(n1024), .Z(n1026) );
  XOR U819 ( .A(n1032), .B(n1033), .Z(n843) );
  AND U820 ( .A(n496), .B(n1034), .Z(n1033) );
  XOR U821 ( .A(n1035), .B(n1032), .Z(n1034) );
  XOR U822 ( .A(n1036), .B(n1037), .Z(n1024) );
  AND U823 ( .A(n1038), .B(n1039), .Z(n1037) );
  XOR U824 ( .A(n1036), .B(n858), .Z(n1039) );
  XOR U825 ( .A(n1040), .B(n1041), .Z(n858) );
  AND U826 ( .A(n498), .B(n1042), .Z(n1041) );
  XOR U827 ( .A(n1043), .B(n1040), .Z(n1042) );
  XNOR U828 ( .A(n855), .B(n1036), .Z(n1038) );
  XOR U829 ( .A(n1044), .B(n1045), .Z(n855) );
  AND U830 ( .A(n496), .B(n1046), .Z(n1045) );
  XOR U831 ( .A(n1047), .B(n1044), .Z(n1046) );
  XOR U832 ( .A(n1048), .B(n1049), .Z(n1036) );
  AND U833 ( .A(n1050), .B(n1051), .Z(n1049) );
  XOR U834 ( .A(n1048), .B(n870), .Z(n1051) );
  XOR U835 ( .A(n1052), .B(n1053), .Z(n870) );
  AND U836 ( .A(n498), .B(n1054), .Z(n1053) );
  XOR U837 ( .A(n1055), .B(n1052), .Z(n1054) );
  XNOR U838 ( .A(n867), .B(n1048), .Z(n1050) );
  XOR U839 ( .A(n1056), .B(n1057), .Z(n867) );
  AND U840 ( .A(n496), .B(n1058), .Z(n1057) );
  XOR U841 ( .A(n1059), .B(n1056), .Z(n1058) );
  XOR U842 ( .A(n1060), .B(n1061), .Z(n1048) );
  AND U843 ( .A(n1062), .B(n1063), .Z(n1061) );
  XOR U844 ( .A(n1060), .B(n882), .Z(n1063) );
  XOR U845 ( .A(n1064), .B(n1065), .Z(n882) );
  AND U846 ( .A(n498), .B(n1066), .Z(n1065) );
  XOR U847 ( .A(n1067), .B(n1064), .Z(n1066) );
  XNOR U848 ( .A(n879), .B(n1060), .Z(n1062) );
  XOR U849 ( .A(n1068), .B(n1069), .Z(n879) );
  AND U850 ( .A(n496), .B(n1070), .Z(n1069) );
  XOR U851 ( .A(n1071), .B(n1068), .Z(n1070) );
  XOR U852 ( .A(n1072), .B(n1073), .Z(n1060) );
  AND U853 ( .A(n1074), .B(n1075), .Z(n1073) );
  XOR U854 ( .A(n1072), .B(n894), .Z(n1075) );
  XOR U855 ( .A(n1076), .B(n1077), .Z(n894) );
  AND U856 ( .A(n498), .B(n1078), .Z(n1077) );
  XOR U857 ( .A(n1079), .B(n1076), .Z(n1078) );
  XNOR U858 ( .A(n891), .B(n1072), .Z(n1074) );
  XOR U859 ( .A(n1080), .B(n1081), .Z(n891) );
  AND U860 ( .A(n496), .B(n1082), .Z(n1081) );
  XOR U861 ( .A(n1083), .B(n1080), .Z(n1082) );
  XOR U862 ( .A(n1084), .B(n1085), .Z(n1072) );
  AND U863 ( .A(n1086), .B(n1087), .Z(n1085) );
  XOR U864 ( .A(n906), .B(n1084), .Z(n1087) );
  XOR U865 ( .A(n1088), .B(n1089), .Z(n906) );
  AND U866 ( .A(n498), .B(n1090), .Z(n1089) );
  XOR U867 ( .A(n1088), .B(n1091), .Z(n1090) );
  XNOR U868 ( .A(n1084), .B(n903), .Z(n1086) );
  XOR U869 ( .A(n1092), .B(n1093), .Z(n903) );
  AND U870 ( .A(n496), .B(n1094), .Z(n1093) );
  XOR U871 ( .A(n1092), .B(n1095), .Z(n1094) );
  XOR U872 ( .A(n1096), .B(n1097), .Z(n1084) );
  AND U873 ( .A(n1098), .B(n1099), .Z(n1097) );
  XNOR U874 ( .A(n1100), .B(n919), .Z(n1099) );
  XOR U875 ( .A(n1101), .B(n1102), .Z(n919) );
  AND U876 ( .A(n498), .B(n1103), .Z(n1102) );
  XOR U877 ( .A(n1104), .B(n1101), .Z(n1103) );
  XNOR U878 ( .A(n916), .B(n1096), .Z(n1098) );
  XOR U879 ( .A(n1105), .B(n1106), .Z(n916) );
  AND U880 ( .A(n496), .B(n1107), .Z(n1106) );
  XOR U881 ( .A(n1108), .B(n1105), .Z(n1107) );
  IV U882 ( .A(n1100), .Z(n1096) );
  AND U883 ( .A(n924), .B(n927), .Z(n1100) );
  XNOR U884 ( .A(n1109), .B(n1110), .Z(n927) );
  AND U885 ( .A(n498), .B(n1111), .Z(n1110) );
  XNOR U886 ( .A(n1112), .B(n1109), .Z(n1111) );
  XOR U887 ( .A(n1113), .B(n1114), .Z(n498) );
  AND U888 ( .A(n1115), .B(n1116), .Z(n1114) );
  XOR U889 ( .A(n935), .B(n1113), .Z(n1116) );
  IV U890 ( .A(n1117), .Z(n935) );
  AND U891 ( .A(n1118), .B(n1119), .Z(n1117) );
  XOR U892 ( .A(n1113), .B(n932), .Z(n1115) );
  AND U893 ( .A(n1120), .B(n1121), .Z(n932) );
  XOR U894 ( .A(n1122), .B(n1123), .Z(n1113) );
  AND U895 ( .A(n1124), .B(n1125), .Z(n1123) );
  XOR U896 ( .A(n1122), .B(n947), .Z(n1125) );
  XOR U897 ( .A(n1126), .B(n1127), .Z(n947) );
  AND U898 ( .A(n410), .B(n1128), .Z(n1127) );
  XOR U899 ( .A(n1129), .B(n1126), .Z(n1128) );
  XNOR U900 ( .A(n944), .B(n1122), .Z(n1124) );
  XOR U901 ( .A(n1130), .B(n1131), .Z(n944) );
  AND U902 ( .A(n408), .B(n1132), .Z(n1131) );
  XOR U903 ( .A(n1133), .B(n1130), .Z(n1132) );
  XOR U904 ( .A(n1134), .B(n1135), .Z(n1122) );
  AND U905 ( .A(n1136), .B(n1137), .Z(n1135) );
  XOR U906 ( .A(n1134), .B(n959), .Z(n1137) );
  XOR U907 ( .A(n1138), .B(n1139), .Z(n959) );
  AND U908 ( .A(n410), .B(n1140), .Z(n1139) );
  XOR U909 ( .A(n1141), .B(n1138), .Z(n1140) );
  XNOR U910 ( .A(n956), .B(n1134), .Z(n1136) );
  XOR U911 ( .A(n1142), .B(n1143), .Z(n956) );
  AND U912 ( .A(n408), .B(n1144), .Z(n1143) );
  XOR U913 ( .A(n1145), .B(n1142), .Z(n1144) );
  XOR U914 ( .A(n1146), .B(n1147), .Z(n1134) );
  AND U915 ( .A(n1148), .B(n1149), .Z(n1147) );
  XOR U916 ( .A(n1146), .B(n971), .Z(n1149) );
  XOR U917 ( .A(n1150), .B(n1151), .Z(n971) );
  AND U918 ( .A(n410), .B(n1152), .Z(n1151) );
  XOR U919 ( .A(n1153), .B(n1150), .Z(n1152) );
  XNOR U920 ( .A(n968), .B(n1146), .Z(n1148) );
  XOR U921 ( .A(n1154), .B(n1155), .Z(n968) );
  AND U922 ( .A(n408), .B(n1156), .Z(n1155) );
  XOR U923 ( .A(n1157), .B(n1154), .Z(n1156) );
  XOR U924 ( .A(n1158), .B(n1159), .Z(n1146) );
  AND U925 ( .A(n1160), .B(n1161), .Z(n1159) );
  XOR U926 ( .A(n1158), .B(n983), .Z(n1161) );
  XOR U927 ( .A(n1162), .B(n1163), .Z(n983) );
  AND U928 ( .A(n410), .B(n1164), .Z(n1163) );
  XOR U929 ( .A(n1165), .B(n1162), .Z(n1164) );
  XNOR U930 ( .A(n980), .B(n1158), .Z(n1160) );
  XOR U931 ( .A(n1166), .B(n1167), .Z(n980) );
  AND U932 ( .A(n408), .B(n1168), .Z(n1167) );
  XOR U933 ( .A(n1169), .B(n1166), .Z(n1168) );
  XOR U934 ( .A(n1170), .B(n1171), .Z(n1158) );
  AND U935 ( .A(n1172), .B(n1173), .Z(n1171) );
  XOR U936 ( .A(n1170), .B(n995), .Z(n1173) );
  XOR U937 ( .A(n1174), .B(n1175), .Z(n995) );
  AND U938 ( .A(n410), .B(n1176), .Z(n1175) );
  XOR U939 ( .A(n1177), .B(n1174), .Z(n1176) );
  XNOR U940 ( .A(n992), .B(n1170), .Z(n1172) );
  XOR U941 ( .A(n1178), .B(n1179), .Z(n992) );
  AND U942 ( .A(n408), .B(n1180), .Z(n1179) );
  XOR U943 ( .A(n1181), .B(n1178), .Z(n1180) );
  XOR U944 ( .A(n1182), .B(n1183), .Z(n1170) );
  AND U945 ( .A(n1184), .B(n1185), .Z(n1183) );
  XOR U946 ( .A(n1182), .B(n1007), .Z(n1185) );
  XOR U947 ( .A(n1186), .B(n1187), .Z(n1007) );
  AND U948 ( .A(n410), .B(n1188), .Z(n1187) );
  XOR U949 ( .A(n1189), .B(n1186), .Z(n1188) );
  XNOR U950 ( .A(n1004), .B(n1182), .Z(n1184) );
  XOR U951 ( .A(n1190), .B(n1191), .Z(n1004) );
  AND U952 ( .A(n408), .B(n1192), .Z(n1191) );
  XOR U953 ( .A(n1193), .B(n1190), .Z(n1192) );
  XOR U954 ( .A(n1194), .B(n1195), .Z(n1182) );
  AND U955 ( .A(n1196), .B(n1197), .Z(n1195) );
  XOR U956 ( .A(n1194), .B(n1019), .Z(n1197) );
  XOR U957 ( .A(n1198), .B(n1199), .Z(n1019) );
  AND U958 ( .A(n410), .B(n1200), .Z(n1199) );
  XOR U959 ( .A(n1201), .B(n1198), .Z(n1200) );
  XNOR U960 ( .A(n1016), .B(n1194), .Z(n1196) );
  XOR U961 ( .A(n1202), .B(n1203), .Z(n1016) );
  AND U962 ( .A(n408), .B(n1204), .Z(n1203) );
  XOR U963 ( .A(n1205), .B(n1202), .Z(n1204) );
  XOR U964 ( .A(n1206), .B(n1207), .Z(n1194) );
  AND U965 ( .A(n1208), .B(n1209), .Z(n1207) );
  XOR U966 ( .A(n1206), .B(n1031), .Z(n1209) );
  XOR U967 ( .A(n1210), .B(n1211), .Z(n1031) );
  AND U968 ( .A(n410), .B(n1212), .Z(n1211) );
  XOR U969 ( .A(n1213), .B(n1210), .Z(n1212) );
  XNOR U970 ( .A(n1028), .B(n1206), .Z(n1208) );
  XOR U971 ( .A(n1214), .B(n1215), .Z(n1028) );
  AND U972 ( .A(n408), .B(n1216), .Z(n1215) );
  XOR U973 ( .A(n1217), .B(n1214), .Z(n1216) );
  XOR U974 ( .A(n1218), .B(n1219), .Z(n1206) );
  AND U975 ( .A(n1220), .B(n1221), .Z(n1219) );
  XOR U976 ( .A(n1218), .B(n1043), .Z(n1221) );
  XOR U977 ( .A(n1222), .B(n1223), .Z(n1043) );
  AND U978 ( .A(n410), .B(n1224), .Z(n1223) );
  XOR U979 ( .A(n1225), .B(n1222), .Z(n1224) );
  XNOR U980 ( .A(n1040), .B(n1218), .Z(n1220) );
  XOR U981 ( .A(n1226), .B(n1227), .Z(n1040) );
  AND U982 ( .A(n408), .B(n1228), .Z(n1227) );
  XOR U983 ( .A(n1229), .B(n1226), .Z(n1228) );
  XOR U984 ( .A(n1230), .B(n1231), .Z(n1218) );
  AND U985 ( .A(n1232), .B(n1233), .Z(n1231) );
  XOR U986 ( .A(n1230), .B(n1055), .Z(n1233) );
  XOR U987 ( .A(n1234), .B(n1235), .Z(n1055) );
  AND U988 ( .A(n410), .B(n1236), .Z(n1235) );
  XOR U989 ( .A(n1237), .B(n1234), .Z(n1236) );
  XNOR U990 ( .A(n1052), .B(n1230), .Z(n1232) );
  XOR U991 ( .A(n1238), .B(n1239), .Z(n1052) );
  AND U992 ( .A(n408), .B(n1240), .Z(n1239) );
  XOR U993 ( .A(n1241), .B(n1238), .Z(n1240) );
  XOR U994 ( .A(n1242), .B(n1243), .Z(n1230) );
  AND U995 ( .A(n1244), .B(n1245), .Z(n1243) );
  XOR U996 ( .A(n1242), .B(n1067), .Z(n1245) );
  XOR U997 ( .A(n1246), .B(n1247), .Z(n1067) );
  AND U998 ( .A(n410), .B(n1248), .Z(n1247) );
  XOR U999 ( .A(n1249), .B(n1246), .Z(n1248) );
  XNOR U1000 ( .A(n1064), .B(n1242), .Z(n1244) );
  XOR U1001 ( .A(n1250), .B(n1251), .Z(n1064) );
  AND U1002 ( .A(n408), .B(n1252), .Z(n1251) );
  XOR U1003 ( .A(n1253), .B(n1250), .Z(n1252) );
  XOR U1004 ( .A(n1254), .B(n1255), .Z(n1242) );
  AND U1005 ( .A(n1256), .B(n1257), .Z(n1255) );
  XOR U1006 ( .A(n1254), .B(n1079), .Z(n1257) );
  XOR U1007 ( .A(n1258), .B(n1259), .Z(n1079) );
  AND U1008 ( .A(n410), .B(n1260), .Z(n1259) );
  XOR U1009 ( .A(n1261), .B(n1258), .Z(n1260) );
  XNOR U1010 ( .A(n1076), .B(n1254), .Z(n1256) );
  XOR U1011 ( .A(n1262), .B(n1263), .Z(n1076) );
  AND U1012 ( .A(n408), .B(n1264), .Z(n1263) );
  XOR U1013 ( .A(n1265), .B(n1262), .Z(n1264) );
  XOR U1014 ( .A(n1266), .B(n1267), .Z(n1254) );
  AND U1015 ( .A(n1268), .B(n1269), .Z(n1267) );
  XOR U1016 ( .A(n1091), .B(n1266), .Z(n1269) );
  XOR U1017 ( .A(n1270), .B(n1271), .Z(n1091) );
  AND U1018 ( .A(n410), .B(n1272), .Z(n1271) );
  XOR U1019 ( .A(n1270), .B(n1273), .Z(n1272) );
  XNOR U1020 ( .A(n1266), .B(n1088), .Z(n1268) );
  XOR U1021 ( .A(n1274), .B(n1275), .Z(n1088) );
  AND U1022 ( .A(n408), .B(n1276), .Z(n1275) );
  XOR U1023 ( .A(n1274), .B(n1277), .Z(n1276) );
  XOR U1024 ( .A(n1278), .B(n1279), .Z(n1266) );
  AND U1025 ( .A(n1280), .B(n1281), .Z(n1279) );
  XNOR U1026 ( .A(n1282), .B(n1104), .Z(n1281) );
  XOR U1027 ( .A(n1283), .B(n1284), .Z(n1104) );
  AND U1028 ( .A(n410), .B(n1285), .Z(n1284) );
  XOR U1029 ( .A(n1286), .B(n1283), .Z(n1285) );
  XNOR U1030 ( .A(n1101), .B(n1278), .Z(n1280) );
  XOR U1031 ( .A(n1287), .B(n1288), .Z(n1101) );
  AND U1032 ( .A(n408), .B(n1289), .Z(n1288) );
  XOR U1033 ( .A(n1290), .B(n1287), .Z(n1289) );
  IV U1034 ( .A(n1282), .Z(n1278) );
  AND U1035 ( .A(n1109), .B(n1112), .Z(n1282) );
  XNOR U1036 ( .A(n1291), .B(n1292), .Z(n1112) );
  AND U1037 ( .A(n410), .B(n1293), .Z(n1292) );
  XNOR U1038 ( .A(n1294), .B(n1291), .Z(n1293) );
  XOR U1039 ( .A(n1295), .B(n1296), .Z(n410) );
  AND U1040 ( .A(n1297), .B(n1298), .Z(n1296) );
  XNOR U1041 ( .A(n1118), .B(n1295), .Z(n1298) );
  AND U1042 ( .A(n1299), .B(n1300), .Z(n1118) );
  XOR U1043 ( .A(n1295), .B(n1119), .Z(n1297) );
  AND U1044 ( .A(n1301), .B(n1302), .Z(n1119) );
  XOR U1045 ( .A(n1303), .B(n1304), .Z(n1295) );
  AND U1046 ( .A(n1305), .B(n1306), .Z(n1304) );
  XOR U1047 ( .A(n1303), .B(n1129), .Z(n1306) );
  XOR U1048 ( .A(n1307), .B(n1308), .Z(n1129) );
  AND U1049 ( .A(n226), .B(n1309), .Z(n1308) );
  XOR U1050 ( .A(n1310), .B(n1307), .Z(n1309) );
  XNOR U1051 ( .A(n1126), .B(n1303), .Z(n1305) );
  XOR U1052 ( .A(n1311), .B(n1312), .Z(n1126) );
  AND U1053 ( .A(n224), .B(n1313), .Z(n1312) );
  XOR U1054 ( .A(n1314), .B(n1311), .Z(n1313) );
  XOR U1055 ( .A(n1315), .B(n1316), .Z(n1303) );
  AND U1056 ( .A(n1317), .B(n1318), .Z(n1316) );
  XOR U1057 ( .A(n1315), .B(n1141), .Z(n1318) );
  XOR U1058 ( .A(n1319), .B(n1320), .Z(n1141) );
  AND U1059 ( .A(n226), .B(n1321), .Z(n1320) );
  XOR U1060 ( .A(n1322), .B(n1319), .Z(n1321) );
  XNOR U1061 ( .A(n1138), .B(n1315), .Z(n1317) );
  XOR U1062 ( .A(n1323), .B(n1324), .Z(n1138) );
  AND U1063 ( .A(n224), .B(n1325), .Z(n1324) );
  XOR U1064 ( .A(n1326), .B(n1323), .Z(n1325) );
  XOR U1065 ( .A(n1327), .B(n1328), .Z(n1315) );
  AND U1066 ( .A(n1329), .B(n1330), .Z(n1328) );
  XOR U1067 ( .A(n1327), .B(n1153), .Z(n1330) );
  XOR U1068 ( .A(n1331), .B(n1332), .Z(n1153) );
  AND U1069 ( .A(n226), .B(n1333), .Z(n1332) );
  XOR U1070 ( .A(n1334), .B(n1331), .Z(n1333) );
  XNOR U1071 ( .A(n1150), .B(n1327), .Z(n1329) );
  XOR U1072 ( .A(n1335), .B(n1336), .Z(n1150) );
  AND U1073 ( .A(n224), .B(n1337), .Z(n1336) );
  XOR U1074 ( .A(n1338), .B(n1335), .Z(n1337) );
  XOR U1075 ( .A(n1339), .B(n1340), .Z(n1327) );
  AND U1076 ( .A(n1341), .B(n1342), .Z(n1340) );
  XOR U1077 ( .A(n1339), .B(n1165), .Z(n1342) );
  XOR U1078 ( .A(n1343), .B(n1344), .Z(n1165) );
  AND U1079 ( .A(n226), .B(n1345), .Z(n1344) );
  XOR U1080 ( .A(n1346), .B(n1343), .Z(n1345) );
  XNOR U1081 ( .A(n1162), .B(n1339), .Z(n1341) );
  XOR U1082 ( .A(n1347), .B(n1348), .Z(n1162) );
  AND U1083 ( .A(n224), .B(n1349), .Z(n1348) );
  XOR U1084 ( .A(n1350), .B(n1347), .Z(n1349) );
  XOR U1085 ( .A(n1351), .B(n1352), .Z(n1339) );
  AND U1086 ( .A(n1353), .B(n1354), .Z(n1352) );
  XOR U1087 ( .A(n1351), .B(n1177), .Z(n1354) );
  XOR U1088 ( .A(n1355), .B(n1356), .Z(n1177) );
  AND U1089 ( .A(n226), .B(n1357), .Z(n1356) );
  XOR U1090 ( .A(n1358), .B(n1355), .Z(n1357) );
  XNOR U1091 ( .A(n1174), .B(n1351), .Z(n1353) );
  XOR U1092 ( .A(n1359), .B(n1360), .Z(n1174) );
  AND U1093 ( .A(n224), .B(n1361), .Z(n1360) );
  XOR U1094 ( .A(n1362), .B(n1359), .Z(n1361) );
  XOR U1095 ( .A(n1363), .B(n1364), .Z(n1351) );
  AND U1096 ( .A(n1365), .B(n1366), .Z(n1364) );
  XOR U1097 ( .A(n1363), .B(n1189), .Z(n1366) );
  XOR U1098 ( .A(n1367), .B(n1368), .Z(n1189) );
  AND U1099 ( .A(n226), .B(n1369), .Z(n1368) );
  XOR U1100 ( .A(n1370), .B(n1367), .Z(n1369) );
  XNOR U1101 ( .A(n1186), .B(n1363), .Z(n1365) );
  XOR U1102 ( .A(n1371), .B(n1372), .Z(n1186) );
  AND U1103 ( .A(n224), .B(n1373), .Z(n1372) );
  XOR U1104 ( .A(n1374), .B(n1371), .Z(n1373) );
  XOR U1105 ( .A(n1375), .B(n1376), .Z(n1363) );
  AND U1106 ( .A(n1377), .B(n1378), .Z(n1376) );
  XOR U1107 ( .A(n1375), .B(n1201), .Z(n1378) );
  XOR U1108 ( .A(n1379), .B(n1380), .Z(n1201) );
  AND U1109 ( .A(n226), .B(n1381), .Z(n1380) );
  XOR U1110 ( .A(n1382), .B(n1379), .Z(n1381) );
  XNOR U1111 ( .A(n1198), .B(n1375), .Z(n1377) );
  XOR U1112 ( .A(n1383), .B(n1384), .Z(n1198) );
  AND U1113 ( .A(n224), .B(n1385), .Z(n1384) );
  XOR U1114 ( .A(n1386), .B(n1383), .Z(n1385) );
  XOR U1115 ( .A(n1387), .B(n1388), .Z(n1375) );
  AND U1116 ( .A(n1389), .B(n1390), .Z(n1388) );
  XOR U1117 ( .A(n1387), .B(n1213), .Z(n1390) );
  XOR U1118 ( .A(n1391), .B(n1392), .Z(n1213) );
  AND U1119 ( .A(n226), .B(n1393), .Z(n1392) );
  XOR U1120 ( .A(n1394), .B(n1391), .Z(n1393) );
  XNOR U1121 ( .A(n1210), .B(n1387), .Z(n1389) );
  XOR U1122 ( .A(n1395), .B(n1396), .Z(n1210) );
  AND U1123 ( .A(n224), .B(n1397), .Z(n1396) );
  XOR U1124 ( .A(n1398), .B(n1395), .Z(n1397) );
  XOR U1125 ( .A(n1399), .B(n1400), .Z(n1387) );
  AND U1126 ( .A(n1401), .B(n1402), .Z(n1400) );
  XOR U1127 ( .A(n1399), .B(n1225), .Z(n1402) );
  XOR U1128 ( .A(n1403), .B(n1404), .Z(n1225) );
  AND U1129 ( .A(n226), .B(n1405), .Z(n1404) );
  XOR U1130 ( .A(n1406), .B(n1403), .Z(n1405) );
  XNOR U1131 ( .A(n1222), .B(n1399), .Z(n1401) );
  XOR U1132 ( .A(n1407), .B(n1408), .Z(n1222) );
  AND U1133 ( .A(n224), .B(n1409), .Z(n1408) );
  XOR U1134 ( .A(n1410), .B(n1407), .Z(n1409) );
  XOR U1135 ( .A(n1411), .B(n1412), .Z(n1399) );
  AND U1136 ( .A(n1413), .B(n1414), .Z(n1412) );
  XOR U1137 ( .A(n1411), .B(n1237), .Z(n1414) );
  XOR U1138 ( .A(n1415), .B(n1416), .Z(n1237) );
  AND U1139 ( .A(n226), .B(n1417), .Z(n1416) );
  XOR U1140 ( .A(n1418), .B(n1415), .Z(n1417) );
  XNOR U1141 ( .A(n1234), .B(n1411), .Z(n1413) );
  XOR U1142 ( .A(n1419), .B(n1420), .Z(n1234) );
  AND U1143 ( .A(n224), .B(n1421), .Z(n1420) );
  XOR U1144 ( .A(n1422), .B(n1419), .Z(n1421) );
  XOR U1145 ( .A(n1423), .B(n1424), .Z(n1411) );
  AND U1146 ( .A(n1425), .B(n1426), .Z(n1424) );
  XOR U1147 ( .A(n1423), .B(n1249), .Z(n1426) );
  XOR U1148 ( .A(n1427), .B(n1428), .Z(n1249) );
  AND U1149 ( .A(n226), .B(n1429), .Z(n1428) );
  XOR U1150 ( .A(n1430), .B(n1427), .Z(n1429) );
  XNOR U1151 ( .A(n1246), .B(n1423), .Z(n1425) );
  XOR U1152 ( .A(n1431), .B(n1432), .Z(n1246) );
  AND U1153 ( .A(n224), .B(n1433), .Z(n1432) );
  XOR U1154 ( .A(n1434), .B(n1431), .Z(n1433) );
  XOR U1155 ( .A(n1435), .B(n1436), .Z(n1423) );
  AND U1156 ( .A(n1437), .B(n1438), .Z(n1436) );
  XOR U1157 ( .A(n1435), .B(n1261), .Z(n1438) );
  XOR U1158 ( .A(n1439), .B(n1440), .Z(n1261) );
  AND U1159 ( .A(n226), .B(n1441), .Z(n1440) );
  XOR U1160 ( .A(n1442), .B(n1439), .Z(n1441) );
  XNOR U1161 ( .A(n1258), .B(n1435), .Z(n1437) );
  XOR U1162 ( .A(n1443), .B(n1444), .Z(n1258) );
  AND U1163 ( .A(n224), .B(n1445), .Z(n1444) );
  XOR U1164 ( .A(n1446), .B(n1443), .Z(n1445) );
  XOR U1165 ( .A(n1447), .B(n1448), .Z(n1435) );
  AND U1166 ( .A(n1449), .B(n1450), .Z(n1448) );
  XOR U1167 ( .A(n1273), .B(n1447), .Z(n1450) );
  XOR U1168 ( .A(n1451), .B(n1452), .Z(n1273) );
  AND U1169 ( .A(n226), .B(n1453), .Z(n1452) );
  XOR U1170 ( .A(n1451), .B(n1454), .Z(n1453) );
  XNOR U1171 ( .A(n1447), .B(n1270), .Z(n1449) );
  XOR U1172 ( .A(n1455), .B(n1456), .Z(n1270) );
  AND U1173 ( .A(n224), .B(n1457), .Z(n1456) );
  XOR U1174 ( .A(n1455), .B(n1458), .Z(n1457) );
  XOR U1175 ( .A(n1459), .B(n1460), .Z(n1447) );
  AND U1176 ( .A(n1461), .B(n1462), .Z(n1460) );
  XNOR U1177 ( .A(n1463), .B(n1286), .Z(n1462) );
  XOR U1178 ( .A(n1464), .B(n1465), .Z(n1286) );
  AND U1179 ( .A(n226), .B(n1466), .Z(n1465) );
  XOR U1180 ( .A(n1467), .B(n1464), .Z(n1466) );
  XNOR U1181 ( .A(n1283), .B(n1459), .Z(n1461) );
  XOR U1182 ( .A(n1468), .B(n1469), .Z(n1283) );
  AND U1183 ( .A(n224), .B(n1470), .Z(n1469) );
  XOR U1184 ( .A(n1471), .B(n1468), .Z(n1470) );
  IV U1185 ( .A(n1463), .Z(n1459) );
  AND U1186 ( .A(n1291), .B(n1294), .Z(n1463) );
  XNOR U1187 ( .A(n1472), .B(n1473), .Z(n1294) );
  AND U1188 ( .A(n226), .B(n1474), .Z(n1473) );
  XNOR U1189 ( .A(n1475), .B(n1472), .Z(n1474) );
  XOR U1190 ( .A(n1476), .B(n1477), .Z(n226) );
  AND U1191 ( .A(n1478), .B(n1479), .Z(n1477) );
  XNOR U1192 ( .A(n1299), .B(n1476), .Z(n1479) );
  AND U1193 ( .A(p_input[2047]), .B(p_input[2031]), .Z(n1299) );
  XOR U1194 ( .A(n1476), .B(n1300), .Z(n1478) );
  AND U1195 ( .A(p_input[2015]), .B(p_input[1999]), .Z(n1300) );
  XOR U1196 ( .A(n1480), .B(n1481), .Z(n1476) );
  AND U1197 ( .A(n1482), .B(n1483), .Z(n1481) );
  XOR U1198 ( .A(n1480), .B(n1310), .Z(n1483) );
  XNOR U1199 ( .A(p_input[2030]), .B(n1484), .Z(n1310) );
  AND U1200 ( .A(n102), .B(n1485), .Z(n1484) );
  XOR U1201 ( .A(p_input[2046]), .B(p_input[2030]), .Z(n1485) );
  XNOR U1202 ( .A(n1307), .B(n1480), .Z(n1482) );
  XOR U1203 ( .A(n1486), .B(n1487), .Z(n1307) );
  AND U1204 ( .A(n100), .B(n1488), .Z(n1487) );
  XOR U1205 ( .A(p_input[2014]), .B(p_input[1998]), .Z(n1488) );
  XOR U1206 ( .A(n1489), .B(n1490), .Z(n1480) );
  AND U1207 ( .A(n1491), .B(n1492), .Z(n1490) );
  XOR U1208 ( .A(n1489), .B(n1322), .Z(n1492) );
  XNOR U1209 ( .A(p_input[2029]), .B(n1493), .Z(n1322) );
  AND U1210 ( .A(n102), .B(n1494), .Z(n1493) );
  XOR U1211 ( .A(p_input[2045]), .B(p_input[2029]), .Z(n1494) );
  XNOR U1212 ( .A(n1319), .B(n1489), .Z(n1491) );
  XOR U1213 ( .A(n1495), .B(n1496), .Z(n1319) );
  AND U1214 ( .A(n100), .B(n1497), .Z(n1496) );
  XOR U1215 ( .A(p_input[2013]), .B(p_input[1997]), .Z(n1497) );
  XOR U1216 ( .A(n1498), .B(n1499), .Z(n1489) );
  AND U1217 ( .A(n1500), .B(n1501), .Z(n1499) );
  XOR U1218 ( .A(n1498), .B(n1334), .Z(n1501) );
  XNOR U1219 ( .A(p_input[2028]), .B(n1502), .Z(n1334) );
  AND U1220 ( .A(n102), .B(n1503), .Z(n1502) );
  XOR U1221 ( .A(p_input[2044]), .B(p_input[2028]), .Z(n1503) );
  XNOR U1222 ( .A(n1331), .B(n1498), .Z(n1500) );
  XOR U1223 ( .A(n1504), .B(n1505), .Z(n1331) );
  AND U1224 ( .A(n100), .B(n1506), .Z(n1505) );
  XOR U1225 ( .A(p_input[2012]), .B(p_input[1996]), .Z(n1506) );
  XOR U1226 ( .A(n1507), .B(n1508), .Z(n1498) );
  AND U1227 ( .A(n1509), .B(n1510), .Z(n1508) );
  XOR U1228 ( .A(n1507), .B(n1346), .Z(n1510) );
  XNOR U1229 ( .A(p_input[2027]), .B(n1511), .Z(n1346) );
  AND U1230 ( .A(n102), .B(n1512), .Z(n1511) );
  XOR U1231 ( .A(p_input[2043]), .B(p_input[2027]), .Z(n1512) );
  XNOR U1232 ( .A(n1343), .B(n1507), .Z(n1509) );
  XOR U1233 ( .A(n1513), .B(n1514), .Z(n1343) );
  AND U1234 ( .A(n100), .B(n1515), .Z(n1514) );
  XOR U1235 ( .A(p_input[2011]), .B(p_input[1995]), .Z(n1515) );
  XOR U1236 ( .A(n1516), .B(n1517), .Z(n1507) );
  AND U1237 ( .A(n1518), .B(n1519), .Z(n1517) );
  XOR U1238 ( .A(n1516), .B(n1358), .Z(n1519) );
  XNOR U1239 ( .A(p_input[2026]), .B(n1520), .Z(n1358) );
  AND U1240 ( .A(n102), .B(n1521), .Z(n1520) );
  XOR U1241 ( .A(p_input[2042]), .B(p_input[2026]), .Z(n1521) );
  XNOR U1242 ( .A(n1355), .B(n1516), .Z(n1518) );
  XOR U1243 ( .A(n1522), .B(n1523), .Z(n1355) );
  AND U1244 ( .A(n100), .B(n1524), .Z(n1523) );
  XOR U1245 ( .A(p_input[2010]), .B(p_input[1994]), .Z(n1524) );
  XOR U1246 ( .A(n1525), .B(n1526), .Z(n1516) );
  AND U1247 ( .A(n1527), .B(n1528), .Z(n1526) );
  XOR U1248 ( .A(n1525), .B(n1370), .Z(n1528) );
  XNOR U1249 ( .A(p_input[2025]), .B(n1529), .Z(n1370) );
  AND U1250 ( .A(n102), .B(n1530), .Z(n1529) );
  XOR U1251 ( .A(p_input[2041]), .B(p_input[2025]), .Z(n1530) );
  XNOR U1252 ( .A(n1367), .B(n1525), .Z(n1527) );
  XOR U1253 ( .A(n1531), .B(n1532), .Z(n1367) );
  AND U1254 ( .A(n100), .B(n1533), .Z(n1532) );
  XOR U1255 ( .A(p_input[2009]), .B(p_input[1993]), .Z(n1533) );
  XOR U1256 ( .A(n1534), .B(n1535), .Z(n1525) );
  AND U1257 ( .A(n1536), .B(n1537), .Z(n1535) );
  XOR U1258 ( .A(n1534), .B(n1382), .Z(n1537) );
  XNOR U1259 ( .A(p_input[2024]), .B(n1538), .Z(n1382) );
  AND U1260 ( .A(n102), .B(n1539), .Z(n1538) );
  XOR U1261 ( .A(p_input[2040]), .B(p_input[2024]), .Z(n1539) );
  XNOR U1262 ( .A(n1379), .B(n1534), .Z(n1536) );
  XOR U1263 ( .A(n1540), .B(n1541), .Z(n1379) );
  AND U1264 ( .A(n100), .B(n1542), .Z(n1541) );
  XOR U1265 ( .A(p_input[2008]), .B(p_input[1992]), .Z(n1542) );
  XOR U1266 ( .A(n1543), .B(n1544), .Z(n1534) );
  AND U1267 ( .A(n1545), .B(n1546), .Z(n1544) );
  XOR U1268 ( .A(n1543), .B(n1394), .Z(n1546) );
  XNOR U1269 ( .A(p_input[2023]), .B(n1547), .Z(n1394) );
  AND U1270 ( .A(n102), .B(n1548), .Z(n1547) );
  XOR U1271 ( .A(p_input[2039]), .B(p_input[2023]), .Z(n1548) );
  XNOR U1272 ( .A(n1391), .B(n1543), .Z(n1545) );
  XOR U1273 ( .A(n1549), .B(n1550), .Z(n1391) );
  AND U1274 ( .A(n100), .B(n1551), .Z(n1550) );
  XOR U1275 ( .A(p_input[2007]), .B(p_input[1991]), .Z(n1551) );
  XOR U1276 ( .A(n1552), .B(n1553), .Z(n1543) );
  AND U1277 ( .A(n1554), .B(n1555), .Z(n1553) );
  XOR U1278 ( .A(n1552), .B(n1406), .Z(n1555) );
  XNOR U1279 ( .A(p_input[2022]), .B(n1556), .Z(n1406) );
  AND U1280 ( .A(n102), .B(n1557), .Z(n1556) );
  XOR U1281 ( .A(p_input[2038]), .B(p_input[2022]), .Z(n1557) );
  XNOR U1282 ( .A(n1403), .B(n1552), .Z(n1554) );
  XOR U1283 ( .A(n1558), .B(n1559), .Z(n1403) );
  AND U1284 ( .A(n100), .B(n1560), .Z(n1559) );
  XOR U1285 ( .A(p_input[2006]), .B(p_input[1990]), .Z(n1560) );
  XOR U1286 ( .A(n1561), .B(n1562), .Z(n1552) );
  AND U1287 ( .A(n1563), .B(n1564), .Z(n1562) );
  XOR U1288 ( .A(n1561), .B(n1418), .Z(n1564) );
  XNOR U1289 ( .A(p_input[2021]), .B(n1565), .Z(n1418) );
  AND U1290 ( .A(n102), .B(n1566), .Z(n1565) );
  XOR U1291 ( .A(p_input[2037]), .B(p_input[2021]), .Z(n1566) );
  XNOR U1292 ( .A(n1415), .B(n1561), .Z(n1563) );
  XOR U1293 ( .A(n1567), .B(n1568), .Z(n1415) );
  AND U1294 ( .A(n100), .B(n1569), .Z(n1568) );
  XOR U1295 ( .A(p_input[2005]), .B(p_input[1989]), .Z(n1569) );
  XOR U1296 ( .A(n1570), .B(n1571), .Z(n1561) );
  AND U1297 ( .A(n1572), .B(n1573), .Z(n1571) );
  XOR U1298 ( .A(n1570), .B(n1430), .Z(n1573) );
  XNOR U1299 ( .A(p_input[2020]), .B(n1574), .Z(n1430) );
  AND U1300 ( .A(n102), .B(n1575), .Z(n1574) );
  XOR U1301 ( .A(p_input[2036]), .B(p_input[2020]), .Z(n1575) );
  XNOR U1302 ( .A(n1427), .B(n1570), .Z(n1572) );
  XOR U1303 ( .A(n1576), .B(n1577), .Z(n1427) );
  AND U1304 ( .A(n100), .B(n1578), .Z(n1577) );
  XOR U1305 ( .A(p_input[2004]), .B(p_input[1988]), .Z(n1578) );
  XOR U1306 ( .A(n1579), .B(n1580), .Z(n1570) );
  AND U1307 ( .A(n1581), .B(n1582), .Z(n1580) );
  XOR U1308 ( .A(n1579), .B(n1442), .Z(n1582) );
  XNOR U1309 ( .A(p_input[2019]), .B(n1583), .Z(n1442) );
  AND U1310 ( .A(n102), .B(n1584), .Z(n1583) );
  XOR U1311 ( .A(p_input[2035]), .B(p_input[2019]), .Z(n1584) );
  XNOR U1312 ( .A(n1439), .B(n1579), .Z(n1581) );
  XOR U1313 ( .A(n1585), .B(n1586), .Z(n1439) );
  AND U1314 ( .A(n100), .B(n1587), .Z(n1586) );
  XOR U1315 ( .A(p_input[2003]), .B(p_input[1987]), .Z(n1587) );
  XOR U1316 ( .A(n1588), .B(n1589), .Z(n1579) );
  AND U1317 ( .A(n1590), .B(n1591), .Z(n1589) );
  XOR U1318 ( .A(n1454), .B(n1588), .Z(n1591) );
  XNOR U1319 ( .A(p_input[2018]), .B(n1592), .Z(n1454) );
  AND U1320 ( .A(n102), .B(n1593), .Z(n1592) );
  XOR U1321 ( .A(p_input[2034]), .B(p_input[2018]), .Z(n1593) );
  XNOR U1322 ( .A(n1588), .B(n1451), .Z(n1590) );
  XOR U1323 ( .A(n1594), .B(n1595), .Z(n1451) );
  AND U1324 ( .A(n100), .B(n1596), .Z(n1595) );
  XOR U1325 ( .A(p_input[2002]), .B(p_input[1986]), .Z(n1596) );
  XOR U1326 ( .A(n1597), .B(n1598), .Z(n1588) );
  AND U1327 ( .A(n1599), .B(n1600), .Z(n1598) );
  XNOR U1328 ( .A(n1601), .B(n1467), .Z(n1600) );
  XNOR U1329 ( .A(p_input[2017]), .B(n1602), .Z(n1467) );
  AND U1330 ( .A(n102), .B(n1603), .Z(n1602) );
  XNOR U1331 ( .A(p_input[2033]), .B(n1604), .Z(n1603) );
  IV U1332 ( .A(p_input[2017]), .Z(n1604) );
  XNOR U1333 ( .A(n1464), .B(n1597), .Z(n1599) );
  XNOR U1334 ( .A(p_input[1985]), .B(n1605), .Z(n1464) );
  AND U1335 ( .A(n100), .B(n1606), .Z(n1605) );
  XOR U1336 ( .A(p_input[2001]), .B(p_input[1985]), .Z(n1606) );
  IV U1337 ( .A(n1601), .Z(n1597) );
  AND U1338 ( .A(n1472), .B(n1475), .Z(n1601) );
  XOR U1339 ( .A(p_input[2016]), .B(n1607), .Z(n1475) );
  AND U1340 ( .A(n102), .B(n1608), .Z(n1607) );
  XOR U1341 ( .A(p_input[2032]), .B(p_input[2016]), .Z(n1608) );
  XOR U1342 ( .A(n1609), .B(n1610), .Z(n102) );
  AND U1343 ( .A(n1611), .B(n1612), .Z(n1610) );
  XNOR U1344 ( .A(p_input[2047]), .B(n1609), .Z(n1612) );
  XOR U1345 ( .A(n1609), .B(p_input[2031]), .Z(n1611) );
  XOR U1346 ( .A(n1613), .B(n1614), .Z(n1609) );
  AND U1347 ( .A(n1615), .B(n1616), .Z(n1614) );
  XNOR U1348 ( .A(p_input[2046]), .B(n1613), .Z(n1616) );
  XOR U1349 ( .A(n1613), .B(p_input[2030]), .Z(n1615) );
  XOR U1350 ( .A(n1617), .B(n1618), .Z(n1613) );
  AND U1351 ( .A(n1619), .B(n1620), .Z(n1618) );
  XNOR U1352 ( .A(p_input[2045]), .B(n1617), .Z(n1620) );
  XOR U1353 ( .A(n1617), .B(p_input[2029]), .Z(n1619) );
  XOR U1354 ( .A(n1621), .B(n1622), .Z(n1617) );
  AND U1355 ( .A(n1623), .B(n1624), .Z(n1622) );
  XNOR U1356 ( .A(p_input[2044]), .B(n1621), .Z(n1624) );
  XOR U1357 ( .A(n1621), .B(p_input[2028]), .Z(n1623) );
  XOR U1358 ( .A(n1625), .B(n1626), .Z(n1621) );
  AND U1359 ( .A(n1627), .B(n1628), .Z(n1626) );
  XNOR U1360 ( .A(p_input[2043]), .B(n1625), .Z(n1628) );
  XOR U1361 ( .A(n1625), .B(p_input[2027]), .Z(n1627) );
  XOR U1362 ( .A(n1629), .B(n1630), .Z(n1625) );
  AND U1363 ( .A(n1631), .B(n1632), .Z(n1630) );
  XNOR U1364 ( .A(p_input[2042]), .B(n1629), .Z(n1632) );
  XOR U1365 ( .A(n1629), .B(p_input[2026]), .Z(n1631) );
  XOR U1366 ( .A(n1633), .B(n1634), .Z(n1629) );
  AND U1367 ( .A(n1635), .B(n1636), .Z(n1634) );
  XNOR U1368 ( .A(p_input[2041]), .B(n1633), .Z(n1636) );
  XOR U1369 ( .A(n1633), .B(p_input[2025]), .Z(n1635) );
  XOR U1370 ( .A(n1637), .B(n1638), .Z(n1633) );
  AND U1371 ( .A(n1639), .B(n1640), .Z(n1638) );
  XNOR U1372 ( .A(p_input[2040]), .B(n1637), .Z(n1640) );
  XOR U1373 ( .A(n1637), .B(p_input[2024]), .Z(n1639) );
  XOR U1374 ( .A(n1641), .B(n1642), .Z(n1637) );
  AND U1375 ( .A(n1643), .B(n1644), .Z(n1642) );
  XNOR U1376 ( .A(p_input[2039]), .B(n1641), .Z(n1644) );
  XOR U1377 ( .A(n1641), .B(p_input[2023]), .Z(n1643) );
  XOR U1378 ( .A(n1645), .B(n1646), .Z(n1641) );
  AND U1379 ( .A(n1647), .B(n1648), .Z(n1646) );
  XNOR U1380 ( .A(p_input[2038]), .B(n1645), .Z(n1648) );
  XOR U1381 ( .A(n1645), .B(p_input[2022]), .Z(n1647) );
  XOR U1382 ( .A(n1649), .B(n1650), .Z(n1645) );
  AND U1383 ( .A(n1651), .B(n1652), .Z(n1650) );
  XNOR U1384 ( .A(p_input[2037]), .B(n1649), .Z(n1652) );
  XOR U1385 ( .A(n1649), .B(p_input[2021]), .Z(n1651) );
  XOR U1386 ( .A(n1653), .B(n1654), .Z(n1649) );
  AND U1387 ( .A(n1655), .B(n1656), .Z(n1654) );
  XNOR U1388 ( .A(p_input[2036]), .B(n1653), .Z(n1656) );
  XOR U1389 ( .A(n1653), .B(p_input[2020]), .Z(n1655) );
  XOR U1390 ( .A(n1657), .B(n1658), .Z(n1653) );
  AND U1391 ( .A(n1659), .B(n1660), .Z(n1658) );
  XNOR U1392 ( .A(p_input[2035]), .B(n1657), .Z(n1660) );
  XOR U1393 ( .A(n1657), .B(p_input[2019]), .Z(n1659) );
  XOR U1394 ( .A(n1661), .B(n1662), .Z(n1657) );
  AND U1395 ( .A(n1663), .B(n1664), .Z(n1662) );
  XNOR U1396 ( .A(p_input[2034]), .B(n1661), .Z(n1664) );
  XOR U1397 ( .A(n1661), .B(p_input[2018]), .Z(n1663) );
  XNOR U1398 ( .A(n1665), .B(n1666), .Z(n1661) );
  AND U1399 ( .A(n1667), .B(n1668), .Z(n1666) );
  XOR U1400 ( .A(p_input[2033]), .B(n1665), .Z(n1668) );
  XNOR U1401 ( .A(p_input[2017]), .B(n1665), .Z(n1667) );
  AND U1402 ( .A(p_input[2032]), .B(n1669), .Z(n1665) );
  IV U1403 ( .A(p_input[2016]), .Z(n1669) );
  XNOR U1404 ( .A(p_input[1984]), .B(n1670), .Z(n1472) );
  AND U1405 ( .A(n100), .B(n1671), .Z(n1670) );
  XOR U1406 ( .A(p_input[2000]), .B(p_input[1984]), .Z(n1671) );
  XOR U1407 ( .A(n1672), .B(n1673), .Z(n100) );
  AND U1408 ( .A(n1674), .B(n1675), .Z(n1673) );
  XNOR U1409 ( .A(p_input[2015]), .B(n1672), .Z(n1675) );
  XOR U1410 ( .A(n1672), .B(p_input[1999]), .Z(n1674) );
  XOR U1411 ( .A(n1676), .B(n1677), .Z(n1672) );
  AND U1412 ( .A(n1678), .B(n1679), .Z(n1677) );
  XNOR U1413 ( .A(p_input[2014]), .B(n1676), .Z(n1679) );
  XNOR U1414 ( .A(n1676), .B(n1486), .Z(n1678) );
  IV U1415 ( .A(p_input[1998]), .Z(n1486) );
  XOR U1416 ( .A(n1680), .B(n1681), .Z(n1676) );
  AND U1417 ( .A(n1682), .B(n1683), .Z(n1681) );
  XNOR U1418 ( .A(p_input[2013]), .B(n1680), .Z(n1683) );
  XNOR U1419 ( .A(n1680), .B(n1495), .Z(n1682) );
  IV U1420 ( .A(p_input[1997]), .Z(n1495) );
  XOR U1421 ( .A(n1684), .B(n1685), .Z(n1680) );
  AND U1422 ( .A(n1686), .B(n1687), .Z(n1685) );
  XNOR U1423 ( .A(p_input[2012]), .B(n1684), .Z(n1687) );
  XNOR U1424 ( .A(n1684), .B(n1504), .Z(n1686) );
  IV U1425 ( .A(p_input[1996]), .Z(n1504) );
  XOR U1426 ( .A(n1688), .B(n1689), .Z(n1684) );
  AND U1427 ( .A(n1690), .B(n1691), .Z(n1689) );
  XNOR U1428 ( .A(p_input[2011]), .B(n1688), .Z(n1691) );
  XNOR U1429 ( .A(n1688), .B(n1513), .Z(n1690) );
  IV U1430 ( .A(p_input[1995]), .Z(n1513) );
  XOR U1431 ( .A(n1692), .B(n1693), .Z(n1688) );
  AND U1432 ( .A(n1694), .B(n1695), .Z(n1693) );
  XNOR U1433 ( .A(p_input[2010]), .B(n1692), .Z(n1695) );
  XNOR U1434 ( .A(n1692), .B(n1522), .Z(n1694) );
  IV U1435 ( .A(p_input[1994]), .Z(n1522) );
  XOR U1436 ( .A(n1696), .B(n1697), .Z(n1692) );
  AND U1437 ( .A(n1698), .B(n1699), .Z(n1697) );
  XNOR U1438 ( .A(p_input[2009]), .B(n1696), .Z(n1699) );
  XNOR U1439 ( .A(n1696), .B(n1531), .Z(n1698) );
  IV U1440 ( .A(p_input[1993]), .Z(n1531) );
  XOR U1441 ( .A(n1700), .B(n1701), .Z(n1696) );
  AND U1442 ( .A(n1702), .B(n1703), .Z(n1701) );
  XNOR U1443 ( .A(p_input[2008]), .B(n1700), .Z(n1703) );
  XNOR U1444 ( .A(n1700), .B(n1540), .Z(n1702) );
  IV U1445 ( .A(p_input[1992]), .Z(n1540) );
  XOR U1446 ( .A(n1704), .B(n1705), .Z(n1700) );
  AND U1447 ( .A(n1706), .B(n1707), .Z(n1705) );
  XNOR U1448 ( .A(p_input[2007]), .B(n1704), .Z(n1707) );
  XNOR U1449 ( .A(n1704), .B(n1549), .Z(n1706) );
  IV U1450 ( .A(p_input[1991]), .Z(n1549) );
  XOR U1451 ( .A(n1708), .B(n1709), .Z(n1704) );
  AND U1452 ( .A(n1710), .B(n1711), .Z(n1709) );
  XNOR U1453 ( .A(p_input[2006]), .B(n1708), .Z(n1711) );
  XNOR U1454 ( .A(n1708), .B(n1558), .Z(n1710) );
  IV U1455 ( .A(p_input[1990]), .Z(n1558) );
  XOR U1456 ( .A(n1712), .B(n1713), .Z(n1708) );
  AND U1457 ( .A(n1714), .B(n1715), .Z(n1713) );
  XNOR U1458 ( .A(p_input[2005]), .B(n1712), .Z(n1715) );
  XNOR U1459 ( .A(n1712), .B(n1567), .Z(n1714) );
  IV U1460 ( .A(p_input[1989]), .Z(n1567) );
  XOR U1461 ( .A(n1716), .B(n1717), .Z(n1712) );
  AND U1462 ( .A(n1718), .B(n1719), .Z(n1717) );
  XNOR U1463 ( .A(p_input[2004]), .B(n1716), .Z(n1719) );
  XNOR U1464 ( .A(n1716), .B(n1576), .Z(n1718) );
  IV U1465 ( .A(p_input[1988]), .Z(n1576) );
  XOR U1466 ( .A(n1720), .B(n1721), .Z(n1716) );
  AND U1467 ( .A(n1722), .B(n1723), .Z(n1721) );
  XNOR U1468 ( .A(p_input[2003]), .B(n1720), .Z(n1723) );
  XNOR U1469 ( .A(n1720), .B(n1585), .Z(n1722) );
  IV U1470 ( .A(p_input[1987]), .Z(n1585) );
  XOR U1471 ( .A(n1724), .B(n1725), .Z(n1720) );
  AND U1472 ( .A(n1726), .B(n1727), .Z(n1725) );
  XNOR U1473 ( .A(p_input[2002]), .B(n1724), .Z(n1727) );
  XNOR U1474 ( .A(n1724), .B(n1594), .Z(n1726) );
  IV U1475 ( .A(p_input[1986]), .Z(n1594) );
  XNOR U1476 ( .A(n1728), .B(n1729), .Z(n1724) );
  AND U1477 ( .A(n1730), .B(n1731), .Z(n1729) );
  XOR U1478 ( .A(p_input[2001]), .B(n1728), .Z(n1731) );
  XNOR U1479 ( .A(p_input[1985]), .B(n1728), .Z(n1730) );
  AND U1480 ( .A(p_input[2000]), .B(n1732), .Z(n1728) );
  IV U1481 ( .A(p_input[1984]), .Z(n1732) );
  XOR U1482 ( .A(n1733), .B(n1734), .Z(n1291) );
  AND U1483 ( .A(n224), .B(n1735), .Z(n1734) );
  XNOR U1484 ( .A(n1736), .B(n1733), .Z(n1735) );
  XOR U1485 ( .A(n1737), .B(n1738), .Z(n224) );
  AND U1486 ( .A(n1739), .B(n1740), .Z(n1738) );
  XNOR U1487 ( .A(n1301), .B(n1737), .Z(n1740) );
  AND U1488 ( .A(p_input[1983]), .B(p_input[1967]), .Z(n1301) );
  XOR U1489 ( .A(n1737), .B(n1302), .Z(n1739) );
  AND U1490 ( .A(p_input[1951]), .B(p_input[1935]), .Z(n1302) );
  XOR U1491 ( .A(n1741), .B(n1742), .Z(n1737) );
  AND U1492 ( .A(n1743), .B(n1744), .Z(n1742) );
  XOR U1493 ( .A(n1741), .B(n1314), .Z(n1744) );
  XNOR U1494 ( .A(p_input[1966]), .B(n1745), .Z(n1314) );
  AND U1495 ( .A(n106), .B(n1746), .Z(n1745) );
  XOR U1496 ( .A(p_input[1982]), .B(p_input[1966]), .Z(n1746) );
  XNOR U1497 ( .A(n1311), .B(n1741), .Z(n1743) );
  XOR U1498 ( .A(n1747), .B(n1748), .Z(n1311) );
  AND U1499 ( .A(n103), .B(n1749), .Z(n1748) );
  XOR U1500 ( .A(p_input[1950]), .B(p_input[1934]), .Z(n1749) );
  XOR U1501 ( .A(n1750), .B(n1751), .Z(n1741) );
  AND U1502 ( .A(n1752), .B(n1753), .Z(n1751) );
  XOR U1503 ( .A(n1750), .B(n1326), .Z(n1753) );
  XNOR U1504 ( .A(p_input[1965]), .B(n1754), .Z(n1326) );
  AND U1505 ( .A(n106), .B(n1755), .Z(n1754) );
  XOR U1506 ( .A(p_input[1981]), .B(p_input[1965]), .Z(n1755) );
  XNOR U1507 ( .A(n1323), .B(n1750), .Z(n1752) );
  XOR U1508 ( .A(n1756), .B(n1757), .Z(n1323) );
  AND U1509 ( .A(n103), .B(n1758), .Z(n1757) );
  XOR U1510 ( .A(p_input[1949]), .B(p_input[1933]), .Z(n1758) );
  XOR U1511 ( .A(n1759), .B(n1760), .Z(n1750) );
  AND U1512 ( .A(n1761), .B(n1762), .Z(n1760) );
  XOR U1513 ( .A(n1759), .B(n1338), .Z(n1762) );
  XNOR U1514 ( .A(p_input[1964]), .B(n1763), .Z(n1338) );
  AND U1515 ( .A(n106), .B(n1764), .Z(n1763) );
  XOR U1516 ( .A(p_input[1980]), .B(p_input[1964]), .Z(n1764) );
  XNOR U1517 ( .A(n1335), .B(n1759), .Z(n1761) );
  XOR U1518 ( .A(n1765), .B(n1766), .Z(n1335) );
  AND U1519 ( .A(n103), .B(n1767), .Z(n1766) );
  XOR U1520 ( .A(p_input[1948]), .B(p_input[1932]), .Z(n1767) );
  XOR U1521 ( .A(n1768), .B(n1769), .Z(n1759) );
  AND U1522 ( .A(n1770), .B(n1771), .Z(n1769) );
  XOR U1523 ( .A(n1768), .B(n1350), .Z(n1771) );
  XNOR U1524 ( .A(p_input[1963]), .B(n1772), .Z(n1350) );
  AND U1525 ( .A(n106), .B(n1773), .Z(n1772) );
  XOR U1526 ( .A(p_input[1979]), .B(p_input[1963]), .Z(n1773) );
  XNOR U1527 ( .A(n1347), .B(n1768), .Z(n1770) );
  XOR U1528 ( .A(n1774), .B(n1775), .Z(n1347) );
  AND U1529 ( .A(n103), .B(n1776), .Z(n1775) );
  XOR U1530 ( .A(p_input[1947]), .B(p_input[1931]), .Z(n1776) );
  XOR U1531 ( .A(n1777), .B(n1778), .Z(n1768) );
  AND U1532 ( .A(n1779), .B(n1780), .Z(n1778) );
  XOR U1533 ( .A(n1777), .B(n1362), .Z(n1780) );
  XNOR U1534 ( .A(p_input[1962]), .B(n1781), .Z(n1362) );
  AND U1535 ( .A(n106), .B(n1782), .Z(n1781) );
  XOR U1536 ( .A(p_input[1978]), .B(p_input[1962]), .Z(n1782) );
  XNOR U1537 ( .A(n1359), .B(n1777), .Z(n1779) );
  XOR U1538 ( .A(n1783), .B(n1784), .Z(n1359) );
  AND U1539 ( .A(n103), .B(n1785), .Z(n1784) );
  XOR U1540 ( .A(p_input[1946]), .B(p_input[1930]), .Z(n1785) );
  XOR U1541 ( .A(n1786), .B(n1787), .Z(n1777) );
  AND U1542 ( .A(n1788), .B(n1789), .Z(n1787) );
  XOR U1543 ( .A(n1786), .B(n1374), .Z(n1789) );
  XNOR U1544 ( .A(p_input[1961]), .B(n1790), .Z(n1374) );
  AND U1545 ( .A(n106), .B(n1791), .Z(n1790) );
  XOR U1546 ( .A(p_input[1977]), .B(p_input[1961]), .Z(n1791) );
  XNOR U1547 ( .A(n1371), .B(n1786), .Z(n1788) );
  XOR U1548 ( .A(n1792), .B(n1793), .Z(n1371) );
  AND U1549 ( .A(n103), .B(n1794), .Z(n1793) );
  XOR U1550 ( .A(p_input[1945]), .B(p_input[1929]), .Z(n1794) );
  XOR U1551 ( .A(n1795), .B(n1796), .Z(n1786) );
  AND U1552 ( .A(n1797), .B(n1798), .Z(n1796) );
  XOR U1553 ( .A(n1795), .B(n1386), .Z(n1798) );
  XNOR U1554 ( .A(p_input[1960]), .B(n1799), .Z(n1386) );
  AND U1555 ( .A(n106), .B(n1800), .Z(n1799) );
  XOR U1556 ( .A(p_input[1976]), .B(p_input[1960]), .Z(n1800) );
  XNOR U1557 ( .A(n1383), .B(n1795), .Z(n1797) );
  XOR U1558 ( .A(n1801), .B(n1802), .Z(n1383) );
  AND U1559 ( .A(n103), .B(n1803), .Z(n1802) );
  XOR U1560 ( .A(p_input[1944]), .B(p_input[1928]), .Z(n1803) );
  XOR U1561 ( .A(n1804), .B(n1805), .Z(n1795) );
  AND U1562 ( .A(n1806), .B(n1807), .Z(n1805) );
  XOR U1563 ( .A(n1804), .B(n1398), .Z(n1807) );
  XNOR U1564 ( .A(p_input[1959]), .B(n1808), .Z(n1398) );
  AND U1565 ( .A(n106), .B(n1809), .Z(n1808) );
  XOR U1566 ( .A(p_input[1975]), .B(p_input[1959]), .Z(n1809) );
  XNOR U1567 ( .A(n1395), .B(n1804), .Z(n1806) );
  XOR U1568 ( .A(n1810), .B(n1811), .Z(n1395) );
  AND U1569 ( .A(n103), .B(n1812), .Z(n1811) );
  XOR U1570 ( .A(p_input[1943]), .B(p_input[1927]), .Z(n1812) );
  XOR U1571 ( .A(n1813), .B(n1814), .Z(n1804) );
  AND U1572 ( .A(n1815), .B(n1816), .Z(n1814) );
  XOR U1573 ( .A(n1813), .B(n1410), .Z(n1816) );
  XNOR U1574 ( .A(p_input[1958]), .B(n1817), .Z(n1410) );
  AND U1575 ( .A(n106), .B(n1818), .Z(n1817) );
  XOR U1576 ( .A(p_input[1974]), .B(p_input[1958]), .Z(n1818) );
  XNOR U1577 ( .A(n1407), .B(n1813), .Z(n1815) );
  XOR U1578 ( .A(n1819), .B(n1820), .Z(n1407) );
  AND U1579 ( .A(n103), .B(n1821), .Z(n1820) );
  XOR U1580 ( .A(p_input[1942]), .B(p_input[1926]), .Z(n1821) );
  XOR U1581 ( .A(n1822), .B(n1823), .Z(n1813) );
  AND U1582 ( .A(n1824), .B(n1825), .Z(n1823) );
  XOR U1583 ( .A(n1822), .B(n1422), .Z(n1825) );
  XNOR U1584 ( .A(p_input[1957]), .B(n1826), .Z(n1422) );
  AND U1585 ( .A(n106), .B(n1827), .Z(n1826) );
  XOR U1586 ( .A(p_input[1973]), .B(p_input[1957]), .Z(n1827) );
  XNOR U1587 ( .A(n1419), .B(n1822), .Z(n1824) );
  XOR U1588 ( .A(n1828), .B(n1829), .Z(n1419) );
  AND U1589 ( .A(n103), .B(n1830), .Z(n1829) );
  XOR U1590 ( .A(p_input[1941]), .B(p_input[1925]), .Z(n1830) );
  XOR U1591 ( .A(n1831), .B(n1832), .Z(n1822) );
  AND U1592 ( .A(n1833), .B(n1834), .Z(n1832) );
  XOR U1593 ( .A(n1831), .B(n1434), .Z(n1834) );
  XNOR U1594 ( .A(p_input[1956]), .B(n1835), .Z(n1434) );
  AND U1595 ( .A(n106), .B(n1836), .Z(n1835) );
  XOR U1596 ( .A(p_input[1972]), .B(p_input[1956]), .Z(n1836) );
  XNOR U1597 ( .A(n1431), .B(n1831), .Z(n1833) );
  XOR U1598 ( .A(n1837), .B(n1838), .Z(n1431) );
  AND U1599 ( .A(n103), .B(n1839), .Z(n1838) );
  XOR U1600 ( .A(p_input[1940]), .B(p_input[1924]), .Z(n1839) );
  XOR U1601 ( .A(n1840), .B(n1841), .Z(n1831) );
  AND U1602 ( .A(n1842), .B(n1843), .Z(n1841) );
  XOR U1603 ( .A(n1840), .B(n1446), .Z(n1843) );
  XNOR U1604 ( .A(p_input[1955]), .B(n1844), .Z(n1446) );
  AND U1605 ( .A(n106), .B(n1845), .Z(n1844) );
  XOR U1606 ( .A(p_input[1971]), .B(p_input[1955]), .Z(n1845) );
  XNOR U1607 ( .A(n1443), .B(n1840), .Z(n1842) );
  XOR U1608 ( .A(n1846), .B(n1847), .Z(n1443) );
  AND U1609 ( .A(n103), .B(n1848), .Z(n1847) );
  XOR U1610 ( .A(p_input[1939]), .B(p_input[1923]), .Z(n1848) );
  XOR U1611 ( .A(n1849), .B(n1850), .Z(n1840) );
  AND U1612 ( .A(n1851), .B(n1852), .Z(n1850) );
  XOR U1613 ( .A(n1458), .B(n1849), .Z(n1852) );
  XNOR U1614 ( .A(p_input[1954]), .B(n1853), .Z(n1458) );
  AND U1615 ( .A(n106), .B(n1854), .Z(n1853) );
  XOR U1616 ( .A(p_input[1970]), .B(p_input[1954]), .Z(n1854) );
  XNOR U1617 ( .A(n1849), .B(n1455), .Z(n1851) );
  XOR U1618 ( .A(n1855), .B(n1856), .Z(n1455) );
  AND U1619 ( .A(n103), .B(n1857), .Z(n1856) );
  XOR U1620 ( .A(p_input[1938]), .B(p_input[1922]), .Z(n1857) );
  XOR U1621 ( .A(n1858), .B(n1859), .Z(n1849) );
  AND U1622 ( .A(n1860), .B(n1861), .Z(n1859) );
  XNOR U1623 ( .A(n1862), .B(n1471), .Z(n1861) );
  XNOR U1624 ( .A(p_input[1953]), .B(n1863), .Z(n1471) );
  AND U1625 ( .A(n106), .B(n1864), .Z(n1863) );
  XNOR U1626 ( .A(p_input[1969]), .B(n1865), .Z(n1864) );
  IV U1627 ( .A(p_input[1953]), .Z(n1865) );
  XNOR U1628 ( .A(n1468), .B(n1858), .Z(n1860) );
  XNOR U1629 ( .A(p_input[1921]), .B(n1866), .Z(n1468) );
  AND U1630 ( .A(n103), .B(n1867), .Z(n1866) );
  XOR U1631 ( .A(p_input[1937]), .B(p_input[1921]), .Z(n1867) );
  IV U1632 ( .A(n1862), .Z(n1858) );
  AND U1633 ( .A(n1733), .B(n1736), .Z(n1862) );
  XOR U1634 ( .A(p_input[1952]), .B(n1868), .Z(n1736) );
  AND U1635 ( .A(n106), .B(n1869), .Z(n1868) );
  XOR U1636 ( .A(p_input[1968]), .B(p_input[1952]), .Z(n1869) );
  XOR U1637 ( .A(n1870), .B(n1871), .Z(n106) );
  AND U1638 ( .A(n1872), .B(n1873), .Z(n1871) );
  XNOR U1639 ( .A(p_input[1983]), .B(n1870), .Z(n1873) );
  XOR U1640 ( .A(n1870), .B(p_input[1967]), .Z(n1872) );
  XOR U1641 ( .A(n1874), .B(n1875), .Z(n1870) );
  AND U1642 ( .A(n1876), .B(n1877), .Z(n1875) );
  XNOR U1643 ( .A(p_input[1982]), .B(n1874), .Z(n1877) );
  XOR U1644 ( .A(n1874), .B(p_input[1966]), .Z(n1876) );
  XOR U1645 ( .A(n1878), .B(n1879), .Z(n1874) );
  AND U1646 ( .A(n1880), .B(n1881), .Z(n1879) );
  XNOR U1647 ( .A(p_input[1981]), .B(n1878), .Z(n1881) );
  XOR U1648 ( .A(n1878), .B(p_input[1965]), .Z(n1880) );
  XOR U1649 ( .A(n1882), .B(n1883), .Z(n1878) );
  AND U1650 ( .A(n1884), .B(n1885), .Z(n1883) );
  XNOR U1651 ( .A(p_input[1980]), .B(n1882), .Z(n1885) );
  XOR U1652 ( .A(n1882), .B(p_input[1964]), .Z(n1884) );
  XOR U1653 ( .A(n1886), .B(n1887), .Z(n1882) );
  AND U1654 ( .A(n1888), .B(n1889), .Z(n1887) );
  XNOR U1655 ( .A(p_input[1979]), .B(n1886), .Z(n1889) );
  XOR U1656 ( .A(n1886), .B(p_input[1963]), .Z(n1888) );
  XOR U1657 ( .A(n1890), .B(n1891), .Z(n1886) );
  AND U1658 ( .A(n1892), .B(n1893), .Z(n1891) );
  XNOR U1659 ( .A(p_input[1978]), .B(n1890), .Z(n1893) );
  XOR U1660 ( .A(n1890), .B(p_input[1962]), .Z(n1892) );
  XOR U1661 ( .A(n1894), .B(n1895), .Z(n1890) );
  AND U1662 ( .A(n1896), .B(n1897), .Z(n1895) );
  XNOR U1663 ( .A(p_input[1977]), .B(n1894), .Z(n1897) );
  XOR U1664 ( .A(n1894), .B(p_input[1961]), .Z(n1896) );
  XOR U1665 ( .A(n1898), .B(n1899), .Z(n1894) );
  AND U1666 ( .A(n1900), .B(n1901), .Z(n1899) );
  XNOR U1667 ( .A(p_input[1976]), .B(n1898), .Z(n1901) );
  XOR U1668 ( .A(n1898), .B(p_input[1960]), .Z(n1900) );
  XOR U1669 ( .A(n1902), .B(n1903), .Z(n1898) );
  AND U1670 ( .A(n1904), .B(n1905), .Z(n1903) );
  XNOR U1671 ( .A(p_input[1975]), .B(n1902), .Z(n1905) );
  XOR U1672 ( .A(n1902), .B(p_input[1959]), .Z(n1904) );
  XOR U1673 ( .A(n1906), .B(n1907), .Z(n1902) );
  AND U1674 ( .A(n1908), .B(n1909), .Z(n1907) );
  XNOR U1675 ( .A(p_input[1974]), .B(n1906), .Z(n1909) );
  XOR U1676 ( .A(n1906), .B(p_input[1958]), .Z(n1908) );
  XOR U1677 ( .A(n1910), .B(n1911), .Z(n1906) );
  AND U1678 ( .A(n1912), .B(n1913), .Z(n1911) );
  XNOR U1679 ( .A(p_input[1973]), .B(n1910), .Z(n1913) );
  XOR U1680 ( .A(n1910), .B(p_input[1957]), .Z(n1912) );
  XOR U1681 ( .A(n1914), .B(n1915), .Z(n1910) );
  AND U1682 ( .A(n1916), .B(n1917), .Z(n1915) );
  XNOR U1683 ( .A(p_input[1972]), .B(n1914), .Z(n1917) );
  XOR U1684 ( .A(n1914), .B(p_input[1956]), .Z(n1916) );
  XOR U1685 ( .A(n1918), .B(n1919), .Z(n1914) );
  AND U1686 ( .A(n1920), .B(n1921), .Z(n1919) );
  XNOR U1687 ( .A(p_input[1971]), .B(n1918), .Z(n1921) );
  XOR U1688 ( .A(n1918), .B(p_input[1955]), .Z(n1920) );
  XOR U1689 ( .A(n1922), .B(n1923), .Z(n1918) );
  AND U1690 ( .A(n1924), .B(n1925), .Z(n1923) );
  XNOR U1691 ( .A(p_input[1970]), .B(n1922), .Z(n1925) );
  XOR U1692 ( .A(n1922), .B(p_input[1954]), .Z(n1924) );
  XNOR U1693 ( .A(n1926), .B(n1927), .Z(n1922) );
  AND U1694 ( .A(n1928), .B(n1929), .Z(n1927) );
  XOR U1695 ( .A(p_input[1969]), .B(n1926), .Z(n1929) );
  XNOR U1696 ( .A(p_input[1953]), .B(n1926), .Z(n1928) );
  AND U1697 ( .A(p_input[1968]), .B(n1930), .Z(n1926) );
  IV U1698 ( .A(p_input[1952]), .Z(n1930) );
  XNOR U1699 ( .A(p_input[1920]), .B(n1931), .Z(n1733) );
  AND U1700 ( .A(n103), .B(n1932), .Z(n1931) );
  XOR U1701 ( .A(p_input[1936]), .B(p_input[1920]), .Z(n1932) );
  XOR U1702 ( .A(n1933), .B(n1934), .Z(n103) );
  AND U1703 ( .A(n1935), .B(n1936), .Z(n1934) );
  XNOR U1704 ( .A(p_input[1951]), .B(n1933), .Z(n1936) );
  XOR U1705 ( .A(n1933), .B(p_input[1935]), .Z(n1935) );
  XOR U1706 ( .A(n1937), .B(n1938), .Z(n1933) );
  AND U1707 ( .A(n1939), .B(n1940), .Z(n1938) );
  XNOR U1708 ( .A(p_input[1950]), .B(n1937), .Z(n1940) );
  XNOR U1709 ( .A(n1937), .B(n1747), .Z(n1939) );
  IV U1710 ( .A(p_input[1934]), .Z(n1747) );
  XOR U1711 ( .A(n1941), .B(n1942), .Z(n1937) );
  AND U1712 ( .A(n1943), .B(n1944), .Z(n1942) );
  XNOR U1713 ( .A(p_input[1949]), .B(n1941), .Z(n1944) );
  XNOR U1714 ( .A(n1941), .B(n1756), .Z(n1943) );
  IV U1715 ( .A(p_input[1933]), .Z(n1756) );
  XOR U1716 ( .A(n1945), .B(n1946), .Z(n1941) );
  AND U1717 ( .A(n1947), .B(n1948), .Z(n1946) );
  XNOR U1718 ( .A(p_input[1948]), .B(n1945), .Z(n1948) );
  XNOR U1719 ( .A(n1945), .B(n1765), .Z(n1947) );
  IV U1720 ( .A(p_input[1932]), .Z(n1765) );
  XOR U1721 ( .A(n1949), .B(n1950), .Z(n1945) );
  AND U1722 ( .A(n1951), .B(n1952), .Z(n1950) );
  XNOR U1723 ( .A(p_input[1947]), .B(n1949), .Z(n1952) );
  XNOR U1724 ( .A(n1949), .B(n1774), .Z(n1951) );
  IV U1725 ( .A(p_input[1931]), .Z(n1774) );
  XOR U1726 ( .A(n1953), .B(n1954), .Z(n1949) );
  AND U1727 ( .A(n1955), .B(n1956), .Z(n1954) );
  XNOR U1728 ( .A(p_input[1946]), .B(n1953), .Z(n1956) );
  XNOR U1729 ( .A(n1953), .B(n1783), .Z(n1955) );
  IV U1730 ( .A(p_input[1930]), .Z(n1783) );
  XOR U1731 ( .A(n1957), .B(n1958), .Z(n1953) );
  AND U1732 ( .A(n1959), .B(n1960), .Z(n1958) );
  XNOR U1733 ( .A(p_input[1945]), .B(n1957), .Z(n1960) );
  XNOR U1734 ( .A(n1957), .B(n1792), .Z(n1959) );
  IV U1735 ( .A(p_input[1929]), .Z(n1792) );
  XOR U1736 ( .A(n1961), .B(n1962), .Z(n1957) );
  AND U1737 ( .A(n1963), .B(n1964), .Z(n1962) );
  XNOR U1738 ( .A(p_input[1944]), .B(n1961), .Z(n1964) );
  XNOR U1739 ( .A(n1961), .B(n1801), .Z(n1963) );
  IV U1740 ( .A(p_input[1928]), .Z(n1801) );
  XOR U1741 ( .A(n1965), .B(n1966), .Z(n1961) );
  AND U1742 ( .A(n1967), .B(n1968), .Z(n1966) );
  XNOR U1743 ( .A(p_input[1943]), .B(n1965), .Z(n1968) );
  XNOR U1744 ( .A(n1965), .B(n1810), .Z(n1967) );
  IV U1745 ( .A(p_input[1927]), .Z(n1810) );
  XOR U1746 ( .A(n1969), .B(n1970), .Z(n1965) );
  AND U1747 ( .A(n1971), .B(n1972), .Z(n1970) );
  XNOR U1748 ( .A(p_input[1942]), .B(n1969), .Z(n1972) );
  XNOR U1749 ( .A(n1969), .B(n1819), .Z(n1971) );
  IV U1750 ( .A(p_input[1926]), .Z(n1819) );
  XOR U1751 ( .A(n1973), .B(n1974), .Z(n1969) );
  AND U1752 ( .A(n1975), .B(n1976), .Z(n1974) );
  XNOR U1753 ( .A(p_input[1941]), .B(n1973), .Z(n1976) );
  XNOR U1754 ( .A(n1973), .B(n1828), .Z(n1975) );
  IV U1755 ( .A(p_input[1925]), .Z(n1828) );
  XOR U1756 ( .A(n1977), .B(n1978), .Z(n1973) );
  AND U1757 ( .A(n1979), .B(n1980), .Z(n1978) );
  XNOR U1758 ( .A(p_input[1940]), .B(n1977), .Z(n1980) );
  XNOR U1759 ( .A(n1977), .B(n1837), .Z(n1979) );
  IV U1760 ( .A(p_input[1924]), .Z(n1837) );
  XOR U1761 ( .A(n1981), .B(n1982), .Z(n1977) );
  AND U1762 ( .A(n1983), .B(n1984), .Z(n1982) );
  XNOR U1763 ( .A(p_input[1939]), .B(n1981), .Z(n1984) );
  XNOR U1764 ( .A(n1981), .B(n1846), .Z(n1983) );
  IV U1765 ( .A(p_input[1923]), .Z(n1846) );
  XOR U1766 ( .A(n1985), .B(n1986), .Z(n1981) );
  AND U1767 ( .A(n1987), .B(n1988), .Z(n1986) );
  XNOR U1768 ( .A(p_input[1938]), .B(n1985), .Z(n1988) );
  XNOR U1769 ( .A(n1985), .B(n1855), .Z(n1987) );
  IV U1770 ( .A(p_input[1922]), .Z(n1855) );
  XNOR U1771 ( .A(n1989), .B(n1990), .Z(n1985) );
  AND U1772 ( .A(n1991), .B(n1992), .Z(n1990) );
  XOR U1773 ( .A(p_input[1937]), .B(n1989), .Z(n1992) );
  XNOR U1774 ( .A(p_input[1921]), .B(n1989), .Z(n1991) );
  AND U1775 ( .A(p_input[1936]), .B(n1993), .Z(n1989) );
  IV U1776 ( .A(p_input[1920]), .Z(n1993) );
  XOR U1777 ( .A(n1994), .B(n1995), .Z(n1109) );
  AND U1778 ( .A(n408), .B(n1996), .Z(n1995) );
  XNOR U1779 ( .A(n1997), .B(n1994), .Z(n1996) );
  XOR U1780 ( .A(n1998), .B(n1999), .Z(n408) );
  AND U1781 ( .A(n2000), .B(n2001), .Z(n1999) );
  XNOR U1782 ( .A(n1121), .B(n1998), .Z(n2001) );
  AND U1783 ( .A(n2002), .B(n2003), .Z(n1121) );
  XOR U1784 ( .A(n1998), .B(n1120), .Z(n2000) );
  AND U1785 ( .A(n2004), .B(n2005), .Z(n1120) );
  XOR U1786 ( .A(n2006), .B(n2007), .Z(n1998) );
  AND U1787 ( .A(n2008), .B(n2009), .Z(n2007) );
  XOR U1788 ( .A(n2006), .B(n1133), .Z(n2009) );
  XOR U1789 ( .A(n2010), .B(n2011), .Z(n1133) );
  AND U1790 ( .A(n230), .B(n2012), .Z(n2011) );
  XOR U1791 ( .A(n2013), .B(n2010), .Z(n2012) );
  XNOR U1792 ( .A(n1130), .B(n2006), .Z(n2008) );
  XOR U1793 ( .A(n2014), .B(n2015), .Z(n1130) );
  AND U1794 ( .A(n227), .B(n2016), .Z(n2015) );
  XOR U1795 ( .A(n2017), .B(n2014), .Z(n2016) );
  XOR U1796 ( .A(n2018), .B(n2019), .Z(n2006) );
  AND U1797 ( .A(n2020), .B(n2021), .Z(n2019) );
  XOR U1798 ( .A(n2018), .B(n1145), .Z(n2021) );
  XOR U1799 ( .A(n2022), .B(n2023), .Z(n1145) );
  AND U1800 ( .A(n230), .B(n2024), .Z(n2023) );
  XOR U1801 ( .A(n2025), .B(n2022), .Z(n2024) );
  XNOR U1802 ( .A(n1142), .B(n2018), .Z(n2020) );
  XOR U1803 ( .A(n2026), .B(n2027), .Z(n1142) );
  AND U1804 ( .A(n227), .B(n2028), .Z(n2027) );
  XOR U1805 ( .A(n2029), .B(n2026), .Z(n2028) );
  XOR U1806 ( .A(n2030), .B(n2031), .Z(n2018) );
  AND U1807 ( .A(n2032), .B(n2033), .Z(n2031) );
  XOR U1808 ( .A(n2030), .B(n1157), .Z(n2033) );
  XOR U1809 ( .A(n2034), .B(n2035), .Z(n1157) );
  AND U1810 ( .A(n230), .B(n2036), .Z(n2035) );
  XOR U1811 ( .A(n2037), .B(n2034), .Z(n2036) );
  XNOR U1812 ( .A(n1154), .B(n2030), .Z(n2032) );
  XOR U1813 ( .A(n2038), .B(n2039), .Z(n1154) );
  AND U1814 ( .A(n227), .B(n2040), .Z(n2039) );
  XOR U1815 ( .A(n2041), .B(n2038), .Z(n2040) );
  XOR U1816 ( .A(n2042), .B(n2043), .Z(n2030) );
  AND U1817 ( .A(n2044), .B(n2045), .Z(n2043) );
  XOR U1818 ( .A(n2042), .B(n1169), .Z(n2045) );
  XOR U1819 ( .A(n2046), .B(n2047), .Z(n1169) );
  AND U1820 ( .A(n230), .B(n2048), .Z(n2047) );
  XOR U1821 ( .A(n2049), .B(n2046), .Z(n2048) );
  XNOR U1822 ( .A(n1166), .B(n2042), .Z(n2044) );
  XOR U1823 ( .A(n2050), .B(n2051), .Z(n1166) );
  AND U1824 ( .A(n227), .B(n2052), .Z(n2051) );
  XOR U1825 ( .A(n2053), .B(n2050), .Z(n2052) );
  XOR U1826 ( .A(n2054), .B(n2055), .Z(n2042) );
  AND U1827 ( .A(n2056), .B(n2057), .Z(n2055) );
  XOR U1828 ( .A(n2054), .B(n1181), .Z(n2057) );
  XOR U1829 ( .A(n2058), .B(n2059), .Z(n1181) );
  AND U1830 ( .A(n230), .B(n2060), .Z(n2059) );
  XOR U1831 ( .A(n2061), .B(n2058), .Z(n2060) );
  XNOR U1832 ( .A(n1178), .B(n2054), .Z(n2056) );
  XOR U1833 ( .A(n2062), .B(n2063), .Z(n1178) );
  AND U1834 ( .A(n227), .B(n2064), .Z(n2063) );
  XOR U1835 ( .A(n2065), .B(n2062), .Z(n2064) );
  XOR U1836 ( .A(n2066), .B(n2067), .Z(n2054) );
  AND U1837 ( .A(n2068), .B(n2069), .Z(n2067) );
  XOR U1838 ( .A(n2066), .B(n1193), .Z(n2069) );
  XOR U1839 ( .A(n2070), .B(n2071), .Z(n1193) );
  AND U1840 ( .A(n230), .B(n2072), .Z(n2071) );
  XOR U1841 ( .A(n2073), .B(n2070), .Z(n2072) );
  XNOR U1842 ( .A(n1190), .B(n2066), .Z(n2068) );
  XOR U1843 ( .A(n2074), .B(n2075), .Z(n1190) );
  AND U1844 ( .A(n227), .B(n2076), .Z(n2075) );
  XOR U1845 ( .A(n2077), .B(n2074), .Z(n2076) );
  XOR U1846 ( .A(n2078), .B(n2079), .Z(n2066) );
  AND U1847 ( .A(n2080), .B(n2081), .Z(n2079) );
  XOR U1848 ( .A(n2078), .B(n1205), .Z(n2081) );
  XOR U1849 ( .A(n2082), .B(n2083), .Z(n1205) );
  AND U1850 ( .A(n230), .B(n2084), .Z(n2083) );
  XOR U1851 ( .A(n2085), .B(n2082), .Z(n2084) );
  XNOR U1852 ( .A(n1202), .B(n2078), .Z(n2080) );
  XOR U1853 ( .A(n2086), .B(n2087), .Z(n1202) );
  AND U1854 ( .A(n227), .B(n2088), .Z(n2087) );
  XOR U1855 ( .A(n2089), .B(n2086), .Z(n2088) );
  XOR U1856 ( .A(n2090), .B(n2091), .Z(n2078) );
  AND U1857 ( .A(n2092), .B(n2093), .Z(n2091) );
  XOR U1858 ( .A(n2090), .B(n1217), .Z(n2093) );
  XOR U1859 ( .A(n2094), .B(n2095), .Z(n1217) );
  AND U1860 ( .A(n230), .B(n2096), .Z(n2095) );
  XOR U1861 ( .A(n2097), .B(n2094), .Z(n2096) );
  XNOR U1862 ( .A(n1214), .B(n2090), .Z(n2092) );
  XOR U1863 ( .A(n2098), .B(n2099), .Z(n1214) );
  AND U1864 ( .A(n227), .B(n2100), .Z(n2099) );
  XOR U1865 ( .A(n2101), .B(n2098), .Z(n2100) );
  XOR U1866 ( .A(n2102), .B(n2103), .Z(n2090) );
  AND U1867 ( .A(n2104), .B(n2105), .Z(n2103) );
  XOR U1868 ( .A(n2102), .B(n1229), .Z(n2105) );
  XOR U1869 ( .A(n2106), .B(n2107), .Z(n1229) );
  AND U1870 ( .A(n230), .B(n2108), .Z(n2107) );
  XOR U1871 ( .A(n2109), .B(n2106), .Z(n2108) );
  XNOR U1872 ( .A(n1226), .B(n2102), .Z(n2104) );
  XOR U1873 ( .A(n2110), .B(n2111), .Z(n1226) );
  AND U1874 ( .A(n227), .B(n2112), .Z(n2111) );
  XOR U1875 ( .A(n2113), .B(n2110), .Z(n2112) );
  XOR U1876 ( .A(n2114), .B(n2115), .Z(n2102) );
  AND U1877 ( .A(n2116), .B(n2117), .Z(n2115) );
  XOR U1878 ( .A(n2114), .B(n1241), .Z(n2117) );
  XOR U1879 ( .A(n2118), .B(n2119), .Z(n1241) );
  AND U1880 ( .A(n230), .B(n2120), .Z(n2119) );
  XOR U1881 ( .A(n2121), .B(n2118), .Z(n2120) );
  XNOR U1882 ( .A(n1238), .B(n2114), .Z(n2116) );
  XOR U1883 ( .A(n2122), .B(n2123), .Z(n1238) );
  AND U1884 ( .A(n227), .B(n2124), .Z(n2123) );
  XOR U1885 ( .A(n2125), .B(n2122), .Z(n2124) );
  XOR U1886 ( .A(n2126), .B(n2127), .Z(n2114) );
  AND U1887 ( .A(n2128), .B(n2129), .Z(n2127) );
  XOR U1888 ( .A(n2126), .B(n1253), .Z(n2129) );
  XOR U1889 ( .A(n2130), .B(n2131), .Z(n1253) );
  AND U1890 ( .A(n230), .B(n2132), .Z(n2131) );
  XOR U1891 ( .A(n2133), .B(n2130), .Z(n2132) );
  XNOR U1892 ( .A(n1250), .B(n2126), .Z(n2128) );
  XOR U1893 ( .A(n2134), .B(n2135), .Z(n1250) );
  AND U1894 ( .A(n227), .B(n2136), .Z(n2135) );
  XOR U1895 ( .A(n2137), .B(n2134), .Z(n2136) );
  XOR U1896 ( .A(n2138), .B(n2139), .Z(n2126) );
  AND U1897 ( .A(n2140), .B(n2141), .Z(n2139) );
  XOR U1898 ( .A(n2138), .B(n1265), .Z(n2141) );
  XOR U1899 ( .A(n2142), .B(n2143), .Z(n1265) );
  AND U1900 ( .A(n230), .B(n2144), .Z(n2143) );
  XOR U1901 ( .A(n2145), .B(n2142), .Z(n2144) );
  XNOR U1902 ( .A(n1262), .B(n2138), .Z(n2140) );
  XOR U1903 ( .A(n2146), .B(n2147), .Z(n1262) );
  AND U1904 ( .A(n227), .B(n2148), .Z(n2147) );
  XOR U1905 ( .A(n2149), .B(n2146), .Z(n2148) );
  XOR U1906 ( .A(n2150), .B(n2151), .Z(n2138) );
  AND U1907 ( .A(n2152), .B(n2153), .Z(n2151) );
  XOR U1908 ( .A(n1277), .B(n2150), .Z(n2153) );
  XOR U1909 ( .A(n2154), .B(n2155), .Z(n1277) );
  AND U1910 ( .A(n230), .B(n2156), .Z(n2155) );
  XOR U1911 ( .A(n2154), .B(n2157), .Z(n2156) );
  XNOR U1912 ( .A(n2150), .B(n1274), .Z(n2152) );
  XOR U1913 ( .A(n2158), .B(n2159), .Z(n1274) );
  AND U1914 ( .A(n227), .B(n2160), .Z(n2159) );
  XOR U1915 ( .A(n2158), .B(n2161), .Z(n2160) );
  XOR U1916 ( .A(n2162), .B(n2163), .Z(n2150) );
  AND U1917 ( .A(n2164), .B(n2165), .Z(n2163) );
  XNOR U1918 ( .A(n2166), .B(n1290), .Z(n2165) );
  XOR U1919 ( .A(n2167), .B(n2168), .Z(n1290) );
  AND U1920 ( .A(n230), .B(n2169), .Z(n2168) );
  XOR U1921 ( .A(n2170), .B(n2167), .Z(n2169) );
  XNOR U1922 ( .A(n1287), .B(n2162), .Z(n2164) );
  XOR U1923 ( .A(n2171), .B(n2172), .Z(n1287) );
  AND U1924 ( .A(n227), .B(n2173), .Z(n2172) );
  XOR U1925 ( .A(n2174), .B(n2171), .Z(n2173) );
  IV U1926 ( .A(n2166), .Z(n2162) );
  AND U1927 ( .A(n1994), .B(n1997), .Z(n2166) );
  XNOR U1928 ( .A(n2175), .B(n2176), .Z(n1997) );
  AND U1929 ( .A(n230), .B(n2177), .Z(n2176) );
  XNOR U1930 ( .A(n2178), .B(n2175), .Z(n2177) );
  XOR U1931 ( .A(n2179), .B(n2180), .Z(n230) );
  AND U1932 ( .A(n2181), .B(n2182), .Z(n2180) );
  XNOR U1933 ( .A(n2002), .B(n2179), .Z(n2182) );
  AND U1934 ( .A(p_input[1919]), .B(p_input[1903]), .Z(n2002) );
  XOR U1935 ( .A(n2179), .B(n2003), .Z(n2181) );
  AND U1936 ( .A(p_input[1887]), .B(p_input[1871]), .Z(n2003) );
  XOR U1937 ( .A(n2183), .B(n2184), .Z(n2179) );
  AND U1938 ( .A(n2185), .B(n2186), .Z(n2184) );
  XOR U1939 ( .A(n2183), .B(n2013), .Z(n2186) );
  XNOR U1940 ( .A(p_input[1902]), .B(n2187), .Z(n2013) );
  AND U1941 ( .A(n114), .B(n2188), .Z(n2187) );
  XOR U1942 ( .A(p_input[1918]), .B(p_input[1902]), .Z(n2188) );
  XNOR U1943 ( .A(n2010), .B(n2183), .Z(n2185) );
  XOR U1944 ( .A(n2189), .B(n2190), .Z(n2010) );
  AND U1945 ( .A(n112), .B(n2191), .Z(n2190) );
  XOR U1946 ( .A(p_input[1886]), .B(p_input[1870]), .Z(n2191) );
  XOR U1947 ( .A(n2192), .B(n2193), .Z(n2183) );
  AND U1948 ( .A(n2194), .B(n2195), .Z(n2193) );
  XOR U1949 ( .A(n2192), .B(n2025), .Z(n2195) );
  XNOR U1950 ( .A(p_input[1901]), .B(n2196), .Z(n2025) );
  AND U1951 ( .A(n114), .B(n2197), .Z(n2196) );
  XOR U1952 ( .A(p_input[1917]), .B(p_input[1901]), .Z(n2197) );
  XNOR U1953 ( .A(n2022), .B(n2192), .Z(n2194) );
  XOR U1954 ( .A(n2198), .B(n2199), .Z(n2022) );
  AND U1955 ( .A(n112), .B(n2200), .Z(n2199) );
  XOR U1956 ( .A(p_input[1885]), .B(p_input[1869]), .Z(n2200) );
  XOR U1957 ( .A(n2201), .B(n2202), .Z(n2192) );
  AND U1958 ( .A(n2203), .B(n2204), .Z(n2202) );
  XOR U1959 ( .A(n2201), .B(n2037), .Z(n2204) );
  XNOR U1960 ( .A(p_input[1900]), .B(n2205), .Z(n2037) );
  AND U1961 ( .A(n114), .B(n2206), .Z(n2205) );
  XOR U1962 ( .A(p_input[1916]), .B(p_input[1900]), .Z(n2206) );
  XNOR U1963 ( .A(n2034), .B(n2201), .Z(n2203) );
  XOR U1964 ( .A(n2207), .B(n2208), .Z(n2034) );
  AND U1965 ( .A(n112), .B(n2209), .Z(n2208) );
  XOR U1966 ( .A(p_input[1884]), .B(p_input[1868]), .Z(n2209) );
  XOR U1967 ( .A(n2210), .B(n2211), .Z(n2201) );
  AND U1968 ( .A(n2212), .B(n2213), .Z(n2211) );
  XOR U1969 ( .A(n2210), .B(n2049), .Z(n2213) );
  XNOR U1970 ( .A(p_input[1899]), .B(n2214), .Z(n2049) );
  AND U1971 ( .A(n114), .B(n2215), .Z(n2214) );
  XOR U1972 ( .A(p_input[1915]), .B(p_input[1899]), .Z(n2215) );
  XNOR U1973 ( .A(n2046), .B(n2210), .Z(n2212) );
  XOR U1974 ( .A(n2216), .B(n2217), .Z(n2046) );
  AND U1975 ( .A(n112), .B(n2218), .Z(n2217) );
  XOR U1976 ( .A(p_input[1883]), .B(p_input[1867]), .Z(n2218) );
  XOR U1977 ( .A(n2219), .B(n2220), .Z(n2210) );
  AND U1978 ( .A(n2221), .B(n2222), .Z(n2220) );
  XOR U1979 ( .A(n2219), .B(n2061), .Z(n2222) );
  XNOR U1980 ( .A(p_input[1898]), .B(n2223), .Z(n2061) );
  AND U1981 ( .A(n114), .B(n2224), .Z(n2223) );
  XOR U1982 ( .A(p_input[1914]), .B(p_input[1898]), .Z(n2224) );
  XNOR U1983 ( .A(n2058), .B(n2219), .Z(n2221) );
  XOR U1984 ( .A(n2225), .B(n2226), .Z(n2058) );
  AND U1985 ( .A(n112), .B(n2227), .Z(n2226) );
  XOR U1986 ( .A(p_input[1882]), .B(p_input[1866]), .Z(n2227) );
  XOR U1987 ( .A(n2228), .B(n2229), .Z(n2219) );
  AND U1988 ( .A(n2230), .B(n2231), .Z(n2229) );
  XOR U1989 ( .A(n2228), .B(n2073), .Z(n2231) );
  XNOR U1990 ( .A(p_input[1897]), .B(n2232), .Z(n2073) );
  AND U1991 ( .A(n114), .B(n2233), .Z(n2232) );
  XOR U1992 ( .A(p_input[1913]), .B(p_input[1897]), .Z(n2233) );
  XNOR U1993 ( .A(n2070), .B(n2228), .Z(n2230) );
  XOR U1994 ( .A(n2234), .B(n2235), .Z(n2070) );
  AND U1995 ( .A(n112), .B(n2236), .Z(n2235) );
  XOR U1996 ( .A(p_input[1881]), .B(p_input[1865]), .Z(n2236) );
  XOR U1997 ( .A(n2237), .B(n2238), .Z(n2228) );
  AND U1998 ( .A(n2239), .B(n2240), .Z(n2238) );
  XOR U1999 ( .A(n2237), .B(n2085), .Z(n2240) );
  XNOR U2000 ( .A(p_input[1896]), .B(n2241), .Z(n2085) );
  AND U2001 ( .A(n114), .B(n2242), .Z(n2241) );
  XOR U2002 ( .A(p_input[1912]), .B(p_input[1896]), .Z(n2242) );
  XNOR U2003 ( .A(n2082), .B(n2237), .Z(n2239) );
  XOR U2004 ( .A(n2243), .B(n2244), .Z(n2082) );
  AND U2005 ( .A(n112), .B(n2245), .Z(n2244) );
  XOR U2006 ( .A(p_input[1880]), .B(p_input[1864]), .Z(n2245) );
  XOR U2007 ( .A(n2246), .B(n2247), .Z(n2237) );
  AND U2008 ( .A(n2248), .B(n2249), .Z(n2247) );
  XOR U2009 ( .A(n2246), .B(n2097), .Z(n2249) );
  XNOR U2010 ( .A(p_input[1895]), .B(n2250), .Z(n2097) );
  AND U2011 ( .A(n114), .B(n2251), .Z(n2250) );
  XOR U2012 ( .A(p_input[1911]), .B(p_input[1895]), .Z(n2251) );
  XNOR U2013 ( .A(n2094), .B(n2246), .Z(n2248) );
  XOR U2014 ( .A(n2252), .B(n2253), .Z(n2094) );
  AND U2015 ( .A(n112), .B(n2254), .Z(n2253) );
  XOR U2016 ( .A(p_input[1879]), .B(p_input[1863]), .Z(n2254) );
  XOR U2017 ( .A(n2255), .B(n2256), .Z(n2246) );
  AND U2018 ( .A(n2257), .B(n2258), .Z(n2256) );
  XOR U2019 ( .A(n2255), .B(n2109), .Z(n2258) );
  XNOR U2020 ( .A(p_input[1894]), .B(n2259), .Z(n2109) );
  AND U2021 ( .A(n114), .B(n2260), .Z(n2259) );
  XOR U2022 ( .A(p_input[1910]), .B(p_input[1894]), .Z(n2260) );
  XNOR U2023 ( .A(n2106), .B(n2255), .Z(n2257) );
  XOR U2024 ( .A(n2261), .B(n2262), .Z(n2106) );
  AND U2025 ( .A(n112), .B(n2263), .Z(n2262) );
  XOR U2026 ( .A(p_input[1878]), .B(p_input[1862]), .Z(n2263) );
  XOR U2027 ( .A(n2264), .B(n2265), .Z(n2255) );
  AND U2028 ( .A(n2266), .B(n2267), .Z(n2265) );
  XOR U2029 ( .A(n2264), .B(n2121), .Z(n2267) );
  XNOR U2030 ( .A(p_input[1893]), .B(n2268), .Z(n2121) );
  AND U2031 ( .A(n114), .B(n2269), .Z(n2268) );
  XOR U2032 ( .A(p_input[1909]), .B(p_input[1893]), .Z(n2269) );
  XNOR U2033 ( .A(n2118), .B(n2264), .Z(n2266) );
  XOR U2034 ( .A(n2270), .B(n2271), .Z(n2118) );
  AND U2035 ( .A(n112), .B(n2272), .Z(n2271) );
  XOR U2036 ( .A(p_input[1877]), .B(p_input[1861]), .Z(n2272) );
  XOR U2037 ( .A(n2273), .B(n2274), .Z(n2264) );
  AND U2038 ( .A(n2275), .B(n2276), .Z(n2274) );
  XOR U2039 ( .A(n2273), .B(n2133), .Z(n2276) );
  XNOR U2040 ( .A(p_input[1892]), .B(n2277), .Z(n2133) );
  AND U2041 ( .A(n114), .B(n2278), .Z(n2277) );
  XOR U2042 ( .A(p_input[1908]), .B(p_input[1892]), .Z(n2278) );
  XNOR U2043 ( .A(n2130), .B(n2273), .Z(n2275) );
  XOR U2044 ( .A(n2279), .B(n2280), .Z(n2130) );
  AND U2045 ( .A(n112), .B(n2281), .Z(n2280) );
  XOR U2046 ( .A(p_input[1876]), .B(p_input[1860]), .Z(n2281) );
  XOR U2047 ( .A(n2282), .B(n2283), .Z(n2273) );
  AND U2048 ( .A(n2284), .B(n2285), .Z(n2283) );
  XOR U2049 ( .A(n2282), .B(n2145), .Z(n2285) );
  XNOR U2050 ( .A(p_input[1891]), .B(n2286), .Z(n2145) );
  AND U2051 ( .A(n114), .B(n2287), .Z(n2286) );
  XOR U2052 ( .A(p_input[1907]), .B(p_input[1891]), .Z(n2287) );
  XNOR U2053 ( .A(n2142), .B(n2282), .Z(n2284) );
  XOR U2054 ( .A(n2288), .B(n2289), .Z(n2142) );
  AND U2055 ( .A(n112), .B(n2290), .Z(n2289) );
  XOR U2056 ( .A(p_input[1875]), .B(p_input[1859]), .Z(n2290) );
  XOR U2057 ( .A(n2291), .B(n2292), .Z(n2282) );
  AND U2058 ( .A(n2293), .B(n2294), .Z(n2292) );
  XOR U2059 ( .A(n2157), .B(n2291), .Z(n2294) );
  XNOR U2060 ( .A(p_input[1890]), .B(n2295), .Z(n2157) );
  AND U2061 ( .A(n114), .B(n2296), .Z(n2295) );
  XOR U2062 ( .A(p_input[1906]), .B(p_input[1890]), .Z(n2296) );
  XNOR U2063 ( .A(n2291), .B(n2154), .Z(n2293) );
  XOR U2064 ( .A(n2297), .B(n2298), .Z(n2154) );
  AND U2065 ( .A(n112), .B(n2299), .Z(n2298) );
  XOR U2066 ( .A(p_input[1874]), .B(p_input[1858]), .Z(n2299) );
  XOR U2067 ( .A(n2300), .B(n2301), .Z(n2291) );
  AND U2068 ( .A(n2302), .B(n2303), .Z(n2301) );
  XNOR U2069 ( .A(n2304), .B(n2170), .Z(n2303) );
  XNOR U2070 ( .A(p_input[1889]), .B(n2305), .Z(n2170) );
  AND U2071 ( .A(n114), .B(n2306), .Z(n2305) );
  XNOR U2072 ( .A(p_input[1905]), .B(n2307), .Z(n2306) );
  IV U2073 ( .A(p_input[1889]), .Z(n2307) );
  XNOR U2074 ( .A(n2167), .B(n2300), .Z(n2302) );
  XNOR U2075 ( .A(p_input[1857]), .B(n2308), .Z(n2167) );
  AND U2076 ( .A(n112), .B(n2309), .Z(n2308) );
  XOR U2077 ( .A(p_input[1873]), .B(p_input[1857]), .Z(n2309) );
  IV U2078 ( .A(n2304), .Z(n2300) );
  AND U2079 ( .A(n2175), .B(n2178), .Z(n2304) );
  XOR U2080 ( .A(p_input[1888]), .B(n2310), .Z(n2178) );
  AND U2081 ( .A(n114), .B(n2311), .Z(n2310) );
  XOR U2082 ( .A(p_input[1904]), .B(p_input[1888]), .Z(n2311) );
  XOR U2083 ( .A(n2312), .B(n2313), .Z(n114) );
  AND U2084 ( .A(n2314), .B(n2315), .Z(n2313) );
  XNOR U2085 ( .A(p_input[1919]), .B(n2312), .Z(n2315) );
  XOR U2086 ( .A(n2312), .B(p_input[1903]), .Z(n2314) );
  XOR U2087 ( .A(n2316), .B(n2317), .Z(n2312) );
  AND U2088 ( .A(n2318), .B(n2319), .Z(n2317) );
  XNOR U2089 ( .A(p_input[1918]), .B(n2316), .Z(n2319) );
  XOR U2090 ( .A(n2316), .B(p_input[1902]), .Z(n2318) );
  XOR U2091 ( .A(n2320), .B(n2321), .Z(n2316) );
  AND U2092 ( .A(n2322), .B(n2323), .Z(n2321) );
  XNOR U2093 ( .A(p_input[1917]), .B(n2320), .Z(n2323) );
  XOR U2094 ( .A(n2320), .B(p_input[1901]), .Z(n2322) );
  XOR U2095 ( .A(n2324), .B(n2325), .Z(n2320) );
  AND U2096 ( .A(n2326), .B(n2327), .Z(n2325) );
  XNOR U2097 ( .A(p_input[1916]), .B(n2324), .Z(n2327) );
  XOR U2098 ( .A(n2324), .B(p_input[1900]), .Z(n2326) );
  XOR U2099 ( .A(n2328), .B(n2329), .Z(n2324) );
  AND U2100 ( .A(n2330), .B(n2331), .Z(n2329) );
  XNOR U2101 ( .A(p_input[1915]), .B(n2328), .Z(n2331) );
  XOR U2102 ( .A(n2328), .B(p_input[1899]), .Z(n2330) );
  XOR U2103 ( .A(n2332), .B(n2333), .Z(n2328) );
  AND U2104 ( .A(n2334), .B(n2335), .Z(n2333) );
  XNOR U2105 ( .A(p_input[1914]), .B(n2332), .Z(n2335) );
  XOR U2106 ( .A(n2332), .B(p_input[1898]), .Z(n2334) );
  XOR U2107 ( .A(n2336), .B(n2337), .Z(n2332) );
  AND U2108 ( .A(n2338), .B(n2339), .Z(n2337) );
  XNOR U2109 ( .A(p_input[1913]), .B(n2336), .Z(n2339) );
  XOR U2110 ( .A(n2336), .B(p_input[1897]), .Z(n2338) );
  XOR U2111 ( .A(n2340), .B(n2341), .Z(n2336) );
  AND U2112 ( .A(n2342), .B(n2343), .Z(n2341) );
  XNOR U2113 ( .A(p_input[1912]), .B(n2340), .Z(n2343) );
  XOR U2114 ( .A(n2340), .B(p_input[1896]), .Z(n2342) );
  XOR U2115 ( .A(n2344), .B(n2345), .Z(n2340) );
  AND U2116 ( .A(n2346), .B(n2347), .Z(n2345) );
  XNOR U2117 ( .A(p_input[1911]), .B(n2344), .Z(n2347) );
  XOR U2118 ( .A(n2344), .B(p_input[1895]), .Z(n2346) );
  XOR U2119 ( .A(n2348), .B(n2349), .Z(n2344) );
  AND U2120 ( .A(n2350), .B(n2351), .Z(n2349) );
  XNOR U2121 ( .A(p_input[1910]), .B(n2348), .Z(n2351) );
  XOR U2122 ( .A(n2348), .B(p_input[1894]), .Z(n2350) );
  XOR U2123 ( .A(n2352), .B(n2353), .Z(n2348) );
  AND U2124 ( .A(n2354), .B(n2355), .Z(n2353) );
  XNOR U2125 ( .A(p_input[1909]), .B(n2352), .Z(n2355) );
  XOR U2126 ( .A(n2352), .B(p_input[1893]), .Z(n2354) );
  XOR U2127 ( .A(n2356), .B(n2357), .Z(n2352) );
  AND U2128 ( .A(n2358), .B(n2359), .Z(n2357) );
  XNOR U2129 ( .A(p_input[1908]), .B(n2356), .Z(n2359) );
  XOR U2130 ( .A(n2356), .B(p_input[1892]), .Z(n2358) );
  XOR U2131 ( .A(n2360), .B(n2361), .Z(n2356) );
  AND U2132 ( .A(n2362), .B(n2363), .Z(n2361) );
  XNOR U2133 ( .A(p_input[1907]), .B(n2360), .Z(n2363) );
  XOR U2134 ( .A(n2360), .B(p_input[1891]), .Z(n2362) );
  XOR U2135 ( .A(n2364), .B(n2365), .Z(n2360) );
  AND U2136 ( .A(n2366), .B(n2367), .Z(n2365) );
  XNOR U2137 ( .A(p_input[1906]), .B(n2364), .Z(n2367) );
  XOR U2138 ( .A(n2364), .B(p_input[1890]), .Z(n2366) );
  XNOR U2139 ( .A(n2368), .B(n2369), .Z(n2364) );
  AND U2140 ( .A(n2370), .B(n2371), .Z(n2369) );
  XOR U2141 ( .A(p_input[1905]), .B(n2368), .Z(n2371) );
  XNOR U2142 ( .A(p_input[1889]), .B(n2368), .Z(n2370) );
  AND U2143 ( .A(p_input[1904]), .B(n2372), .Z(n2368) );
  IV U2144 ( .A(p_input[1888]), .Z(n2372) );
  XNOR U2145 ( .A(p_input[1856]), .B(n2373), .Z(n2175) );
  AND U2146 ( .A(n112), .B(n2374), .Z(n2373) );
  XOR U2147 ( .A(p_input[1872]), .B(p_input[1856]), .Z(n2374) );
  XOR U2148 ( .A(n2375), .B(n2376), .Z(n112) );
  AND U2149 ( .A(n2377), .B(n2378), .Z(n2376) );
  XNOR U2150 ( .A(p_input[1887]), .B(n2375), .Z(n2378) );
  XOR U2151 ( .A(n2375), .B(p_input[1871]), .Z(n2377) );
  XOR U2152 ( .A(n2379), .B(n2380), .Z(n2375) );
  AND U2153 ( .A(n2381), .B(n2382), .Z(n2380) );
  XNOR U2154 ( .A(p_input[1886]), .B(n2379), .Z(n2382) );
  XNOR U2155 ( .A(n2379), .B(n2189), .Z(n2381) );
  IV U2156 ( .A(p_input[1870]), .Z(n2189) );
  XOR U2157 ( .A(n2383), .B(n2384), .Z(n2379) );
  AND U2158 ( .A(n2385), .B(n2386), .Z(n2384) );
  XNOR U2159 ( .A(p_input[1885]), .B(n2383), .Z(n2386) );
  XNOR U2160 ( .A(n2383), .B(n2198), .Z(n2385) );
  IV U2161 ( .A(p_input[1869]), .Z(n2198) );
  XOR U2162 ( .A(n2387), .B(n2388), .Z(n2383) );
  AND U2163 ( .A(n2389), .B(n2390), .Z(n2388) );
  XNOR U2164 ( .A(p_input[1884]), .B(n2387), .Z(n2390) );
  XNOR U2165 ( .A(n2387), .B(n2207), .Z(n2389) );
  IV U2166 ( .A(p_input[1868]), .Z(n2207) );
  XOR U2167 ( .A(n2391), .B(n2392), .Z(n2387) );
  AND U2168 ( .A(n2393), .B(n2394), .Z(n2392) );
  XNOR U2169 ( .A(p_input[1883]), .B(n2391), .Z(n2394) );
  XNOR U2170 ( .A(n2391), .B(n2216), .Z(n2393) );
  IV U2171 ( .A(p_input[1867]), .Z(n2216) );
  XOR U2172 ( .A(n2395), .B(n2396), .Z(n2391) );
  AND U2173 ( .A(n2397), .B(n2398), .Z(n2396) );
  XNOR U2174 ( .A(p_input[1882]), .B(n2395), .Z(n2398) );
  XNOR U2175 ( .A(n2395), .B(n2225), .Z(n2397) );
  IV U2176 ( .A(p_input[1866]), .Z(n2225) );
  XOR U2177 ( .A(n2399), .B(n2400), .Z(n2395) );
  AND U2178 ( .A(n2401), .B(n2402), .Z(n2400) );
  XNOR U2179 ( .A(p_input[1881]), .B(n2399), .Z(n2402) );
  XNOR U2180 ( .A(n2399), .B(n2234), .Z(n2401) );
  IV U2181 ( .A(p_input[1865]), .Z(n2234) );
  XOR U2182 ( .A(n2403), .B(n2404), .Z(n2399) );
  AND U2183 ( .A(n2405), .B(n2406), .Z(n2404) );
  XNOR U2184 ( .A(p_input[1880]), .B(n2403), .Z(n2406) );
  XNOR U2185 ( .A(n2403), .B(n2243), .Z(n2405) );
  IV U2186 ( .A(p_input[1864]), .Z(n2243) );
  XOR U2187 ( .A(n2407), .B(n2408), .Z(n2403) );
  AND U2188 ( .A(n2409), .B(n2410), .Z(n2408) );
  XNOR U2189 ( .A(p_input[1879]), .B(n2407), .Z(n2410) );
  XNOR U2190 ( .A(n2407), .B(n2252), .Z(n2409) );
  IV U2191 ( .A(p_input[1863]), .Z(n2252) );
  XOR U2192 ( .A(n2411), .B(n2412), .Z(n2407) );
  AND U2193 ( .A(n2413), .B(n2414), .Z(n2412) );
  XNOR U2194 ( .A(p_input[1878]), .B(n2411), .Z(n2414) );
  XNOR U2195 ( .A(n2411), .B(n2261), .Z(n2413) );
  IV U2196 ( .A(p_input[1862]), .Z(n2261) );
  XOR U2197 ( .A(n2415), .B(n2416), .Z(n2411) );
  AND U2198 ( .A(n2417), .B(n2418), .Z(n2416) );
  XNOR U2199 ( .A(p_input[1877]), .B(n2415), .Z(n2418) );
  XNOR U2200 ( .A(n2415), .B(n2270), .Z(n2417) );
  IV U2201 ( .A(p_input[1861]), .Z(n2270) );
  XOR U2202 ( .A(n2419), .B(n2420), .Z(n2415) );
  AND U2203 ( .A(n2421), .B(n2422), .Z(n2420) );
  XNOR U2204 ( .A(p_input[1876]), .B(n2419), .Z(n2422) );
  XNOR U2205 ( .A(n2419), .B(n2279), .Z(n2421) );
  IV U2206 ( .A(p_input[1860]), .Z(n2279) );
  XOR U2207 ( .A(n2423), .B(n2424), .Z(n2419) );
  AND U2208 ( .A(n2425), .B(n2426), .Z(n2424) );
  XNOR U2209 ( .A(p_input[1875]), .B(n2423), .Z(n2426) );
  XNOR U2210 ( .A(n2423), .B(n2288), .Z(n2425) );
  IV U2211 ( .A(p_input[1859]), .Z(n2288) );
  XOR U2212 ( .A(n2427), .B(n2428), .Z(n2423) );
  AND U2213 ( .A(n2429), .B(n2430), .Z(n2428) );
  XNOR U2214 ( .A(p_input[1874]), .B(n2427), .Z(n2430) );
  XNOR U2215 ( .A(n2427), .B(n2297), .Z(n2429) );
  IV U2216 ( .A(p_input[1858]), .Z(n2297) );
  XNOR U2217 ( .A(n2431), .B(n2432), .Z(n2427) );
  AND U2218 ( .A(n2433), .B(n2434), .Z(n2432) );
  XOR U2219 ( .A(p_input[1873]), .B(n2431), .Z(n2434) );
  XNOR U2220 ( .A(p_input[1857]), .B(n2431), .Z(n2433) );
  AND U2221 ( .A(p_input[1872]), .B(n2435), .Z(n2431) );
  IV U2222 ( .A(p_input[1856]), .Z(n2435) );
  XOR U2223 ( .A(n2436), .B(n2437), .Z(n1994) );
  AND U2224 ( .A(n227), .B(n2438), .Z(n2437) );
  XNOR U2225 ( .A(n2439), .B(n2436), .Z(n2438) );
  XOR U2226 ( .A(n2440), .B(n2441), .Z(n227) );
  AND U2227 ( .A(n2442), .B(n2443), .Z(n2441) );
  XNOR U2228 ( .A(n2005), .B(n2440), .Z(n2443) );
  AND U2229 ( .A(p_input[1855]), .B(p_input[1839]), .Z(n2005) );
  XOR U2230 ( .A(n2440), .B(n2004), .Z(n2442) );
  AND U2231 ( .A(p_input[1807]), .B(p_input[1823]), .Z(n2004) );
  XOR U2232 ( .A(n2444), .B(n2445), .Z(n2440) );
  AND U2233 ( .A(n2446), .B(n2447), .Z(n2445) );
  XOR U2234 ( .A(n2444), .B(n2017), .Z(n2447) );
  XNOR U2235 ( .A(p_input[1838]), .B(n2448), .Z(n2017) );
  AND U2236 ( .A(n118), .B(n2449), .Z(n2448) );
  XOR U2237 ( .A(p_input[1854]), .B(p_input[1838]), .Z(n2449) );
  XNOR U2238 ( .A(n2014), .B(n2444), .Z(n2446) );
  XOR U2239 ( .A(n2450), .B(n2451), .Z(n2014) );
  AND U2240 ( .A(n115), .B(n2452), .Z(n2451) );
  XOR U2241 ( .A(p_input[1822]), .B(p_input[1806]), .Z(n2452) );
  XOR U2242 ( .A(n2453), .B(n2454), .Z(n2444) );
  AND U2243 ( .A(n2455), .B(n2456), .Z(n2454) );
  XOR U2244 ( .A(n2453), .B(n2029), .Z(n2456) );
  XNOR U2245 ( .A(p_input[1837]), .B(n2457), .Z(n2029) );
  AND U2246 ( .A(n118), .B(n2458), .Z(n2457) );
  XOR U2247 ( .A(p_input[1853]), .B(p_input[1837]), .Z(n2458) );
  XNOR U2248 ( .A(n2026), .B(n2453), .Z(n2455) );
  XOR U2249 ( .A(n2459), .B(n2460), .Z(n2026) );
  AND U2250 ( .A(n115), .B(n2461), .Z(n2460) );
  XOR U2251 ( .A(p_input[1821]), .B(p_input[1805]), .Z(n2461) );
  XOR U2252 ( .A(n2462), .B(n2463), .Z(n2453) );
  AND U2253 ( .A(n2464), .B(n2465), .Z(n2463) );
  XOR U2254 ( .A(n2462), .B(n2041), .Z(n2465) );
  XNOR U2255 ( .A(p_input[1836]), .B(n2466), .Z(n2041) );
  AND U2256 ( .A(n118), .B(n2467), .Z(n2466) );
  XOR U2257 ( .A(p_input[1852]), .B(p_input[1836]), .Z(n2467) );
  XNOR U2258 ( .A(n2038), .B(n2462), .Z(n2464) );
  XOR U2259 ( .A(n2468), .B(n2469), .Z(n2038) );
  AND U2260 ( .A(n115), .B(n2470), .Z(n2469) );
  XOR U2261 ( .A(p_input[1820]), .B(p_input[1804]), .Z(n2470) );
  XOR U2262 ( .A(n2471), .B(n2472), .Z(n2462) );
  AND U2263 ( .A(n2473), .B(n2474), .Z(n2472) );
  XOR U2264 ( .A(n2471), .B(n2053), .Z(n2474) );
  XNOR U2265 ( .A(p_input[1835]), .B(n2475), .Z(n2053) );
  AND U2266 ( .A(n118), .B(n2476), .Z(n2475) );
  XOR U2267 ( .A(p_input[1851]), .B(p_input[1835]), .Z(n2476) );
  XNOR U2268 ( .A(n2050), .B(n2471), .Z(n2473) );
  XOR U2269 ( .A(n2477), .B(n2478), .Z(n2050) );
  AND U2270 ( .A(n115), .B(n2479), .Z(n2478) );
  XOR U2271 ( .A(p_input[1819]), .B(p_input[1803]), .Z(n2479) );
  XOR U2272 ( .A(n2480), .B(n2481), .Z(n2471) );
  AND U2273 ( .A(n2482), .B(n2483), .Z(n2481) );
  XOR U2274 ( .A(n2480), .B(n2065), .Z(n2483) );
  XNOR U2275 ( .A(p_input[1834]), .B(n2484), .Z(n2065) );
  AND U2276 ( .A(n118), .B(n2485), .Z(n2484) );
  XOR U2277 ( .A(p_input[1850]), .B(p_input[1834]), .Z(n2485) );
  XNOR U2278 ( .A(n2062), .B(n2480), .Z(n2482) );
  XOR U2279 ( .A(n2486), .B(n2487), .Z(n2062) );
  AND U2280 ( .A(n115), .B(n2488), .Z(n2487) );
  XOR U2281 ( .A(p_input[1818]), .B(p_input[1802]), .Z(n2488) );
  XOR U2282 ( .A(n2489), .B(n2490), .Z(n2480) );
  AND U2283 ( .A(n2491), .B(n2492), .Z(n2490) );
  XOR U2284 ( .A(n2489), .B(n2077), .Z(n2492) );
  XNOR U2285 ( .A(p_input[1833]), .B(n2493), .Z(n2077) );
  AND U2286 ( .A(n118), .B(n2494), .Z(n2493) );
  XOR U2287 ( .A(p_input[1849]), .B(p_input[1833]), .Z(n2494) );
  XNOR U2288 ( .A(n2074), .B(n2489), .Z(n2491) );
  XOR U2289 ( .A(n2495), .B(n2496), .Z(n2074) );
  AND U2290 ( .A(n115), .B(n2497), .Z(n2496) );
  XOR U2291 ( .A(p_input[1817]), .B(p_input[1801]), .Z(n2497) );
  XOR U2292 ( .A(n2498), .B(n2499), .Z(n2489) );
  AND U2293 ( .A(n2500), .B(n2501), .Z(n2499) );
  XOR U2294 ( .A(n2498), .B(n2089), .Z(n2501) );
  XNOR U2295 ( .A(p_input[1832]), .B(n2502), .Z(n2089) );
  AND U2296 ( .A(n118), .B(n2503), .Z(n2502) );
  XOR U2297 ( .A(p_input[1848]), .B(p_input[1832]), .Z(n2503) );
  XNOR U2298 ( .A(n2086), .B(n2498), .Z(n2500) );
  XOR U2299 ( .A(n2504), .B(n2505), .Z(n2086) );
  AND U2300 ( .A(n115), .B(n2506), .Z(n2505) );
  XOR U2301 ( .A(p_input[1816]), .B(p_input[1800]), .Z(n2506) );
  XOR U2302 ( .A(n2507), .B(n2508), .Z(n2498) );
  AND U2303 ( .A(n2509), .B(n2510), .Z(n2508) );
  XOR U2304 ( .A(n2507), .B(n2101), .Z(n2510) );
  XNOR U2305 ( .A(p_input[1831]), .B(n2511), .Z(n2101) );
  AND U2306 ( .A(n118), .B(n2512), .Z(n2511) );
  XOR U2307 ( .A(p_input[1847]), .B(p_input[1831]), .Z(n2512) );
  XNOR U2308 ( .A(n2098), .B(n2507), .Z(n2509) );
  XOR U2309 ( .A(n2513), .B(n2514), .Z(n2098) );
  AND U2310 ( .A(n115), .B(n2515), .Z(n2514) );
  XOR U2311 ( .A(p_input[1815]), .B(p_input[1799]), .Z(n2515) );
  XOR U2312 ( .A(n2516), .B(n2517), .Z(n2507) );
  AND U2313 ( .A(n2518), .B(n2519), .Z(n2517) );
  XOR U2314 ( .A(n2516), .B(n2113), .Z(n2519) );
  XNOR U2315 ( .A(p_input[1830]), .B(n2520), .Z(n2113) );
  AND U2316 ( .A(n118), .B(n2521), .Z(n2520) );
  XOR U2317 ( .A(p_input[1846]), .B(p_input[1830]), .Z(n2521) );
  XNOR U2318 ( .A(n2110), .B(n2516), .Z(n2518) );
  XOR U2319 ( .A(n2522), .B(n2523), .Z(n2110) );
  AND U2320 ( .A(n115), .B(n2524), .Z(n2523) );
  XOR U2321 ( .A(p_input[1814]), .B(p_input[1798]), .Z(n2524) );
  XOR U2322 ( .A(n2525), .B(n2526), .Z(n2516) );
  AND U2323 ( .A(n2527), .B(n2528), .Z(n2526) );
  XOR U2324 ( .A(n2525), .B(n2125), .Z(n2528) );
  XNOR U2325 ( .A(p_input[1829]), .B(n2529), .Z(n2125) );
  AND U2326 ( .A(n118), .B(n2530), .Z(n2529) );
  XOR U2327 ( .A(p_input[1845]), .B(p_input[1829]), .Z(n2530) );
  XNOR U2328 ( .A(n2122), .B(n2525), .Z(n2527) );
  XOR U2329 ( .A(n2531), .B(n2532), .Z(n2122) );
  AND U2330 ( .A(n115), .B(n2533), .Z(n2532) );
  XOR U2331 ( .A(p_input[1813]), .B(p_input[1797]), .Z(n2533) );
  XOR U2332 ( .A(n2534), .B(n2535), .Z(n2525) );
  AND U2333 ( .A(n2536), .B(n2537), .Z(n2535) );
  XOR U2334 ( .A(n2534), .B(n2137), .Z(n2537) );
  XNOR U2335 ( .A(p_input[1828]), .B(n2538), .Z(n2137) );
  AND U2336 ( .A(n118), .B(n2539), .Z(n2538) );
  XOR U2337 ( .A(p_input[1844]), .B(p_input[1828]), .Z(n2539) );
  XNOR U2338 ( .A(n2134), .B(n2534), .Z(n2536) );
  XOR U2339 ( .A(n2540), .B(n2541), .Z(n2134) );
  AND U2340 ( .A(n115), .B(n2542), .Z(n2541) );
  XOR U2341 ( .A(p_input[1812]), .B(p_input[1796]), .Z(n2542) );
  XOR U2342 ( .A(n2543), .B(n2544), .Z(n2534) );
  AND U2343 ( .A(n2545), .B(n2546), .Z(n2544) );
  XOR U2344 ( .A(n2543), .B(n2149), .Z(n2546) );
  XNOR U2345 ( .A(p_input[1827]), .B(n2547), .Z(n2149) );
  AND U2346 ( .A(n118), .B(n2548), .Z(n2547) );
  XOR U2347 ( .A(p_input[1843]), .B(p_input[1827]), .Z(n2548) );
  XNOR U2348 ( .A(n2146), .B(n2543), .Z(n2545) );
  XOR U2349 ( .A(n2549), .B(n2550), .Z(n2146) );
  AND U2350 ( .A(n115), .B(n2551), .Z(n2550) );
  XOR U2351 ( .A(p_input[1811]), .B(p_input[1795]), .Z(n2551) );
  XOR U2352 ( .A(n2552), .B(n2553), .Z(n2543) );
  AND U2353 ( .A(n2554), .B(n2555), .Z(n2553) );
  XOR U2354 ( .A(n2161), .B(n2552), .Z(n2555) );
  XNOR U2355 ( .A(p_input[1826]), .B(n2556), .Z(n2161) );
  AND U2356 ( .A(n118), .B(n2557), .Z(n2556) );
  XOR U2357 ( .A(p_input[1842]), .B(p_input[1826]), .Z(n2557) );
  XNOR U2358 ( .A(n2552), .B(n2158), .Z(n2554) );
  XOR U2359 ( .A(n2558), .B(n2559), .Z(n2158) );
  AND U2360 ( .A(n115), .B(n2560), .Z(n2559) );
  XOR U2361 ( .A(p_input[1810]), .B(p_input[1794]), .Z(n2560) );
  XOR U2362 ( .A(n2561), .B(n2562), .Z(n2552) );
  AND U2363 ( .A(n2563), .B(n2564), .Z(n2562) );
  XNOR U2364 ( .A(n2565), .B(n2174), .Z(n2564) );
  XNOR U2365 ( .A(p_input[1825]), .B(n2566), .Z(n2174) );
  AND U2366 ( .A(n118), .B(n2567), .Z(n2566) );
  XNOR U2367 ( .A(p_input[1841]), .B(n2568), .Z(n2567) );
  IV U2368 ( .A(p_input[1825]), .Z(n2568) );
  XNOR U2369 ( .A(n2171), .B(n2561), .Z(n2563) );
  XNOR U2370 ( .A(p_input[1793]), .B(n2569), .Z(n2171) );
  AND U2371 ( .A(n115), .B(n2570), .Z(n2569) );
  XOR U2372 ( .A(p_input[1809]), .B(p_input[1793]), .Z(n2570) );
  IV U2373 ( .A(n2565), .Z(n2561) );
  AND U2374 ( .A(n2436), .B(n2439), .Z(n2565) );
  XOR U2375 ( .A(p_input[1824]), .B(n2571), .Z(n2439) );
  AND U2376 ( .A(n118), .B(n2572), .Z(n2571) );
  XOR U2377 ( .A(p_input[1840]), .B(p_input[1824]), .Z(n2572) );
  XOR U2378 ( .A(n2573), .B(n2574), .Z(n118) );
  AND U2379 ( .A(n2575), .B(n2576), .Z(n2574) );
  XNOR U2380 ( .A(p_input[1855]), .B(n2573), .Z(n2576) );
  XOR U2381 ( .A(n2573), .B(p_input[1839]), .Z(n2575) );
  XOR U2382 ( .A(n2577), .B(n2578), .Z(n2573) );
  AND U2383 ( .A(n2579), .B(n2580), .Z(n2578) );
  XNOR U2384 ( .A(p_input[1854]), .B(n2577), .Z(n2580) );
  XOR U2385 ( .A(n2577), .B(p_input[1838]), .Z(n2579) );
  XOR U2386 ( .A(n2581), .B(n2582), .Z(n2577) );
  AND U2387 ( .A(n2583), .B(n2584), .Z(n2582) );
  XNOR U2388 ( .A(p_input[1853]), .B(n2581), .Z(n2584) );
  XOR U2389 ( .A(n2581), .B(p_input[1837]), .Z(n2583) );
  XOR U2390 ( .A(n2585), .B(n2586), .Z(n2581) );
  AND U2391 ( .A(n2587), .B(n2588), .Z(n2586) );
  XNOR U2392 ( .A(p_input[1852]), .B(n2585), .Z(n2588) );
  XOR U2393 ( .A(n2585), .B(p_input[1836]), .Z(n2587) );
  XOR U2394 ( .A(n2589), .B(n2590), .Z(n2585) );
  AND U2395 ( .A(n2591), .B(n2592), .Z(n2590) );
  XNOR U2396 ( .A(p_input[1851]), .B(n2589), .Z(n2592) );
  XOR U2397 ( .A(n2589), .B(p_input[1835]), .Z(n2591) );
  XOR U2398 ( .A(n2593), .B(n2594), .Z(n2589) );
  AND U2399 ( .A(n2595), .B(n2596), .Z(n2594) );
  XNOR U2400 ( .A(p_input[1850]), .B(n2593), .Z(n2596) );
  XOR U2401 ( .A(n2593), .B(p_input[1834]), .Z(n2595) );
  XOR U2402 ( .A(n2597), .B(n2598), .Z(n2593) );
  AND U2403 ( .A(n2599), .B(n2600), .Z(n2598) );
  XNOR U2404 ( .A(p_input[1849]), .B(n2597), .Z(n2600) );
  XOR U2405 ( .A(n2597), .B(p_input[1833]), .Z(n2599) );
  XOR U2406 ( .A(n2601), .B(n2602), .Z(n2597) );
  AND U2407 ( .A(n2603), .B(n2604), .Z(n2602) );
  XNOR U2408 ( .A(p_input[1848]), .B(n2601), .Z(n2604) );
  XOR U2409 ( .A(n2601), .B(p_input[1832]), .Z(n2603) );
  XOR U2410 ( .A(n2605), .B(n2606), .Z(n2601) );
  AND U2411 ( .A(n2607), .B(n2608), .Z(n2606) );
  XNOR U2412 ( .A(p_input[1847]), .B(n2605), .Z(n2608) );
  XOR U2413 ( .A(n2605), .B(p_input[1831]), .Z(n2607) );
  XOR U2414 ( .A(n2609), .B(n2610), .Z(n2605) );
  AND U2415 ( .A(n2611), .B(n2612), .Z(n2610) );
  XNOR U2416 ( .A(p_input[1846]), .B(n2609), .Z(n2612) );
  XOR U2417 ( .A(n2609), .B(p_input[1830]), .Z(n2611) );
  XOR U2418 ( .A(n2613), .B(n2614), .Z(n2609) );
  AND U2419 ( .A(n2615), .B(n2616), .Z(n2614) );
  XNOR U2420 ( .A(p_input[1845]), .B(n2613), .Z(n2616) );
  XOR U2421 ( .A(n2613), .B(p_input[1829]), .Z(n2615) );
  XOR U2422 ( .A(n2617), .B(n2618), .Z(n2613) );
  AND U2423 ( .A(n2619), .B(n2620), .Z(n2618) );
  XNOR U2424 ( .A(p_input[1844]), .B(n2617), .Z(n2620) );
  XOR U2425 ( .A(n2617), .B(p_input[1828]), .Z(n2619) );
  XOR U2426 ( .A(n2621), .B(n2622), .Z(n2617) );
  AND U2427 ( .A(n2623), .B(n2624), .Z(n2622) );
  XNOR U2428 ( .A(p_input[1843]), .B(n2621), .Z(n2624) );
  XOR U2429 ( .A(n2621), .B(p_input[1827]), .Z(n2623) );
  XOR U2430 ( .A(n2625), .B(n2626), .Z(n2621) );
  AND U2431 ( .A(n2627), .B(n2628), .Z(n2626) );
  XNOR U2432 ( .A(p_input[1842]), .B(n2625), .Z(n2628) );
  XOR U2433 ( .A(n2625), .B(p_input[1826]), .Z(n2627) );
  XNOR U2434 ( .A(n2629), .B(n2630), .Z(n2625) );
  AND U2435 ( .A(n2631), .B(n2632), .Z(n2630) );
  XOR U2436 ( .A(p_input[1841]), .B(n2629), .Z(n2632) );
  XNOR U2437 ( .A(p_input[1825]), .B(n2629), .Z(n2631) );
  AND U2438 ( .A(p_input[1840]), .B(n2633), .Z(n2629) );
  IV U2439 ( .A(p_input[1824]), .Z(n2633) );
  XNOR U2440 ( .A(p_input[1792]), .B(n2634), .Z(n2436) );
  AND U2441 ( .A(n115), .B(n2635), .Z(n2634) );
  XOR U2442 ( .A(p_input[1808]), .B(p_input[1792]), .Z(n2635) );
  XOR U2443 ( .A(n2636), .B(n2637), .Z(n115) );
  AND U2444 ( .A(n2638), .B(n2639), .Z(n2637) );
  XNOR U2445 ( .A(p_input[1823]), .B(n2636), .Z(n2639) );
  XOR U2446 ( .A(n2636), .B(p_input[1807]), .Z(n2638) );
  XOR U2447 ( .A(n2640), .B(n2641), .Z(n2636) );
  AND U2448 ( .A(n2642), .B(n2643), .Z(n2641) );
  XNOR U2449 ( .A(p_input[1822]), .B(n2640), .Z(n2643) );
  XNOR U2450 ( .A(n2640), .B(n2450), .Z(n2642) );
  IV U2451 ( .A(p_input[1806]), .Z(n2450) );
  XOR U2452 ( .A(n2644), .B(n2645), .Z(n2640) );
  AND U2453 ( .A(n2646), .B(n2647), .Z(n2645) );
  XNOR U2454 ( .A(p_input[1821]), .B(n2644), .Z(n2647) );
  XNOR U2455 ( .A(n2644), .B(n2459), .Z(n2646) );
  IV U2456 ( .A(p_input[1805]), .Z(n2459) );
  XOR U2457 ( .A(n2648), .B(n2649), .Z(n2644) );
  AND U2458 ( .A(n2650), .B(n2651), .Z(n2649) );
  XNOR U2459 ( .A(p_input[1820]), .B(n2648), .Z(n2651) );
  XNOR U2460 ( .A(n2648), .B(n2468), .Z(n2650) );
  IV U2461 ( .A(p_input[1804]), .Z(n2468) );
  XOR U2462 ( .A(n2652), .B(n2653), .Z(n2648) );
  AND U2463 ( .A(n2654), .B(n2655), .Z(n2653) );
  XNOR U2464 ( .A(p_input[1819]), .B(n2652), .Z(n2655) );
  XNOR U2465 ( .A(n2652), .B(n2477), .Z(n2654) );
  IV U2466 ( .A(p_input[1803]), .Z(n2477) );
  XOR U2467 ( .A(n2656), .B(n2657), .Z(n2652) );
  AND U2468 ( .A(n2658), .B(n2659), .Z(n2657) );
  XNOR U2469 ( .A(p_input[1818]), .B(n2656), .Z(n2659) );
  XNOR U2470 ( .A(n2656), .B(n2486), .Z(n2658) );
  IV U2471 ( .A(p_input[1802]), .Z(n2486) );
  XOR U2472 ( .A(n2660), .B(n2661), .Z(n2656) );
  AND U2473 ( .A(n2662), .B(n2663), .Z(n2661) );
  XNOR U2474 ( .A(p_input[1817]), .B(n2660), .Z(n2663) );
  XNOR U2475 ( .A(n2660), .B(n2495), .Z(n2662) );
  IV U2476 ( .A(p_input[1801]), .Z(n2495) );
  XOR U2477 ( .A(n2664), .B(n2665), .Z(n2660) );
  AND U2478 ( .A(n2666), .B(n2667), .Z(n2665) );
  XNOR U2479 ( .A(p_input[1816]), .B(n2664), .Z(n2667) );
  XNOR U2480 ( .A(n2664), .B(n2504), .Z(n2666) );
  IV U2481 ( .A(p_input[1800]), .Z(n2504) );
  XOR U2482 ( .A(n2668), .B(n2669), .Z(n2664) );
  AND U2483 ( .A(n2670), .B(n2671), .Z(n2669) );
  XNOR U2484 ( .A(p_input[1815]), .B(n2668), .Z(n2671) );
  XNOR U2485 ( .A(n2668), .B(n2513), .Z(n2670) );
  IV U2486 ( .A(p_input[1799]), .Z(n2513) );
  XOR U2487 ( .A(n2672), .B(n2673), .Z(n2668) );
  AND U2488 ( .A(n2674), .B(n2675), .Z(n2673) );
  XNOR U2489 ( .A(p_input[1814]), .B(n2672), .Z(n2675) );
  XNOR U2490 ( .A(n2672), .B(n2522), .Z(n2674) );
  IV U2491 ( .A(p_input[1798]), .Z(n2522) );
  XOR U2492 ( .A(n2676), .B(n2677), .Z(n2672) );
  AND U2493 ( .A(n2678), .B(n2679), .Z(n2677) );
  XNOR U2494 ( .A(p_input[1813]), .B(n2676), .Z(n2679) );
  XNOR U2495 ( .A(n2676), .B(n2531), .Z(n2678) );
  IV U2496 ( .A(p_input[1797]), .Z(n2531) );
  XOR U2497 ( .A(n2680), .B(n2681), .Z(n2676) );
  AND U2498 ( .A(n2682), .B(n2683), .Z(n2681) );
  XNOR U2499 ( .A(p_input[1812]), .B(n2680), .Z(n2683) );
  XNOR U2500 ( .A(n2680), .B(n2540), .Z(n2682) );
  IV U2501 ( .A(p_input[1796]), .Z(n2540) );
  XOR U2502 ( .A(n2684), .B(n2685), .Z(n2680) );
  AND U2503 ( .A(n2686), .B(n2687), .Z(n2685) );
  XNOR U2504 ( .A(p_input[1811]), .B(n2684), .Z(n2687) );
  XNOR U2505 ( .A(n2684), .B(n2549), .Z(n2686) );
  IV U2506 ( .A(p_input[1795]), .Z(n2549) );
  XOR U2507 ( .A(n2688), .B(n2689), .Z(n2684) );
  AND U2508 ( .A(n2690), .B(n2691), .Z(n2689) );
  XNOR U2509 ( .A(p_input[1810]), .B(n2688), .Z(n2691) );
  XNOR U2510 ( .A(n2688), .B(n2558), .Z(n2690) );
  IV U2511 ( .A(p_input[1794]), .Z(n2558) );
  XNOR U2512 ( .A(n2692), .B(n2693), .Z(n2688) );
  AND U2513 ( .A(n2694), .B(n2695), .Z(n2693) );
  XOR U2514 ( .A(p_input[1809]), .B(n2692), .Z(n2695) );
  XNOR U2515 ( .A(p_input[1793]), .B(n2692), .Z(n2694) );
  AND U2516 ( .A(p_input[1808]), .B(n2696), .Z(n2692) );
  IV U2517 ( .A(p_input[1792]), .Z(n2696) );
  XOR U2518 ( .A(n2697), .B(n2698), .Z(n924) );
  AND U2519 ( .A(n496), .B(n2699), .Z(n2698) );
  XNOR U2520 ( .A(n2700), .B(n2697), .Z(n2699) );
  XOR U2521 ( .A(n2701), .B(n2702), .Z(n496) );
  AND U2522 ( .A(n2703), .B(n2704), .Z(n2702) );
  XNOR U2523 ( .A(n939), .B(n2701), .Z(n2704) );
  AND U2524 ( .A(n2705), .B(n2706), .Z(n939) );
  XNOR U2525 ( .A(n2701), .B(n936), .Z(n2703) );
  IV U2526 ( .A(n2707), .Z(n936) );
  AND U2527 ( .A(n2708), .B(n2709), .Z(n2707) );
  XOR U2528 ( .A(n2710), .B(n2711), .Z(n2701) );
  AND U2529 ( .A(n2712), .B(n2713), .Z(n2711) );
  XOR U2530 ( .A(n2710), .B(n951), .Z(n2713) );
  XOR U2531 ( .A(n2714), .B(n2715), .Z(n951) );
  AND U2532 ( .A(n414), .B(n2716), .Z(n2715) );
  XOR U2533 ( .A(n2717), .B(n2714), .Z(n2716) );
  XNOR U2534 ( .A(n948), .B(n2710), .Z(n2712) );
  XOR U2535 ( .A(n2718), .B(n2719), .Z(n948) );
  AND U2536 ( .A(n411), .B(n2720), .Z(n2719) );
  XOR U2537 ( .A(n2721), .B(n2718), .Z(n2720) );
  XOR U2538 ( .A(n2722), .B(n2723), .Z(n2710) );
  AND U2539 ( .A(n2724), .B(n2725), .Z(n2723) );
  XOR U2540 ( .A(n2722), .B(n963), .Z(n2725) );
  XOR U2541 ( .A(n2726), .B(n2727), .Z(n963) );
  AND U2542 ( .A(n414), .B(n2728), .Z(n2727) );
  XOR U2543 ( .A(n2729), .B(n2726), .Z(n2728) );
  XNOR U2544 ( .A(n960), .B(n2722), .Z(n2724) );
  XOR U2545 ( .A(n2730), .B(n2731), .Z(n960) );
  AND U2546 ( .A(n411), .B(n2732), .Z(n2731) );
  XOR U2547 ( .A(n2733), .B(n2730), .Z(n2732) );
  XOR U2548 ( .A(n2734), .B(n2735), .Z(n2722) );
  AND U2549 ( .A(n2736), .B(n2737), .Z(n2735) );
  XOR U2550 ( .A(n2734), .B(n975), .Z(n2737) );
  XOR U2551 ( .A(n2738), .B(n2739), .Z(n975) );
  AND U2552 ( .A(n414), .B(n2740), .Z(n2739) );
  XOR U2553 ( .A(n2741), .B(n2738), .Z(n2740) );
  XNOR U2554 ( .A(n972), .B(n2734), .Z(n2736) );
  XOR U2555 ( .A(n2742), .B(n2743), .Z(n972) );
  AND U2556 ( .A(n411), .B(n2744), .Z(n2743) );
  XOR U2557 ( .A(n2745), .B(n2742), .Z(n2744) );
  XOR U2558 ( .A(n2746), .B(n2747), .Z(n2734) );
  AND U2559 ( .A(n2748), .B(n2749), .Z(n2747) );
  XOR U2560 ( .A(n2746), .B(n987), .Z(n2749) );
  XOR U2561 ( .A(n2750), .B(n2751), .Z(n987) );
  AND U2562 ( .A(n414), .B(n2752), .Z(n2751) );
  XOR U2563 ( .A(n2753), .B(n2750), .Z(n2752) );
  XNOR U2564 ( .A(n984), .B(n2746), .Z(n2748) );
  XOR U2565 ( .A(n2754), .B(n2755), .Z(n984) );
  AND U2566 ( .A(n411), .B(n2756), .Z(n2755) );
  XOR U2567 ( .A(n2757), .B(n2754), .Z(n2756) );
  XOR U2568 ( .A(n2758), .B(n2759), .Z(n2746) );
  AND U2569 ( .A(n2760), .B(n2761), .Z(n2759) );
  XOR U2570 ( .A(n2758), .B(n999), .Z(n2761) );
  XOR U2571 ( .A(n2762), .B(n2763), .Z(n999) );
  AND U2572 ( .A(n414), .B(n2764), .Z(n2763) );
  XOR U2573 ( .A(n2765), .B(n2762), .Z(n2764) );
  XNOR U2574 ( .A(n996), .B(n2758), .Z(n2760) );
  XOR U2575 ( .A(n2766), .B(n2767), .Z(n996) );
  AND U2576 ( .A(n411), .B(n2768), .Z(n2767) );
  XOR U2577 ( .A(n2769), .B(n2766), .Z(n2768) );
  XOR U2578 ( .A(n2770), .B(n2771), .Z(n2758) );
  AND U2579 ( .A(n2772), .B(n2773), .Z(n2771) );
  XOR U2580 ( .A(n2770), .B(n1011), .Z(n2773) );
  XOR U2581 ( .A(n2774), .B(n2775), .Z(n1011) );
  AND U2582 ( .A(n414), .B(n2776), .Z(n2775) );
  XOR U2583 ( .A(n2777), .B(n2774), .Z(n2776) );
  XNOR U2584 ( .A(n1008), .B(n2770), .Z(n2772) );
  XOR U2585 ( .A(n2778), .B(n2779), .Z(n1008) );
  AND U2586 ( .A(n411), .B(n2780), .Z(n2779) );
  XOR U2587 ( .A(n2781), .B(n2778), .Z(n2780) );
  XOR U2588 ( .A(n2782), .B(n2783), .Z(n2770) );
  AND U2589 ( .A(n2784), .B(n2785), .Z(n2783) );
  XOR U2590 ( .A(n2782), .B(n1023), .Z(n2785) );
  XOR U2591 ( .A(n2786), .B(n2787), .Z(n1023) );
  AND U2592 ( .A(n414), .B(n2788), .Z(n2787) );
  XOR U2593 ( .A(n2789), .B(n2786), .Z(n2788) );
  XNOR U2594 ( .A(n1020), .B(n2782), .Z(n2784) );
  XOR U2595 ( .A(n2790), .B(n2791), .Z(n1020) );
  AND U2596 ( .A(n411), .B(n2792), .Z(n2791) );
  XOR U2597 ( .A(n2793), .B(n2790), .Z(n2792) );
  XOR U2598 ( .A(n2794), .B(n2795), .Z(n2782) );
  AND U2599 ( .A(n2796), .B(n2797), .Z(n2795) );
  XOR U2600 ( .A(n2794), .B(n1035), .Z(n2797) );
  XOR U2601 ( .A(n2798), .B(n2799), .Z(n1035) );
  AND U2602 ( .A(n414), .B(n2800), .Z(n2799) );
  XOR U2603 ( .A(n2801), .B(n2798), .Z(n2800) );
  XNOR U2604 ( .A(n1032), .B(n2794), .Z(n2796) );
  XOR U2605 ( .A(n2802), .B(n2803), .Z(n1032) );
  AND U2606 ( .A(n411), .B(n2804), .Z(n2803) );
  XOR U2607 ( .A(n2805), .B(n2802), .Z(n2804) );
  XOR U2608 ( .A(n2806), .B(n2807), .Z(n2794) );
  AND U2609 ( .A(n2808), .B(n2809), .Z(n2807) );
  XOR U2610 ( .A(n2806), .B(n1047), .Z(n2809) );
  XOR U2611 ( .A(n2810), .B(n2811), .Z(n1047) );
  AND U2612 ( .A(n414), .B(n2812), .Z(n2811) );
  XOR U2613 ( .A(n2813), .B(n2810), .Z(n2812) );
  XNOR U2614 ( .A(n1044), .B(n2806), .Z(n2808) );
  XOR U2615 ( .A(n2814), .B(n2815), .Z(n1044) );
  AND U2616 ( .A(n411), .B(n2816), .Z(n2815) );
  XOR U2617 ( .A(n2817), .B(n2814), .Z(n2816) );
  XOR U2618 ( .A(n2818), .B(n2819), .Z(n2806) );
  AND U2619 ( .A(n2820), .B(n2821), .Z(n2819) );
  XOR U2620 ( .A(n2818), .B(n1059), .Z(n2821) );
  XOR U2621 ( .A(n2822), .B(n2823), .Z(n1059) );
  AND U2622 ( .A(n414), .B(n2824), .Z(n2823) );
  XOR U2623 ( .A(n2825), .B(n2822), .Z(n2824) );
  XNOR U2624 ( .A(n1056), .B(n2818), .Z(n2820) );
  XOR U2625 ( .A(n2826), .B(n2827), .Z(n1056) );
  AND U2626 ( .A(n411), .B(n2828), .Z(n2827) );
  XOR U2627 ( .A(n2829), .B(n2826), .Z(n2828) );
  XOR U2628 ( .A(n2830), .B(n2831), .Z(n2818) );
  AND U2629 ( .A(n2832), .B(n2833), .Z(n2831) );
  XOR U2630 ( .A(n2830), .B(n1071), .Z(n2833) );
  XOR U2631 ( .A(n2834), .B(n2835), .Z(n1071) );
  AND U2632 ( .A(n414), .B(n2836), .Z(n2835) );
  XOR U2633 ( .A(n2837), .B(n2834), .Z(n2836) );
  XNOR U2634 ( .A(n1068), .B(n2830), .Z(n2832) );
  XOR U2635 ( .A(n2838), .B(n2839), .Z(n1068) );
  AND U2636 ( .A(n411), .B(n2840), .Z(n2839) );
  XOR U2637 ( .A(n2841), .B(n2838), .Z(n2840) );
  XOR U2638 ( .A(n2842), .B(n2843), .Z(n2830) );
  AND U2639 ( .A(n2844), .B(n2845), .Z(n2843) );
  XOR U2640 ( .A(n2842), .B(n1083), .Z(n2845) );
  XOR U2641 ( .A(n2846), .B(n2847), .Z(n1083) );
  AND U2642 ( .A(n414), .B(n2848), .Z(n2847) );
  XOR U2643 ( .A(n2849), .B(n2846), .Z(n2848) );
  XNOR U2644 ( .A(n1080), .B(n2842), .Z(n2844) );
  XOR U2645 ( .A(n2850), .B(n2851), .Z(n1080) );
  AND U2646 ( .A(n411), .B(n2852), .Z(n2851) );
  XOR U2647 ( .A(n2853), .B(n2850), .Z(n2852) );
  XOR U2648 ( .A(n2854), .B(n2855), .Z(n2842) );
  AND U2649 ( .A(n2856), .B(n2857), .Z(n2855) );
  XOR U2650 ( .A(n1095), .B(n2854), .Z(n2857) );
  XOR U2651 ( .A(n2858), .B(n2859), .Z(n1095) );
  AND U2652 ( .A(n414), .B(n2860), .Z(n2859) );
  XOR U2653 ( .A(n2858), .B(n2861), .Z(n2860) );
  XNOR U2654 ( .A(n2854), .B(n1092), .Z(n2856) );
  XOR U2655 ( .A(n2862), .B(n2863), .Z(n1092) );
  AND U2656 ( .A(n411), .B(n2864), .Z(n2863) );
  XOR U2657 ( .A(n2862), .B(n2865), .Z(n2864) );
  XOR U2658 ( .A(n2866), .B(n2867), .Z(n2854) );
  AND U2659 ( .A(n2868), .B(n2869), .Z(n2867) );
  XNOR U2660 ( .A(n2870), .B(n1108), .Z(n2869) );
  XOR U2661 ( .A(n2871), .B(n2872), .Z(n1108) );
  AND U2662 ( .A(n414), .B(n2873), .Z(n2872) );
  XOR U2663 ( .A(n2874), .B(n2871), .Z(n2873) );
  XNOR U2664 ( .A(n1105), .B(n2866), .Z(n2868) );
  XOR U2665 ( .A(n2875), .B(n2876), .Z(n1105) );
  AND U2666 ( .A(n411), .B(n2877), .Z(n2876) );
  XOR U2667 ( .A(n2878), .B(n2875), .Z(n2877) );
  IV U2668 ( .A(n2870), .Z(n2866) );
  AND U2669 ( .A(n2697), .B(n2700), .Z(n2870) );
  XNOR U2670 ( .A(n2879), .B(n2880), .Z(n2700) );
  AND U2671 ( .A(n414), .B(n2881), .Z(n2880) );
  XNOR U2672 ( .A(n2882), .B(n2879), .Z(n2881) );
  XOR U2673 ( .A(n2883), .B(n2884), .Z(n414) );
  AND U2674 ( .A(n2885), .B(n2886), .Z(n2884) );
  XNOR U2675 ( .A(n2705), .B(n2883), .Z(n2886) );
  AND U2676 ( .A(n2887), .B(n2888), .Z(n2705) );
  XOR U2677 ( .A(n2883), .B(n2706), .Z(n2885) );
  AND U2678 ( .A(n2889), .B(n2890), .Z(n2706) );
  XOR U2679 ( .A(n2891), .B(n2892), .Z(n2883) );
  AND U2680 ( .A(n2893), .B(n2894), .Z(n2892) );
  XOR U2681 ( .A(n2891), .B(n2717), .Z(n2894) );
  XOR U2682 ( .A(n2895), .B(n2896), .Z(n2717) );
  AND U2683 ( .A(n238), .B(n2897), .Z(n2896) );
  XOR U2684 ( .A(n2898), .B(n2895), .Z(n2897) );
  XNOR U2685 ( .A(n2714), .B(n2891), .Z(n2893) );
  XOR U2686 ( .A(n2899), .B(n2900), .Z(n2714) );
  AND U2687 ( .A(n236), .B(n2901), .Z(n2900) );
  XOR U2688 ( .A(n2902), .B(n2899), .Z(n2901) );
  XOR U2689 ( .A(n2903), .B(n2904), .Z(n2891) );
  AND U2690 ( .A(n2905), .B(n2906), .Z(n2904) );
  XOR U2691 ( .A(n2903), .B(n2729), .Z(n2906) );
  XOR U2692 ( .A(n2907), .B(n2908), .Z(n2729) );
  AND U2693 ( .A(n238), .B(n2909), .Z(n2908) );
  XOR U2694 ( .A(n2910), .B(n2907), .Z(n2909) );
  XNOR U2695 ( .A(n2726), .B(n2903), .Z(n2905) );
  XOR U2696 ( .A(n2911), .B(n2912), .Z(n2726) );
  AND U2697 ( .A(n236), .B(n2913), .Z(n2912) );
  XOR U2698 ( .A(n2914), .B(n2911), .Z(n2913) );
  XOR U2699 ( .A(n2915), .B(n2916), .Z(n2903) );
  AND U2700 ( .A(n2917), .B(n2918), .Z(n2916) );
  XOR U2701 ( .A(n2915), .B(n2741), .Z(n2918) );
  XOR U2702 ( .A(n2919), .B(n2920), .Z(n2741) );
  AND U2703 ( .A(n238), .B(n2921), .Z(n2920) );
  XOR U2704 ( .A(n2922), .B(n2919), .Z(n2921) );
  XNOR U2705 ( .A(n2738), .B(n2915), .Z(n2917) );
  XOR U2706 ( .A(n2923), .B(n2924), .Z(n2738) );
  AND U2707 ( .A(n236), .B(n2925), .Z(n2924) );
  XOR U2708 ( .A(n2926), .B(n2923), .Z(n2925) );
  XOR U2709 ( .A(n2927), .B(n2928), .Z(n2915) );
  AND U2710 ( .A(n2929), .B(n2930), .Z(n2928) );
  XOR U2711 ( .A(n2927), .B(n2753), .Z(n2930) );
  XOR U2712 ( .A(n2931), .B(n2932), .Z(n2753) );
  AND U2713 ( .A(n238), .B(n2933), .Z(n2932) );
  XOR U2714 ( .A(n2934), .B(n2931), .Z(n2933) );
  XNOR U2715 ( .A(n2750), .B(n2927), .Z(n2929) );
  XOR U2716 ( .A(n2935), .B(n2936), .Z(n2750) );
  AND U2717 ( .A(n236), .B(n2937), .Z(n2936) );
  XOR U2718 ( .A(n2938), .B(n2935), .Z(n2937) );
  XOR U2719 ( .A(n2939), .B(n2940), .Z(n2927) );
  AND U2720 ( .A(n2941), .B(n2942), .Z(n2940) );
  XOR U2721 ( .A(n2939), .B(n2765), .Z(n2942) );
  XOR U2722 ( .A(n2943), .B(n2944), .Z(n2765) );
  AND U2723 ( .A(n238), .B(n2945), .Z(n2944) );
  XOR U2724 ( .A(n2946), .B(n2943), .Z(n2945) );
  XNOR U2725 ( .A(n2762), .B(n2939), .Z(n2941) );
  XOR U2726 ( .A(n2947), .B(n2948), .Z(n2762) );
  AND U2727 ( .A(n236), .B(n2949), .Z(n2948) );
  XOR U2728 ( .A(n2950), .B(n2947), .Z(n2949) );
  XOR U2729 ( .A(n2951), .B(n2952), .Z(n2939) );
  AND U2730 ( .A(n2953), .B(n2954), .Z(n2952) );
  XOR U2731 ( .A(n2951), .B(n2777), .Z(n2954) );
  XOR U2732 ( .A(n2955), .B(n2956), .Z(n2777) );
  AND U2733 ( .A(n238), .B(n2957), .Z(n2956) );
  XOR U2734 ( .A(n2958), .B(n2955), .Z(n2957) );
  XNOR U2735 ( .A(n2774), .B(n2951), .Z(n2953) );
  XOR U2736 ( .A(n2959), .B(n2960), .Z(n2774) );
  AND U2737 ( .A(n236), .B(n2961), .Z(n2960) );
  XOR U2738 ( .A(n2962), .B(n2959), .Z(n2961) );
  XOR U2739 ( .A(n2963), .B(n2964), .Z(n2951) );
  AND U2740 ( .A(n2965), .B(n2966), .Z(n2964) );
  XOR U2741 ( .A(n2963), .B(n2789), .Z(n2966) );
  XOR U2742 ( .A(n2967), .B(n2968), .Z(n2789) );
  AND U2743 ( .A(n238), .B(n2969), .Z(n2968) );
  XOR U2744 ( .A(n2970), .B(n2967), .Z(n2969) );
  XNOR U2745 ( .A(n2786), .B(n2963), .Z(n2965) );
  XOR U2746 ( .A(n2971), .B(n2972), .Z(n2786) );
  AND U2747 ( .A(n236), .B(n2973), .Z(n2972) );
  XOR U2748 ( .A(n2974), .B(n2971), .Z(n2973) );
  XOR U2749 ( .A(n2975), .B(n2976), .Z(n2963) );
  AND U2750 ( .A(n2977), .B(n2978), .Z(n2976) );
  XOR U2751 ( .A(n2975), .B(n2801), .Z(n2978) );
  XOR U2752 ( .A(n2979), .B(n2980), .Z(n2801) );
  AND U2753 ( .A(n238), .B(n2981), .Z(n2980) );
  XOR U2754 ( .A(n2982), .B(n2979), .Z(n2981) );
  XNOR U2755 ( .A(n2798), .B(n2975), .Z(n2977) );
  XOR U2756 ( .A(n2983), .B(n2984), .Z(n2798) );
  AND U2757 ( .A(n236), .B(n2985), .Z(n2984) );
  XOR U2758 ( .A(n2986), .B(n2983), .Z(n2985) );
  XOR U2759 ( .A(n2987), .B(n2988), .Z(n2975) );
  AND U2760 ( .A(n2989), .B(n2990), .Z(n2988) );
  XOR U2761 ( .A(n2987), .B(n2813), .Z(n2990) );
  XOR U2762 ( .A(n2991), .B(n2992), .Z(n2813) );
  AND U2763 ( .A(n238), .B(n2993), .Z(n2992) );
  XOR U2764 ( .A(n2994), .B(n2991), .Z(n2993) );
  XNOR U2765 ( .A(n2810), .B(n2987), .Z(n2989) );
  XOR U2766 ( .A(n2995), .B(n2996), .Z(n2810) );
  AND U2767 ( .A(n236), .B(n2997), .Z(n2996) );
  XOR U2768 ( .A(n2998), .B(n2995), .Z(n2997) );
  XOR U2769 ( .A(n2999), .B(n3000), .Z(n2987) );
  AND U2770 ( .A(n3001), .B(n3002), .Z(n3000) );
  XOR U2771 ( .A(n2999), .B(n2825), .Z(n3002) );
  XOR U2772 ( .A(n3003), .B(n3004), .Z(n2825) );
  AND U2773 ( .A(n238), .B(n3005), .Z(n3004) );
  XOR U2774 ( .A(n3006), .B(n3003), .Z(n3005) );
  XNOR U2775 ( .A(n2822), .B(n2999), .Z(n3001) );
  XOR U2776 ( .A(n3007), .B(n3008), .Z(n2822) );
  AND U2777 ( .A(n236), .B(n3009), .Z(n3008) );
  XOR U2778 ( .A(n3010), .B(n3007), .Z(n3009) );
  XOR U2779 ( .A(n3011), .B(n3012), .Z(n2999) );
  AND U2780 ( .A(n3013), .B(n3014), .Z(n3012) );
  XOR U2781 ( .A(n3011), .B(n2837), .Z(n3014) );
  XOR U2782 ( .A(n3015), .B(n3016), .Z(n2837) );
  AND U2783 ( .A(n238), .B(n3017), .Z(n3016) );
  XOR U2784 ( .A(n3018), .B(n3015), .Z(n3017) );
  XNOR U2785 ( .A(n2834), .B(n3011), .Z(n3013) );
  XOR U2786 ( .A(n3019), .B(n3020), .Z(n2834) );
  AND U2787 ( .A(n236), .B(n3021), .Z(n3020) );
  XOR U2788 ( .A(n3022), .B(n3019), .Z(n3021) );
  XOR U2789 ( .A(n3023), .B(n3024), .Z(n3011) );
  AND U2790 ( .A(n3025), .B(n3026), .Z(n3024) );
  XOR U2791 ( .A(n3023), .B(n2849), .Z(n3026) );
  XOR U2792 ( .A(n3027), .B(n3028), .Z(n2849) );
  AND U2793 ( .A(n238), .B(n3029), .Z(n3028) );
  XOR U2794 ( .A(n3030), .B(n3027), .Z(n3029) );
  XNOR U2795 ( .A(n2846), .B(n3023), .Z(n3025) );
  XOR U2796 ( .A(n3031), .B(n3032), .Z(n2846) );
  AND U2797 ( .A(n236), .B(n3033), .Z(n3032) );
  XOR U2798 ( .A(n3034), .B(n3031), .Z(n3033) );
  XOR U2799 ( .A(n3035), .B(n3036), .Z(n3023) );
  AND U2800 ( .A(n3037), .B(n3038), .Z(n3036) );
  XOR U2801 ( .A(n2861), .B(n3035), .Z(n3038) );
  XOR U2802 ( .A(n3039), .B(n3040), .Z(n2861) );
  AND U2803 ( .A(n238), .B(n3041), .Z(n3040) );
  XOR U2804 ( .A(n3039), .B(n3042), .Z(n3041) );
  XNOR U2805 ( .A(n3035), .B(n2858), .Z(n3037) );
  XOR U2806 ( .A(n3043), .B(n3044), .Z(n2858) );
  AND U2807 ( .A(n236), .B(n3045), .Z(n3044) );
  XOR U2808 ( .A(n3043), .B(n3046), .Z(n3045) );
  XOR U2809 ( .A(n3047), .B(n3048), .Z(n3035) );
  AND U2810 ( .A(n3049), .B(n3050), .Z(n3048) );
  XNOR U2811 ( .A(n3051), .B(n2874), .Z(n3050) );
  XOR U2812 ( .A(n3052), .B(n3053), .Z(n2874) );
  AND U2813 ( .A(n238), .B(n3054), .Z(n3053) );
  XOR U2814 ( .A(n3055), .B(n3052), .Z(n3054) );
  XNOR U2815 ( .A(n2871), .B(n3047), .Z(n3049) );
  XOR U2816 ( .A(n3056), .B(n3057), .Z(n2871) );
  AND U2817 ( .A(n236), .B(n3058), .Z(n3057) );
  XOR U2818 ( .A(n3059), .B(n3056), .Z(n3058) );
  IV U2819 ( .A(n3051), .Z(n3047) );
  AND U2820 ( .A(n2879), .B(n2882), .Z(n3051) );
  XNOR U2821 ( .A(n3060), .B(n3061), .Z(n2882) );
  AND U2822 ( .A(n238), .B(n3062), .Z(n3061) );
  XNOR U2823 ( .A(n3063), .B(n3060), .Z(n3062) );
  XOR U2824 ( .A(n3064), .B(n3065), .Z(n238) );
  AND U2825 ( .A(n3066), .B(n3067), .Z(n3065) );
  XNOR U2826 ( .A(n2887), .B(n3064), .Z(n3067) );
  AND U2827 ( .A(p_input[1791]), .B(p_input[1775]), .Z(n2887) );
  XOR U2828 ( .A(n3064), .B(n2888), .Z(n3066) );
  AND U2829 ( .A(p_input[1759]), .B(p_input[1743]), .Z(n2888) );
  XOR U2830 ( .A(n3068), .B(n3069), .Z(n3064) );
  AND U2831 ( .A(n3070), .B(n3071), .Z(n3069) );
  XOR U2832 ( .A(n3068), .B(n2898), .Z(n3071) );
  XNOR U2833 ( .A(p_input[1774]), .B(n3072), .Z(n2898) );
  AND U2834 ( .A(n130), .B(n3073), .Z(n3072) );
  XOR U2835 ( .A(p_input[1790]), .B(p_input[1774]), .Z(n3073) );
  XNOR U2836 ( .A(n2895), .B(n3068), .Z(n3070) );
  XOR U2837 ( .A(n3074), .B(n3075), .Z(n2895) );
  AND U2838 ( .A(n128), .B(n3076), .Z(n3075) );
  XOR U2839 ( .A(p_input[1758]), .B(p_input[1742]), .Z(n3076) );
  XOR U2840 ( .A(n3077), .B(n3078), .Z(n3068) );
  AND U2841 ( .A(n3079), .B(n3080), .Z(n3078) );
  XOR U2842 ( .A(n3077), .B(n2910), .Z(n3080) );
  XNOR U2843 ( .A(p_input[1773]), .B(n3081), .Z(n2910) );
  AND U2844 ( .A(n130), .B(n3082), .Z(n3081) );
  XOR U2845 ( .A(p_input[1789]), .B(p_input[1773]), .Z(n3082) );
  XNOR U2846 ( .A(n2907), .B(n3077), .Z(n3079) );
  XOR U2847 ( .A(n3083), .B(n3084), .Z(n2907) );
  AND U2848 ( .A(n128), .B(n3085), .Z(n3084) );
  XOR U2849 ( .A(p_input[1757]), .B(p_input[1741]), .Z(n3085) );
  XOR U2850 ( .A(n3086), .B(n3087), .Z(n3077) );
  AND U2851 ( .A(n3088), .B(n3089), .Z(n3087) );
  XOR U2852 ( .A(n3086), .B(n2922), .Z(n3089) );
  XNOR U2853 ( .A(p_input[1772]), .B(n3090), .Z(n2922) );
  AND U2854 ( .A(n130), .B(n3091), .Z(n3090) );
  XOR U2855 ( .A(p_input[1788]), .B(p_input[1772]), .Z(n3091) );
  XNOR U2856 ( .A(n2919), .B(n3086), .Z(n3088) );
  XOR U2857 ( .A(n3092), .B(n3093), .Z(n2919) );
  AND U2858 ( .A(n128), .B(n3094), .Z(n3093) );
  XOR U2859 ( .A(p_input[1756]), .B(p_input[1740]), .Z(n3094) );
  XOR U2860 ( .A(n3095), .B(n3096), .Z(n3086) );
  AND U2861 ( .A(n3097), .B(n3098), .Z(n3096) );
  XOR U2862 ( .A(n3095), .B(n2934), .Z(n3098) );
  XNOR U2863 ( .A(p_input[1771]), .B(n3099), .Z(n2934) );
  AND U2864 ( .A(n130), .B(n3100), .Z(n3099) );
  XOR U2865 ( .A(p_input[1787]), .B(p_input[1771]), .Z(n3100) );
  XNOR U2866 ( .A(n2931), .B(n3095), .Z(n3097) );
  XOR U2867 ( .A(n3101), .B(n3102), .Z(n2931) );
  AND U2868 ( .A(n128), .B(n3103), .Z(n3102) );
  XOR U2869 ( .A(p_input[1755]), .B(p_input[1739]), .Z(n3103) );
  XOR U2870 ( .A(n3104), .B(n3105), .Z(n3095) );
  AND U2871 ( .A(n3106), .B(n3107), .Z(n3105) );
  XOR U2872 ( .A(n3104), .B(n2946), .Z(n3107) );
  XNOR U2873 ( .A(p_input[1770]), .B(n3108), .Z(n2946) );
  AND U2874 ( .A(n130), .B(n3109), .Z(n3108) );
  XOR U2875 ( .A(p_input[1786]), .B(p_input[1770]), .Z(n3109) );
  XNOR U2876 ( .A(n2943), .B(n3104), .Z(n3106) );
  XOR U2877 ( .A(n3110), .B(n3111), .Z(n2943) );
  AND U2878 ( .A(n128), .B(n3112), .Z(n3111) );
  XOR U2879 ( .A(p_input[1754]), .B(p_input[1738]), .Z(n3112) );
  XOR U2880 ( .A(n3113), .B(n3114), .Z(n3104) );
  AND U2881 ( .A(n3115), .B(n3116), .Z(n3114) );
  XOR U2882 ( .A(n3113), .B(n2958), .Z(n3116) );
  XNOR U2883 ( .A(p_input[1769]), .B(n3117), .Z(n2958) );
  AND U2884 ( .A(n130), .B(n3118), .Z(n3117) );
  XOR U2885 ( .A(p_input[1785]), .B(p_input[1769]), .Z(n3118) );
  XNOR U2886 ( .A(n2955), .B(n3113), .Z(n3115) );
  XOR U2887 ( .A(n3119), .B(n3120), .Z(n2955) );
  AND U2888 ( .A(n128), .B(n3121), .Z(n3120) );
  XOR U2889 ( .A(p_input[1753]), .B(p_input[1737]), .Z(n3121) );
  XOR U2890 ( .A(n3122), .B(n3123), .Z(n3113) );
  AND U2891 ( .A(n3124), .B(n3125), .Z(n3123) );
  XOR U2892 ( .A(n3122), .B(n2970), .Z(n3125) );
  XNOR U2893 ( .A(p_input[1768]), .B(n3126), .Z(n2970) );
  AND U2894 ( .A(n130), .B(n3127), .Z(n3126) );
  XOR U2895 ( .A(p_input[1784]), .B(p_input[1768]), .Z(n3127) );
  XNOR U2896 ( .A(n2967), .B(n3122), .Z(n3124) );
  XOR U2897 ( .A(n3128), .B(n3129), .Z(n2967) );
  AND U2898 ( .A(n128), .B(n3130), .Z(n3129) );
  XOR U2899 ( .A(p_input[1752]), .B(p_input[1736]), .Z(n3130) );
  XOR U2900 ( .A(n3131), .B(n3132), .Z(n3122) );
  AND U2901 ( .A(n3133), .B(n3134), .Z(n3132) );
  XOR U2902 ( .A(n3131), .B(n2982), .Z(n3134) );
  XNOR U2903 ( .A(p_input[1767]), .B(n3135), .Z(n2982) );
  AND U2904 ( .A(n130), .B(n3136), .Z(n3135) );
  XOR U2905 ( .A(p_input[1783]), .B(p_input[1767]), .Z(n3136) );
  XNOR U2906 ( .A(n2979), .B(n3131), .Z(n3133) );
  XOR U2907 ( .A(n3137), .B(n3138), .Z(n2979) );
  AND U2908 ( .A(n128), .B(n3139), .Z(n3138) );
  XOR U2909 ( .A(p_input[1751]), .B(p_input[1735]), .Z(n3139) );
  XOR U2910 ( .A(n3140), .B(n3141), .Z(n3131) );
  AND U2911 ( .A(n3142), .B(n3143), .Z(n3141) );
  XOR U2912 ( .A(n3140), .B(n2994), .Z(n3143) );
  XNOR U2913 ( .A(p_input[1766]), .B(n3144), .Z(n2994) );
  AND U2914 ( .A(n130), .B(n3145), .Z(n3144) );
  XOR U2915 ( .A(p_input[1782]), .B(p_input[1766]), .Z(n3145) );
  XNOR U2916 ( .A(n2991), .B(n3140), .Z(n3142) );
  XOR U2917 ( .A(n3146), .B(n3147), .Z(n2991) );
  AND U2918 ( .A(n128), .B(n3148), .Z(n3147) );
  XOR U2919 ( .A(p_input[1750]), .B(p_input[1734]), .Z(n3148) );
  XOR U2920 ( .A(n3149), .B(n3150), .Z(n3140) );
  AND U2921 ( .A(n3151), .B(n3152), .Z(n3150) );
  XOR U2922 ( .A(n3149), .B(n3006), .Z(n3152) );
  XNOR U2923 ( .A(p_input[1765]), .B(n3153), .Z(n3006) );
  AND U2924 ( .A(n130), .B(n3154), .Z(n3153) );
  XOR U2925 ( .A(p_input[1781]), .B(p_input[1765]), .Z(n3154) );
  XNOR U2926 ( .A(n3003), .B(n3149), .Z(n3151) );
  XOR U2927 ( .A(n3155), .B(n3156), .Z(n3003) );
  AND U2928 ( .A(n128), .B(n3157), .Z(n3156) );
  XOR U2929 ( .A(p_input[1749]), .B(p_input[1733]), .Z(n3157) );
  XOR U2930 ( .A(n3158), .B(n3159), .Z(n3149) );
  AND U2931 ( .A(n3160), .B(n3161), .Z(n3159) );
  XOR U2932 ( .A(n3158), .B(n3018), .Z(n3161) );
  XNOR U2933 ( .A(p_input[1764]), .B(n3162), .Z(n3018) );
  AND U2934 ( .A(n130), .B(n3163), .Z(n3162) );
  XOR U2935 ( .A(p_input[1780]), .B(p_input[1764]), .Z(n3163) );
  XNOR U2936 ( .A(n3015), .B(n3158), .Z(n3160) );
  XOR U2937 ( .A(n3164), .B(n3165), .Z(n3015) );
  AND U2938 ( .A(n128), .B(n3166), .Z(n3165) );
  XOR U2939 ( .A(p_input[1748]), .B(p_input[1732]), .Z(n3166) );
  XOR U2940 ( .A(n3167), .B(n3168), .Z(n3158) );
  AND U2941 ( .A(n3169), .B(n3170), .Z(n3168) );
  XOR U2942 ( .A(n3167), .B(n3030), .Z(n3170) );
  XNOR U2943 ( .A(p_input[1763]), .B(n3171), .Z(n3030) );
  AND U2944 ( .A(n130), .B(n3172), .Z(n3171) );
  XOR U2945 ( .A(p_input[1779]), .B(p_input[1763]), .Z(n3172) );
  XNOR U2946 ( .A(n3027), .B(n3167), .Z(n3169) );
  XOR U2947 ( .A(n3173), .B(n3174), .Z(n3027) );
  AND U2948 ( .A(n128), .B(n3175), .Z(n3174) );
  XOR U2949 ( .A(p_input[1747]), .B(p_input[1731]), .Z(n3175) );
  XOR U2950 ( .A(n3176), .B(n3177), .Z(n3167) );
  AND U2951 ( .A(n3178), .B(n3179), .Z(n3177) );
  XOR U2952 ( .A(n3042), .B(n3176), .Z(n3179) );
  XNOR U2953 ( .A(p_input[1762]), .B(n3180), .Z(n3042) );
  AND U2954 ( .A(n130), .B(n3181), .Z(n3180) );
  XOR U2955 ( .A(p_input[1778]), .B(p_input[1762]), .Z(n3181) );
  XNOR U2956 ( .A(n3176), .B(n3039), .Z(n3178) );
  XOR U2957 ( .A(n3182), .B(n3183), .Z(n3039) );
  AND U2958 ( .A(n128), .B(n3184), .Z(n3183) );
  XOR U2959 ( .A(p_input[1746]), .B(p_input[1730]), .Z(n3184) );
  XOR U2960 ( .A(n3185), .B(n3186), .Z(n3176) );
  AND U2961 ( .A(n3187), .B(n3188), .Z(n3186) );
  XNOR U2962 ( .A(n3189), .B(n3055), .Z(n3188) );
  XNOR U2963 ( .A(p_input[1761]), .B(n3190), .Z(n3055) );
  AND U2964 ( .A(n130), .B(n3191), .Z(n3190) );
  XNOR U2965 ( .A(p_input[1777]), .B(n3192), .Z(n3191) );
  IV U2966 ( .A(p_input[1761]), .Z(n3192) );
  XNOR U2967 ( .A(n3052), .B(n3185), .Z(n3187) );
  XNOR U2968 ( .A(p_input[1729]), .B(n3193), .Z(n3052) );
  AND U2969 ( .A(n128), .B(n3194), .Z(n3193) );
  XOR U2970 ( .A(p_input[1745]), .B(p_input[1729]), .Z(n3194) );
  IV U2971 ( .A(n3189), .Z(n3185) );
  AND U2972 ( .A(n3060), .B(n3063), .Z(n3189) );
  XOR U2973 ( .A(p_input[1760]), .B(n3195), .Z(n3063) );
  AND U2974 ( .A(n130), .B(n3196), .Z(n3195) );
  XOR U2975 ( .A(p_input[1776]), .B(p_input[1760]), .Z(n3196) );
  XOR U2976 ( .A(n3197), .B(n3198), .Z(n130) );
  AND U2977 ( .A(n3199), .B(n3200), .Z(n3198) );
  XNOR U2978 ( .A(p_input[1791]), .B(n3197), .Z(n3200) );
  XOR U2979 ( .A(n3197), .B(p_input[1775]), .Z(n3199) );
  XOR U2980 ( .A(n3201), .B(n3202), .Z(n3197) );
  AND U2981 ( .A(n3203), .B(n3204), .Z(n3202) );
  XNOR U2982 ( .A(p_input[1790]), .B(n3201), .Z(n3204) );
  XOR U2983 ( .A(n3201), .B(p_input[1774]), .Z(n3203) );
  XOR U2984 ( .A(n3205), .B(n3206), .Z(n3201) );
  AND U2985 ( .A(n3207), .B(n3208), .Z(n3206) );
  XNOR U2986 ( .A(p_input[1789]), .B(n3205), .Z(n3208) );
  XOR U2987 ( .A(n3205), .B(p_input[1773]), .Z(n3207) );
  XOR U2988 ( .A(n3209), .B(n3210), .Z(n3205) );
  AND U2989 ( .A(n3211), .B(n3212), .Z(n3210) );
  XNOR U2990 ( .A(p_input[1788]), .B(n3209), .Z(n3212) );
  XOR U2991 ( .A(n3209), .B(p_input[1772]), .Z(n3211) );
  XOR U2992 ( .A(n3213), .B(n3214), .Z(n3209) );
  AND U2993 ( .A(n3215), .B(n3216), .Z(n3214) );
  XNOR U2994 ( .A(p_input[1787]), .B(n3213), .Z(n3216) );
  XOR U2995 ( .A(n3213), .B(p_input[1771]), .Z(n3215) );
  XOR U2996 ( .A(n3217), .B(n3218), .Z(n3213) );
  AND U2997 ( .A(n3219), .B(n3220), .Z(n3218) );
  XNOR U2998 ( .A(p_input[1786]), .B(n3217), .Z(n3220) );
  XOR U2999 ( .A(n3217), .B(p_input[1770]), .Z(n3219) );
  XOR U3000 ( .A(n3221), .B(n3222), .Z(n3217) );
  AND U3001 ( .A(n3223), .B(n3224), .Z(n3222) );
  XNOR U3002 ( .A(p_input[1785]), .B(n3221), .Z(n3224) );
  XOR U3003 ( .A(n3221), .B(p_input[1769]), .Z(n3223) );
  XOR U3004 ( .A(n3225), .B(n3226), .Z(n3221) );
  AND U3005 ( .A(n3227), .B(n3228), .Z(n3226) );
  XNOR U3006 ( .A(p_input[1784]), .B(n3225), .Z(n3228) );
  XOR U3007 ( .A(n3225), .B(p_input[1768]), .Z(n3227) );
  XOR U3008 ( .A(n3229), .B(n3230), .Z(n3225) );
  AND U3009 ( .A(n3231), .B(n3232), .Z(n3230) );
  XNOR U3010 ( .A(p_input[1783]), .B(n3229), .Z(n3232) );
  XOR U3011 ( .A(n3229), .B(p_input[1767]), .Z(n3231) );
  XOR U3012 ( .A(n3233), .B(n3234), .Z(n3229) );
  AND U3013 ( .A(n3235), .B(n3236), .Z(n3234) );
  XNOR U3014 ( .A(p_input[1782]), .B(n3233), .Z(n3236) );
  XOR U3015 ( .A(n3233), .B(p_input[1766]), .Z(n3235) );
  XOR U3016 ( .A(n3237), .B(n3238), .Z(n3233) );
  AND U3017 ( .A(n3239), .B(n3240), .Z(n3238) );
  XNOR U3018 ( .A(p_input[1781]), .B(n3237), .Z(n3240) );
  XOR U3019 ( .A(n3237), .B(p_input[1765]), .Z(n3239) );
  XOR U3020 ( .A(n3241), .B(n3242), .Z(n3237) );
  AND U3021 ( .A(n3243), .B(n3244), .Z(n3242) );
  XNOR U3022 ( .A(p_input[1780]), .B(n3241), .Z(n3244) );
  XOR U3023 ( .A(n3241), .B(p_input[1764]), .Z(n3243) );
  XOR U3024 ( .A(n3245), .B(n3246), .Z(n3241) );
  AND U3025 ( .A(n3247), .B(n3248), .Z(n3246) );
  XNOR U3026 ( .A(p_input[1779]), .B(n3245), .Z(n3248) );
  XOR U3027 ( .A(n3245), .B(p_input[1763]), .Z(n3247) );
  XOR U3028 ( .A(n3249), .B(n3250), .Z(n3245) );
  AND U3029 ( .A(n3251), .B(n3252), .Z(n3250) );
  XNOR U3030 ( .A(p_input[1778]), .B(n3249), .Z(n3252) );
  XOR U3031 ( .A(n3249), .B(p_input[1762]), .Z(n3251) );
  XNOR U3032 ( .A(n3253), .B(n3254), .Z(n3249) );
  AND U3033 ( .A(n3255), .B(n3256), .Z(n3254) );
  XOR U3034 ( .A(p_input[1777]), .B(n3253), .Z(n3256) );
  XNOR U3035 ( .A(p_input[1761]), .B(n3253), .Z(n3255) );
  AND U3036 ( .A(p_input[1776]), .B(n3257), .Z(n3253) );
  IV U3037 ( .A(p_input[1760]), .Z(n3257) );
  XNOR U3038 ( .A(p_input[1728]), .B(n3258), .Z(n3060) );
  AND U3039 ( .A(n128), .B(n3259), .Z(n3258) );
  XOR U3040 ( .A(p_input[1744]), .B(p_input[1728]), .Z(n3259) );
  XOR U3041 ( .A(n3260), .B(n3261), .Z(n128) );
  AND U3042 ( .A(n3262), .B(n3263), .Z(n3261) );
  XNOR U3043 ( .A(p_input[1759]), .B(n3260), .Z(n3263) );
  XOR U3044 ( .A(n3260), .B(p_input[1743]), .Z(n3262) );
  XOR U3045 ( .A(n3264), .B(n3265), .Z(n3260) );
  AND U3046 ( .A(n3266), .B(n3267), .Z(n3265) );
  XNOR U3047 ( .A(p_input[1758]), .B(n3264), .Z(n3267) );
  XNOR U3048 ( .A(n3264), .B(n3074), .Z(n3266) );
  IV U3049 ( .A(p_input[1742]), .Z(n3074) );
  XOR U3050 ( .A(n3268), .B(n3269), .Z(n3264) );
  AND U3051 ( .A(n3270), .B(n3271), .Z(n3269) );
  XNOR U3052 ( .A(p_input[1757]), .B(n3268), .Z(n3271) );
  XNOR U3053 ( .A(n3268), .B(n3083), .Z(n3270) );
  IV U3054 ( .A(p_input[1741]), .Z(n3083) );
  XOR U3055 ( .A(n3272), .B(n3273), .Z(n3268) );
  AND U3056 ( .A(n3274), .B(n3275), .Z(n3273) );
  XNOR U3057 ( .A(p_input[1756]), .B(n3272), .Z(n3275) );
  XNOR U3058 ( .A(n3272), .B(n3092), .Z(n3274) );
  IV U3059 ( .A(p_input[1740]), .Z(n3092) );
  XOR U3060 ( .A(n3276), .B(n3277), .Z(n3272) );
  AND U3061 ( .A(n3278), .B(n3279), .Z(n3277) );
  XNOR U3062 ( .A(p_input[1755]), .B(n3276), .Z(n3279) );
  XNOR U3063 ( .A(n3276), .B(n3101), .Z(n3278) );
  IV U3064 ( .A(p_input[1739]), .Z(n3101) );
  XOR U3065 ( .A(n3280), .B(n3281), .Z(n3276) );
  AND U3066 ( .A(n3282), .B(n3283), .Z(n3281) );
  XNOR U3067 ( .A(p_input[1754]), .B(n3280), .Z(n3283) );
  XNOR U3068 ( .A(n3280), .B(n3110), .Z(n3282) );
  IV U3069 ( .A(p_input[1738]), .Z(n3110) );
  XOR U3070 ( .A(n3284), .B(n3285), .Z(n3280) );
  AND U3071 ( .A(n3286), .B(n3287), .Z(n3285) );
  XNOR U3072 ( .A(p_input[1753]), .B(n3284), .Z(n3287) );
  XNOR U3073 ( .A(n3284), .B(n3119), .Z(n3286) );
  IV U3074 ( .A(p_input[1737]), .Z(n3119) );
  XOR U3075 ( .A(n3288), .B(n3289), .Z(n3284) );
  AND U3076 ( .A(n3290), .B(n3291), .Z(n3289) );
  XNOR U3077 ( .A(p_input[1752]), .B(n3288), .Z(n3291) );
  XNOR U3078 ( .A(n3288), .B(n3128), .Z(n3290) );
  IV U3079 ( .A(p_input[1736]), .Z(n3128) );
  XOR U3080 ( .A(n3292), .B(n3293), .Z(n3288) );
  AND U3081 ( .A(n3294), .B(n3295), .Z(n3293) );
  XNOR U3082 ( .A(p_input[1751]), .B(n3292), .Z(n3295) );
  XNOR U3083 ( .A(n3292), .B(n3137), .Z(n3294) );
  IV U3084 ( .A(p_input[1735]), .Z(n3137) );
  XOR U3085 ( .A(n3296), .B(n3297), .Z(n3292) );
  AND U3086 ( .A(n3298), .B(n3299), .Z(n3297) );
  XNOR U3087 ( .A(p_input[1750]), .B(n3296), .Z(n3299) );
  XNOR U3088 ( .A(n3296), .B(n3146), .Z(n3298) );
  IV U3089 ( .A(p_input[1734]), .Z(n3146) );
  XOR U3090 ( .A(n3300), .B(n3301), .Z(n3296) );
  AND U3091 ( .A(n3302), .B(n3303), .Z(n3301) );
  XNOR U3092 ( .A(p_input[1749]), .B(n3300), .Z(n3303) );
  XNOR U3093 ( .A(n3300), .B(n3155), .Z(n3302) );
  IV U3094 ( .A(p_input[1733]), .Z(n3155) );
  XOR U3095 ( .A(n3304), .B(n3305), .Z(n3300) );
  AND U3096 ( .A(n3306), .B(n3307), .Z(n3305) );
  XNOR U3097 ( .A(p_input[1748]), .B(n3304), .Z(n3307) );
  XNOR U3098 ( .A(n3304), .B(n3164), .Z(n3306) );
  IV U3099 ( .A(p_input[1732]), .Z(n3164) );
  XOR U3100 ( .A(n3308), .B(n3309), .Z(n3304) );
  AND U3101 ( .A(n3310), .B(n3311), .Z(n3309) );
  XNOR U3102 ( .A(p_input[1747]), .B(n3308), .Z(n3311) );
  XNOR U3103 ( .A(n3308), .B(n3173), .Z(n3310) );
  IV U3104 ( .A(p_input[1731]), .Z(n3173) );
  XOR U3105 ( .A(n3312), .B(n3313), .Z(n3308) );
  AND U3106 ( .A(n3314), .B(n3315), .Z(n3313) );
  XNOR U3107 ( .A(p_input[1746]), .B(n3312), .Z(n3315) );
  XNOR U3108 ( .A(n3312), .B(n3182), .Z(n3314) );
  IV U3109 ( .A(p_input[1730]), .Z(n3182) );
  XNOR U3110 ( .A(n3316), .B(n3317), .Z(n3312) );
  AND U3111 ( .A(n3318), .B(n3319), .Z(n3317) );
  XOR U3112 ( .A(p_input[1745]), .B(n3316), .Z(n3319) );
  XNOR U3113 ( .A(p_input[1729]), .B(n3316), .Z(n3318) );
  AND U3114 ( .A(p_input[1744]), .B(n3320), .Z(n3316) );
  IV U3115 ( .A(p_input[1728]), .Z(n3320) );
  XOR U3116 ( .A(n3321), .B(n3322), .Z(n2879) );
  AND U3117 ( .A(n236), .B(n3323), .Z(n3322) );
  XNOR U3118 ( .A(n3324), .B(n3321), .Z(n3323) );
  XOR U3119 ( .A(n3325), .B(n3326), .Z(n236) );
  AND U3120 ( .A(n3327), .B(n3328), .Z(n3326) );
  XNOR U3121 ( .A(n2889), .B(n3325), .Z(n3328) );
  AND U3122 ( .A(p_input[1727]), .B(p_input[1711]), .Z(n2889) );
  XOR U3123 ( .A(n3325), .B(n2890), .Z(n3327) );
  AND U3124 ( .A(p_input[1695]), .B(p_input[1679]), .Z(n2890) );
  XOR U3125 ( .A(n3329), .B(n3330), .Z(n3325) );
  AND U3126 ( .A(n3331), .B(n3332), .Z(n3330) );
  XOR U3127 ( .A(n3329), .B(n2902), .Z(n3332) );
  XNOR U3128 ( .A(p_input[1710]), .B(n3333), .Z(n2902) );
  AND U3129 ( .A(n134), .B(n3334), .Z(n3333) );
  XOR U3130 ( .A(p_input[1726]), .B(p_input[1710]), .Z(n3334) );
  XNOR U3131 ( .A(n2899), .B(n3329), .Z(n3331) );
  XOR U3132 ( .A(n3335), .B(n3336), .Z(n2899) );
  AND U3133 ( .A(n131), .B(n3337), .Z(n3336) );
  XOR U3134 ( .A(p_input[1694]), .B(p_input[1678]), .Z(n3337) );
  XOR U3135 ( .A(n3338), .B(n3339), .Z(n3329) );
  AND U3136 ( .A(n3340), .B(n3341), .Z(n3339) );
  XOR U3137 ( .A(n3338), .B(n2914), .Z(n3341) );
  XNOR U3138 ( .A(p_input[1709]), .B(n3342), .Z(n2914) );
  AND U3139 ( .A(n134), .B(n3343), .Z(n3342) );
  XOR U3140 ( .A(p_input[1725]), .B(p_input[1709]), .Z(n3343) );
  XNOR U3141 ( .A(n2911), .B(n3338), .Z(n3340) );
  XOR U3142 ( .A(n3344), .B(n3345), .Z(n2911) );
  AND U3143 ( .A(n131), .B(n3346), .Z(n3345) );
  XOR U3144 ( .A(p_input[1693]), .B(p_input[1677]), .Z(n3346) );
  XOR U3145 ( .A(n3347), .B(n3348), .Z(n3338) );
  AND U3146 ( .A(n3349), .B(n3350), .Z(n3348) );
  XOR U3147 ( .A(n3347), .B(n2926), .Z(n3350) );
  XNOR U3148 ( .A(p_input[1708]), .B(n3351), .Z(n2926) );
  AND U3149 ( .A(n134), .B(n3352), .Z(n3351) );
  XOR U3150 ( .A(p_input[1724]), .B(p_input[1708]), .Z(n3352) );
  XNOR U3151 ( .A(n2923), .B(n3347), .Z(n3349) );
  XOR U3152 ( .A(n3353), .B(n3354), .Z(n2923) );
  AND U3153 ( .A(n131), .B(n3355), .Z(n3354) );
  XOR U3154 ( .A(p_input[1692]), .B(p_input[1676]), .Z(n3355) );
  XOR U3155 ( .A(n3356), .B(n3357), .Z(n3347) );
  AND U3156 ( .A(n3358), .B(n3359), .Z(n3357) );
  XOR U3157 ( .A(n3356), .B(n2938), .Z(n3359) );
  XNOR U3158 ( .A(p_input[1707]), .B(n3360), .Z(n2938) );
  AND U3159 ( .A(n134), .B(n3361), .Z(n3360) );
  XOR U3160 ( .A(p_input[1723]), .B(p_input[1707]), .Z(n3361) );
  XNOR U3161 ( .A(n2935), .B(n3356), .Z(n3358) );
  XOR U3162 ( .A(n3362), .B(n3363), .Z(n2935) );
  AND U3163 ( .A(n131), .B(n3364), .Z(n3363) );
  XOR U3164 ( .A(p_input[1691]), .B(p_input[1675]), .Z(n3364) );
  XOR U3165 ( .A(n3365), .B(n3366), .Z(n3356) );
  AND U3166 ( .A(n3367), .B(n3368), .Z(n3366) );
  XOR U3167 ( .A(n3365), .B(n2950), .Z(n3368) );
  XNOR U3168 ( .A(p_input[1706]), .B(n3369), .Z(n2950) );
  AND U3169 ( .A(n134), .B(n3370), .Z(n3369) );
  XOR U3170 ( .A(p_input[1722]), .B(p_input[1706]), .Z(n3370) );
  XNOR U3171 ( .A(n2947), .B(n3365), .Z(n3367) );
  XOR U3172 ( .A(n3371), .B(n3372), .Z(n2947) );
  AND U3173 ( .A(n131), .B(n3373), .Z(n3372) );
  XOR U3174 ( .A(p_input[1690]), .B(p_input[1674]), .Z(n3373) );
  XOR U3175 ( .A(n3374), .B(n3375), .Z(n3365) );
  AND U3176 ( .A(n3376), .B(n3377), .Z(n3375) );
  XOR U3177 ( .A(n3374), .B(n2962), .Z(n3377) );
  XNOR U3178 ( .A(p_input[1705]), .B(n3378), .Z(n2962) );
  AND U3179 ( .A(n134), .B(n3379), .Z(n3378) );
  XOR U3180 ( .A(p_input[1721]), .B(p_input[1705]), .Z(n3379) );
  XNOR U3181 ( .A(n2959), .B(n3374), .Z(n3376) );
  XOR U3182 ( .A(n3380), .B(n3381), .Z(n2959) );
  AND U3183 ( .A(n131), .B(n3382), .Z(n3381) );
  XOR U3184 ( .A(p_input[1689]), .B(p_input[1673]), .Z(n3382) );
  XOR U3185 ( .A(n3383), .B(n3384), .Z(n3374) );
  AND U3186 ( .A(n3385), .B(n3386), .Z(n3384) );
  XOR U3187 ( .A(n3383), .B(n2974), .Z(n3386) );
  XNOR U3188 ( .A(p_input[1704]), .B(n3387), .Z(n2974) );
  AND U3189 ( .A(n134), .B(n3388), .Z(n3387) );
  XOR U3190 ( .A(p_input[1720]), .B(p_input[1704]), .Z(n3388) );
  XNOR U3191 ( .A(n2971), .B(n3383), .Z(n3385) );
  XOR U3192 ( .A(n3389), .B(n3390), .Z(n2971) );
  AND U3193 ( .A(n131), .B(n3391), .Z(n3390) );
  XOR U3194 ( .A(p_input[1688]), .B(p_input[1672]), .Z(n3391) );
  XOR U3195 ( .A(n3392), .B(n3393), .Z(n3383) );
  AND U3196 ( .A(n3394), .B(n3395), .Z(n3393) );
  XOR U3197 ( .A(n3392), .B(n2986), .Z(n3395) );
  XNOR U3198 ( .A(p_input[1703]), .B(n3396), .Z(n2986) );
  AND U3199 ( .A(n134), .B(n3397), .Z(n3396) );
  XOR U3200 ( .A(p_input[1719]), .B(p_input[1703]), .Z(n3397) );
  XNOR U3201 ( .A(n2983), .B(n3392), .Z(n3394) );
  XOR U3202 ( .A(n3398), .B(n3399), .Z(n2983) );
  AND U3203 ( .A(n131), .B(n3400), .Z(n3399) );
  XOR U3204 ( .A(p_input[1687]), .B(p_input[1671]), .Z(n3400) );
  XOR U3205 ( .A(n3401), .B(n3402), .Z(n3392) );
  AND U3206 ( .A(n3403), .B(n3404), .Z(n3402) );
  XOR U3207 ( .A(n3401), .B(n2998), .Z(n3404) );
  XNOR U3208 ( .A(p_input[1702]), .B(n3405), .Z(n2998) );
  AND U3209 ( .A(n134), .B(n3406), .Z(n3405) );
  XOR U3210 ( .A(p_input[1718]), .B(p_input[1702]), .Z(n3406) );
  XNOR U3211 ( .A(n2995), .B(n3401), .Z(n3403) );
  XOR U3212 ( .A(n3407), .B(n3408), .Z(n2995) );
  AND U3213 ( .A(n131), .B(n3409), .Z(n3408) );
  XOR U3214 ( .A(p_input[1686]), .B(p_input[1670]), .Z(n3409) );
  XOR U3215 ( .A(n3410), .B(n3411), .Z(n3401) );
  AND U3216 ( .A(n3412), .B(n3413), .Z(n3411) );
  XOR U3217 ( .A(n3410), .B(n3010), .Z(n3413) );
  XNOR U3218 ( .A(p_input[1701]), .B(n3414), .Z(n3010) );
  AND U3219 ( .A(n134), .B(n3415), .Z(n3414) );
  XOR U3220 ( .A(p_input[1717]), .B(p_input[1701]), .Z(n3415) );
  XNOR U3221 ( .A(n3007), .B(n3410), .Z(n3412) );
  XOR U3222 ( .A(n3416), .B(n3417), .Z(n3007) );
  AND U3223 ( .A(n131), .B(n3418), .Z(n3417) );
  XOR U3224 ( .A(p_input[1685]), .B(p_input[1669]), .Z(n3418) );
  XOR U3225 ( .A(n3419), .B(n3420), .Z(n3410) );
  AND U3226 ( .A(n3421), .B(n3422), .Z(n3420) );
  XOR U3227 ( .A(n3419), .B(n3022), .Z(n3422) );
  XNOR U3228 ( .A(p_input[1700]), .B(n3423), .Z(n3022) );
  AND U3229 ( .A(n134), .B(n3424), .Z(n3423) );
  XOR U3230 ( .A(p_input[1716]), .B(p_input[1700]), .Z(n3424) );
  XNOR U3231 ( .A(n3019), .B(n3419), .Z(n3421) );
  XOR U3232 ( .A(n3425), .B(n3426), .Z(n3019) );
  AND U3233 ( .A(n131), .B(n3427), .Z(n3426) );
  XOR U3234 ( .A(p_input[1684]), .B(p_input[1668]), .Z(n3427) );
  XOR U3235 ( .A(n3428), .B(n3429), .Z(n3419) );
  AND U3236 ( .A(n3430), .B(n3431), .Z(n3429) );
  XOR U3237 ( .A(n3428), .B(n3034), .Z(n3431) );
  XNOR U3238 ( .A(p_input[1699]), .B(n3432), .Z(n3034) );
  AND U3239 ( .A(n134), .B(n3433), .Z(n3432) );
  XOR U3240 ( .A(p_input[1715]), .B(p_input[1699]), .Z(n3433) );
  XNOR U3241 ( .A(n3031), .B(n3428), .Z(n3430) );
  XOR U3242 ( .A(n3434), .B(n3435), .Z(n3031) );
  AND U3243 ( .A(n131), .B(n3436), .Z(n3435) );
  XOR U3244 ( .A(p_input[1683]), .B(p_input[1667]), .Z(n3436) );
  XOR U3245 ( .A(n3437), .B(n3438), .Z(n3428) );
  AND U3246 ( .A(n3439), .B(n3440), .Z(n3438) );
  XOR U3247 ( .A(n3046), .B(n3437), .Z(n3440) );
  XNOR U3248 ( .A(p_input[1698]), .B(n3441), .Z(n3046) );
  AND U3249 ( .A(n134), .B(n3442), .Z(n3441) );
  XOR U3250 ( .A(p_input[1714]), .B(p_input[1698]), .Z(n3442) );
  XNOR U3251 ( .A(n3437), .B(n3043), .Z(n3439) );
  XOR U3252 ( .A(n3443), .B(n3444), .Z(n3043) );
  AND U3253 ( .A(n131), .B(n3445), .Z(n3444) );
  XOR U3254 ( .A(p_input[1682]), .B(p_input[1666]), .Z(n3445) );
  XOR U3255 ( .A(n3446), .B(n3447), .Z(n3437) );
  AND U3256 ( .A(n3448), .B(n3449), .Z(n3447) );
  XNOR U3257 ( .A(n3450), .B(n3059), .Z(n3449) );
  XNOR U3258 ( .A(p_input[1697]), .B(n3451), .Z(n3059) );
  AND U3259 ( .A(n134), .B(n3452), .Z(n3451) );
  XNOR U3260 ( .A(p_input[1713]), .B(n3453), .Z(n3452) );
  IV U3261 ( .A(p_input[1697]), .Z(n3453) );
  XNOR U3262 ( .A(n3056), .B(n3446), .Z(n3448) );
  XNOR U3263 ( .A(p_input[1665]), .B(n3454), .Z(n3056) );
  AND U3264 ( .A(n131), .B(n3455), .Z(n3454) );
  XOR U3265 ( .A(p_input[1681]), .B(p_input[1665]), .Z(n3455) );
  IV U3266 ( .A(n3450), .Z(n3446) );
  AND U3267 ( .A(n3321), .B(n3324), .Z(n3450) );
  XOR U3268 ( .A(p_input[1696]), .B(n3456), .Z(n3324) );
  AND U3269 ( .A(n134), .B(n3457), .Z(n3456) );
  XOR U3270 ( .A(p_input[1712]), .B(p_input[1696]), .Z(n3457) );
  XOR U3271 ( .A(n3458), .B(n3459), .Z(n134) );
  AND U3272 ( .A(n3460), .B(n3461), .Z(n3459) );
  XNOR U3273 ( .A(p_input[1727]), .B(n3458), .Z(n3461) );
  XOR U3274 ( .A(n3458), .B(p_input[1711]), .Z(n3460) );
  XOR U3275 ( .A(n3462), .B(n3463), .Z(n3458) );
  AND U3276 ( .A(n3464), .B(n3465), .Z(n3463) );
  XNOR U3277 ( .A(p_input[1726]), .B(n3462), .Z(n3465) );
  XOR U3278 ( .A(n3462), .B(p_input[1710]), .Z(n3464) );
  XOR U3279 ( .A(n3466), .B(n3467), .Z(n3462) );
  AND U3280 ( .A(n3468), .B(n3469), .Z(n3467) );
  XNOR U3281 ( .A(p_input[1725]), .B(n3466), .Z(n3469) );
  XOR U3282 ( .A(n3466), .B(p_input[1709]), .Z(n3468) );
  XOR U3283 ( .A(n3470), .B(n3471), .Z(n3466) );
  AND U3284 ( .A(n3472), .B(n3473), .Z(n3471) );
  XNOR U3285 ( .A(p_input[1724]), .B(n3470), .Z(n3473) );
  XOR U3286 ( .A(n3470), .B(p_input[1708]), .Z(n3472) );
  XOR U3287 ( .A(n3474), .B(n3475), .Z(n3470) );
  AND U3288 ( .A(n3476), .B(n3477), .Z(n3475) );
  XNOR U3289 ( .A(p_input[1723]), .B(n3474), .Z(n3477) );
  XOR U3290 ( .A(n3474), .B(p_input[1707]), .Z(n3476) );
  XOR U3291 ( .A(n3478), .B(n3479), .Z(n3474) );
  AND U3292 ( .A(n3480), .B(n3481), .Z(n3479) );
  XNOR U3293 ( .A(p_input[1722]), .B(n3478), .Z(n3481) );
  XOR U3294 ( .A(n3478), .B(p_input[1706]), .Z(n3480) );
  XOR U3295 ( .A(n3482), .B(n3483), .Z(n3478) );
  AND U3296 ( .A(n3484), .B(n3485), .Z(n3483) );
  XNOR U3297 ( .A(p_input[1721]), .B(n3482), .Z(n3485) );
  XOR U3298 ( .A(n3482), .B(p_input[1705]), .Z(n3484) );
  XOR U3299 ( .A(n3486), .B(n3487), .Z(n3482) );
  AND U3300 ( .A(n3488), .B(n3489), .Z(n3487) );
  XNOR U3301 ( .A(p_input[1720]), .B(n3486), .Z(n3489) );
  XOR U3302 ( .A(n3486), .B(p_input[1704]), .Z(n3488) );
  XOR U3303 ( .A(n3490), .B(n3491), .Z(n3486) );
  AND U3304 ( .A(n3492), .B(n3493), .Z(n3491) );
  XNOR U3305 ( .A(p_input[1719]), .B(n3490), .Z(n3493) );
  XOR U3306 ( .A(n3490), .B(p_input[1703]), .Z(n3492) );
  XOR U3307 ( .A(n3494), .B(n3495), .Z(n3490) );
  AND U3308 ( .A(n3496), .B(n3497), .Z(n3495) );
  XNOR U3309 ( .A(p_input[1718]), .B(n3494), .Z(n3497) );
  XOR U3310 ( .A(n3494), .B(p_input[1702]), .Z(n3496) );
  XOR U3311 ( .A(n3498), .B(n3499), .Z(n3494) );
  AND U3312 ( .A(n3500), .B(n3501), .Z(n3499) );
  XNOR U3313 ( .A(p_input[1717]), .B(n3498), .Z(n3501) );
  XOR U3314 ( .A(n3498), .B(p_input[1701]), .Z(n3500) );
  XOR U3315 ( .A(n3502), .B(n3503), .Z(n3498) );
  AND U3316 ( .A(n3504), .B(n3505), .Z(n3503) );
  XNOR U3317 ( .A(p_input[1716]), .B(n3502), .Z(n3505) );
  XOR U3318 ( .A(n3502), .B(p_input[1700]), .Z(n3504) );
  XOR U3319 ( .A(n3506), .B(n3507), .Z(n3502) );
  AND U3320 ( .A(n3508), .B(n3509), .Z(n3507) );
  XNOR U3321 ( .A(p_input[1715]), .B(n3506), .Z(n3509) );
  XOR U3322 ( .A(n3506), .B(p_input[1699]), .Z(n3508) );
  XOR U3323 ( .A(n3510), .B(n3511), .Z(n3506) );
  AND U3324 ( .A(n3512), .B(n3513), .Z(n3511) );
  XNOR U3325 ( .A(p_input[1714]), .B(n3510), .Z(n3513) );
  XOR U3326 ( .A(n3510), .B(p_input[1698]), .Z(n3512) );
  XNOR U3327 ( .A(n3514), .B(n3515), .Z(n3510) );
  AND U3328 ( .A(n3516), .B(n3517), .Z(n3515) );
  XOR U3329 ( .A(p_input[1713]), .B(n3514), .Z(n3517) );
  XNOR U3330 ( .A(p_input[1697]), .B(n3514), .Z(n3516) );
  AND U3331 ( .A(p_input[1712]), .B(n3518), .Z(n3514) );
  IV U3332 ( .A(p_input[1696]), .Z(n3518) );
  XNOR U3333 ( .A(p_input[1664]), .B(n3519), .Z(n3321) );
  AND U3334 ( .A(n131), .B(n3520), .Z(n3519) );
  XOR U3335 ( .A(p_input[1680]), .B(p_input[1664]), .Z(n3520) );
  XOR U3336 ( .A(n3521), .B(n3522), .Z(n131) );
  AND U3337 ( .A(n3523), .B(n3524), .Z(n3522) );
  XNOR U3338 ( .A(p_input[1695]), .B(n3521), .Z(n3524) );
  XOR U3339 ( .A(n3521), .B(p_input[1679]), .Z(n3523) );
  XOR U3340 ( .A(n3525), .B(n3526), .Z(n3521) );
  AND U3341 ( .A(n3527), .B(n3528), .Z(n3526) );
  XNOR U3342 ( .A(p_input[1694]), .B(n3525), .Z(n3528) );
  XNOR U3343 ( .A(n3525), .B(n3335), .Z(n3527) );
  IV U3344 ( .A(p_input[1678]), .Z(n3335) );
  XOR U3345 ( .A(n3529), .B(n3530), .Z(n3525) );
  AND U3346 ( .A(n3531), .B(n3532), .Z(n3530) );
  XNOR U3347 ( .A(p_input[1693]), .B(n3529), .Z(n3532) );
  XNOR U3348 ( .A(n3529), .B(n3344), .Z(n3531) );
  IV U3349 ( .A(p_input[1677]), .Z(n3344) );
  XOR U3350 ( .A(n3533), .B(n3534), .Z(n3529) );
  AND U3351 ( .A(n3535), .B(n3536), .Z(n3534) );
  XNOR U3352 ( .A(p_input[1692]), .B(n3533), .Z(n3536) );
  XNOR U3353 ( .A(n3533), .B(n3353), .Z(n3535) );
  IV U3354 ( .A(p_input[1676]), .Z(n3353) );
  XOR U3355 ( .A(n3537), .B(n3538), .Z(n3533) );
  AND U3356 ( .A(n3539), .B(n3540), .Z(n3538) );
  XNOR U3357 ( .A(p_input[1691]), .B(n3537), .Z(n3540) );
  XNOR U3358 ( .A(n3537), .B(n3362), .Z(n3539) );
  IV U3359 ( .A(p_input[1675]), .Z(n3362) );
  XOR U3360 ( .A(n3541), .B(n3542), .Z(n3537) );
  AND U3361 ( .A(n3543), .B(n3544), .Z(n3542) );
  XNOR U3362 ( .A(p_input[1690]), .B(n3541), .Z(n3544) );
  XNOR U3363 ( .A(n3541), .B(n3371), .Z(n3543) );
  IV U3364 ( .A(p_input[1674]), .Z(n3371) );
  XOR U3365 ( .A(n3545), .B(n3546), .Z(n3541) );
  AND U3366 ( .A(n3547), .B(n3548), .Z(n3546) );
  XNOR U3367 ( .A(p_input[1689]), .B(n3545), .Z(n3548) );
  XNOR U3368 ( .A(n3545), .B(n3380), .Z(n3547) );
  IV U3369 ( .A(p_input[1673]), .Z(n3380) );
  XOR U3370 ( .A(n3549), .B(n3550), .Z(n3545) );
  AND U3371 ( .A(n3551), .B(n3552), .Z(n3550) );
  XNOR U3372 ( .A(p_input[1688]), .B(n3549), .Z(n3552) );
  XNOR U3373 ( .A(n3549), .B(n3389), .Z(n3551) );
  IV U3374 ( .A(p_input[1672]), .Z(n3389) );
  XOR U3375 ( .A(n3553), .B(n3554), .Z(n3549) );
  AND U3376 ( .A(n3555), .B(n3556), .Z(n3554) );
  XNOR U3377 ( .A(p_input[1687]), .B(n3553), .Z(n3556) );
  XNOR U3378 ( .A(n3553), .B(n3398), .Z(n3555) );
  IV U3379 ( .A(p_input[1671]), .Z(n3398) );
  XOR U3380 ( .A(n3557), .B(n3558), .Z(n3553) );
  AND U3381 ( .A(n3559), .B(n3560), .Z(n3558) );
  XNOR U3382 ( .A(p_input[1686]), .B(n3557), .Z(n3560) );
  XNOR U3383 ( .A(n3557), .B(n3407), .Z(n3559) );
  IV U3384 ( .A(p_input[1670]), .Z(n3407) );
  XOR U3385 ( .A(n3561), .B(n3562), .Z(n3557) );
  AND U3386 ( .A(n3563), .B(n3564), .Z(n3562) );
  XNOR U3387 ( .A(p_input[1685]), .B(n3561), .Z(n3564) );
  XNOR U3388 ( .A(n3561), .B(n3416), .Z(n3563) );
  IV U3389 ( .A(p_input[1669]), .Z(n3416) );
  XOR U3390 ( .A(n3565), .B(n3566), .Z(n3561) );
  AND U3391 ( .A(n3567), .B(n3568), .Z(n3566) );
  XNOR U3392 ( .A(p_input[1684]), .B(n3565), .Z(n3568) );
  XNOR U3393 ( .A(n3565), .B(n3425), .Z(n3567) );
  IV U3394 ( .A(p_input[1668]), .Z(n3425) );
  XOR U3395 ( .A(n3569), .B(n3570), .Z(n3565) );
  AND U3396 ( .A(n3571), .B(n3572), .Z(n3570) );
  XNOR U3397 ( .A(p_input[1683]), .B(n3569), .Z(n3572) );
  XNOR U3398 ( .A(n3569), .B(n3434), .Z(n3571) );
  IV U3399 ( .A(p_input[1667]), .Z(n3434) );
  XOR U3400 ( .A(n3573), .B(n3574), .Z(n3569) );
  AND U3401 ( .A(n3575), .B(n3576), .Z(n3574) );
  XNOR U3402 ( .A(p_input[1682]), .B(n3573), .Z(n3576) );
  XNOR U3403 ( .A(n3573), .B(n3443), .Z(n3575) );
  IV U3404 ( .A(p_input[1666]), .Z(n3443) );
  XNOR U3405 ( .A(n3577), .B(n3578), .Z(n3573) );
  AND U3406 ( .A(n3579), .B(n3580), .Z(n3578) );
  XOR U3407 ( .A(p_input[1681]), .B(n3577), .Z(n3580) );
  XNOR U3408 ( .A(p_input[1665]), .B(n3577), .Z(n3579) );
  AND U3409 ( .A(p_input[1680]), .B(n3581), .Z(n3577) );
  IV U3410 ( .A(p_input[1664]), .Z(n3581) );
  XOR U3411 ( .A(n3582), .B(n3583), .Z(n2697) );
  AND U3412 ( .A(n411), .B(n3584), .Z(n3583) );
  XNOR U3413 ( .A(n3585), .B(n3582), .Z(n3584) );
  XOR U3414 ( .A(n3586), .B(n3587), .Z(n411) );
  AND U3415 ( .A(n3588), .B(n3589), .Z(n3587) );
  XNOR U3416 ( .A(n2709), .B(n3586), .Z(n3589) );
  AND U3417 ( .A(n3590), .B(n3591), .Z(n2709) );
  XOR U3418 ( .A(n3586), .B(n2708), .Z(n3588) );
  AND U3419 ( .A(n3592), .B(n3593), .Z(n2708) );
  XOR U3420 ( .A(n3594), .B(n3595), .Z(n3586) );
  AND U3421 ( .A(n3596), .B(n3597), .Z(n3595) );
  XOR U3422 ( .A(n3594), .B(n2721), .Z(n3597) );
  XOR U3423 ( .A(n3598), .B(n3599), .Z(n2721) );
  AND U3424 ( .A(n242), .B(n3600), .Z(n3599) );
  XOR U3425 ( .A(n3601), .B(n3598), .Z(n3600) );
  XNOR U3426 ( .A(n2718), .B(n3594), .Z(n3596) );
  XOR U3427 ( .A(n3602), .B(n3603), .Z(n2718) );
  AND U3428 ( .A(n239), .B(n3604), .Z(n3603) );
  XOR U3429 ( .A(n3605), .B(n3602), .Z(n3604) );
  XOR U3430 ( .A(n3606), .B(n3607), .Z(n3594) );
  AND U3431 ( .A(n3608), .B(n3609), .Z(n3607) );
  XOR U3432 ( .A(n3606), .B(n2733), .Z(n3609) );
  XOR U3433 ( .A(n3610), .B(n3611), .Z(n2733) );
  AND U3434 ( .A(n242), .B(n3612), .Z(n3611) );
  XOR U3435 ( .A(n3613), .B(n3610), .Z(n3612) );
  XNOR U3436 ( .A(n2730), .B(n3606), .Z(n3608) );
  XOR U3437 ( .A(n3614), .B(n3615), .Z(n2730) );
  AND U3438 ( .A(n239), .B(n3616), .Z(n3615) );
  XOR U3439 ( .A(n3617), .B(n3614), .Z(n3616) );
  XOR U3440 ( .A(n3618), .B(n3619), .Z(n3606) );
  AND U3441 ( .A(n3620), .B(n3621), .Z(n3619) );
  XOR U3442 ( .A(n3618), .B(n2745), .Z(n3621) );
  XOR U3443 ( .A(n3622), .B(n3623), .Z(n2745) );
  AND U3444 ( .A(n242), .B(n3624), .Z(n3623) );
  XOR U3445 ( .A(n3625), .B(n3622), .Z(n3624) );
  XNOR U3446 ( .A(n2742), .B(n3618), .Z(n3620) );
  XOR U3447 ( .A(n3626), .B(n3627), .Z(n2742) );
  AND U3448 ( .A(n239), .B(n3628), .Z(n3627) );
  XOR U3449 ( .A(n3629), .B(n3626), .Z(n3628) );
  XOR U3450 ( .A(n3630), .B(n3631), .Z(n3618) );
  AND U3451 ( .A(n3632), .B(n3633), .Z(n3631) );
  XOR U3452 ( .A(n3630), .B(n2757), .Z(n3633) );
  XOR U3453 ( .A(n3634), .B(n3635), .Z(n2757) );
  AND U3454 ( .A(n242), .B(n3636), .Z(n3635) );
  XOR U3455 ( .A(n3637), .B(n3634), .Z(n3636) );
  XNOR U3456 ( .A(n2754), .B(n3630), .Z(n3632) );
  XOR U3457 ( .A(n3638), .B(n3639), .Z(n2754) );
  AND U3458 ( .A(n239), .B(n3640), .Z(n3639) );
  XOR U3459 ( .A(n3641), .B(n3638), .Z(n3640) );
  XOR U3460 ( .A(n3642), .B(n3643), .Z(n3630) );
  AND U3461 ( .A(n3644), .B(n3645), .Z(n3643) );
  XOR U3462 ( .A(n3642), .B(n2769), .Z(n3645) );
  XOR U3463 ( .A(n3646), .B(n3647), .Z(n2769) );
  AND U3464 ( .A(n242), .B(n3648), .Z(n3647) );
  XOR U3465 ( .A(n3649), .B(n3646), .Z(n3648) );
  XNOR U3466 ( .A(n2766), .B(n3642), .Z(n3644) );
  XOR U3467 ( .A(n3650), .B(n3651), .Z(n2766) );
  AND U3468 ( .A(n239), .B(n3652), .Z(n3651) );
  XOR U3469 ( .A(n3653), .B(n3650), .Z(n3652) );
  XOR U3470 ( .A(n3654), .B(n3655), .Z(n3642) );
  AND U3471 ( .A(n3656), .B(n3657), .Z(n3655) );
  XOR U3472 ( .A(n3654), .B(n2781), .Z(n3657) );
  XOR U3473 ( .A(n3658), .B(n3659), .Z(n2781) );
  AND U3474 ( .A(n242), .B(n3660), .Z(n3659) );
  XOR U3475 ( .A(n3661), .B(n3658), .Z(n3660) );
  XNOR U3476 ( .A(n2778), .B(n3654), .Z(n3656) );
  XOR U3477 ( .A(n3662), .B(n3663), .Z(n2778) );
  AND U3478 ( .A(n239), .B(n3664), .Z(n3663) );
  XOR U3479 ( .A(n3665), .B(n3662), .Z(n3664) );
  XOR U3480 ( .A(n3666), .B(n3667), .Z(n3654) );
  AND U3481 ( .A(n3668), .B(n3669), .Z(n3667) );
  XOR U3482 ( .A(n3666), .B(n2793), .Z(n3669) );
  XOR U3483 ( .A(n3670), .B(n3671), .Z(n2793) );
  AND U3484 ( .A(n242), .B(n3672), .Z(n3671) );
  XOR U3485 ( .A(n3673), .B(n3670), .Z(n3672) );
  XNOR U3486 ( .A(n2790), .B(n3666), .Z(n3668) );
  XOR U3487 ( .A(n3674), .B(n3675), .Z(n2790) );
  AND U3488 ( .A(n239), .B(n3676), .Z(n3675) );
  XOR U3489 ( .A(n3677), .B(n3674), .Z(n3676) );
  XOR U3490 ( .A(n3678), .B(n3679), .Z(n3666) );
  AND U3491 ( .A(n3680), .B(n3681), .Z(n3679) );
  XOR U3492 ( .A(n3678), .B(n2805), .Z(n3681) );
  XOR U3493 ( .A(n3682), .B(n3683), .Z(n2805) );
  AND U3494 ( .A(n242), .B(n3684), .Z(n3683) );
  XOR U3495 ( .A(n3685), .B(n3682), .Z(n3684) );
  XNOR U3496 ( .A(n2802), .B(n3678), .Z(n3680) );
  XOR U3497 ( .A(n3686), .B(n3687), .Z(n2802) );
  AND U3498 ( .A(n239), .B(n3688), .Z(n3687) );
  XOR U3499 ( .A(n3689), .B(n3686), .Z(n3688) );
  XOR U3500 ( .A(n3690), .B(n3691), .Z(n3678) );
  AND U3501 ( .A(n3692), .B(n3693), .Z(n3691) );
  XOR U3502 ( .A(n3690), .B(n2817), .Z(n3693) );
  XOR U3503 ( .A(n3694), .B(n3695), .Z(n2817) );
  AND U3504 ( .A(n242), .B(n3696), .Z(n3695) );
  XOR U3505 ( .A(n3697), .B(n3694), .Z(n3696) );
  XNOR U3506 ( .A(n2814), .B(n3690), .Z(n3692) );
  XOR U3507 ( .A(n3698), .B(n3699), .Z(n2814) );
  AND U3508 ( .A(n239), .B(n3700), .Z(n3699) );
  XOR U3509 ( .A(n3701), .B(n3698), .Z(n3700) );
  XOR U3510 ( .A(n3702), .B(n3703), .Z(n3690) );
  AND U3511 ( .A(n3704), .B(n3705), .Z(n3703) );
  XOR U3512 ( .A(n3702), .B(n2829), .Z(n3705) );
  XOR U3513 ( .A(n3706), .B(n3707), .Z(n2829) );
  AND U3514 ( .A(n242), .B(n3708), .Z(n3707) );
  XOR U3515 ( .A(n3709), .B(n3706), .Z(n3708) );
  XNOR U3516 ( .A(n2826), .B(n3702), .Z(n3704) );
  XOR U3517 ( .A(n3710), .B(n3711), .Z(n2826) );
  AND U3518 ( .A(n239), .B(n3712), .Z(n3711) );
  XOR U3519 ( .A(n3713), .B(n3710), .Z(n3712) );
  XOR U3520 ( .A(n3714), .B(n3715), .Z(n3702) );
  AND U3521 ( .A(n3716), .B(n3717), .Z(n3715) );
  XOR U3522 ( .A(n3714), .B(n2841), .Z(n3717) );
  XOR U3523 ( .A(n3718), .B(n3719), .Z(n2841) );
  AND U3524 ( .A(n242), .B(n3720), .Z(n3719) );
  XOR U3525 ( .A(n3721), .B(n3718), .Z(n3720) );
  XNOR U3526 ( .A(n2838), .B(n3714), .Z(n3716) );
  XOR U3527 ( .A(n3722), .B(n3723), .Z(n2838) );
  AND U3528 ( .A(n239), .B(n3724), .Z(n3723) );
  XOR U3529 ( .A(n3725), .B(n3722), .Z(n3724) );
  XOR U3530 ( .A(n3726), .B(n3727), .Z(n3714) );
  AND U3531 ( .A(n3728), .B(n3729), .Z(n3727) );
  XOR U3532 ( .A(n3726), .B(n2853), .Z(n3729) );
  XOR U3533 ( .A(n3730), .B(n3731), .Z(n2853) );
  AND U3534 ( .A(n242), .B(n3732), .Z(n3731) );
  XOR U3535 ( .A(n3733), .B(n3730), .Z(n3732) );
  XNOR U3536 ( .A(n2850), .B(n3726), .Z(n3728) );
  XOR U3537 ( .A(n3734), .B(n3735), .Z(n2850) );
  AND U3538 ( .A(n239), .B(n3736), .Z(n3735) );
  XOR U3539 ( .A(n3737), .B(n3734), .Z(n3736) );
  XOR U3540 ( .A(n3738), .B(n3739), .Z(n3726) );
  AND U3541 ( .A(n3740), .B(n3741), .Z(n3739) );
  XOR U3542 ( .A(n2865), .B(n3738), .Z(n3741) );
  XOR U3543 ( .A(n3742), .B(n3743), .Z(n2865) );
  AND U3544 ( .A(n242), .B(n3744), .Z(n3743) );
  XOR U3545 ( .A(n3742), .B(n3745), .Z(n3744) );
  XNOR U3546 ( .A(n3738), .B(n2862), .Z(n3740) );
  XOR U3547 ( .A(n3746), .B(n3747), .Z(n2862) );
  AND U3548 ( .A(n239), .B(n3748), .Z(n3747) );
  XOR U3549 ( .A(n3746), .B(n3749), .Z(n3748) );
  XOR U3550 ( .A(n3750), .B(n3751), .Z(n3738) );
  AND U3551 ( .A(n3752), .B(n3753), .Z(n3751) );
  XNOR U3552 ( .A(n3754), .B(n2878), .Z(n3753) );
  XOR U3553 ( .A(n3755), .B(n3756), .Z(n2878) );
  AND U3554 ( .A(n242), .B(n3757), .Z(n3756) );
  XOR U3555 ( .A(n3758), .B(n3755), .Z(n3757) );
  XNOR U3556 ( .A(n2875), .B(n3750), .Z(n3752) );
  XOR U3557 ( .A(n3759), .B(n3760), .Z(n2875) );
  AND U3558 ( .A(n239), .B(n3761), .Z(n3760) );
  XOR U3559 ( .A(n3762), .B(n3759), .Z(n3761) );
  IV U3560 ( .A(n3754), .Z(n3750) );
  AND U3561 ( .A(n3582), .B(n3585), .Z(n3754) );
  XNOR U3562 ( .A(n3763), .B(n3764), .Z(n3585) );
  AND U3563 ( .A(n242), .B(n3765), .Z(n3764) );
  XNOR U3564 ( .A(n3766), .B(n3763), .Z(n3765) );
  XOR U3565 ( .A(n3767), .B(n3768), .Z(n242) );
  AND U3566 ( .A(n3769), .B(n3770), .Z(n3768) );
  XNOR U3567 ( .A(n3590), .B(n3767), .Z(n3770) );
  AND U3568 ( .A(p_input[1663]), .B(p_input[1647]), .Z(n3590) );
  XOR U3569 ( .A(n3767), .B(n3591), .Z(n3769) );
  AND U3570 ( .A(p_input[1631]), .B(p_input[1615]), .Z(n3591) );
  XOR U3571 ( .A(n3771), .B(n3772), .Z(n3767) );
  AND U3572 ( .A(n3773), .B(n3774), .Z(n3772) );
  XOR U3573 ( .A(n3771), .B(n3601), .Z(n3774) );
  XNOR U3574 ( .A(p_input[1646]), .B(n3775), .Z(n3601) );
  AND U3575 ( .A(n142), .B(n3776), .Z(n3775) );
  XOR U3576 ( .A(p_input[1662]), .B(p_input[1646]), .Z(n3776) );
  XNOR U3577 ( .A(n3598), .B(n3771), .Z(n3773) );
  XOR U3578 ( .A(n3777), .B(n3778), .Z(n3598) );
  AND U3579 ( .A(n140), .B(n3779), .Z(n3778) );
  XOR U3580 ( .A(p_input[1630]), .B(p_input[1614]), .Z(n3779) );
  XOR U3581 ( .A(n3780), .B(n3781), .Z(n3771) );
  AND U3582 ( .A(n3782), .B(n3783), .Z(n3781) );
  XOR U3583 ( .A(n3780), .B(n3613), .Z(n3783) );
  XNOR U3584 ( .A(p_input[1645]), .B(n3784), .Z(n3613) );
  AND U3585 ( .A(n142), .B(n3785), .Z(n3784) );
  XOR U3586 ( .A(p_input[1661]), .B(p_input[1645]), .Z(n3785) );
  XNOR U3587 ( .A(n3610), .B(n3780), .Z(n3782) );
  XOR U3588 ( .A(n3786), .B(n3787), .Z(n3610) );
  AND U3589 ( .A(n140), .B(n3788), .Z(n3787) );
  XOR U3590 ( .A(p_input[1629]), .B(p_input[1613]), .Z(n3788) );
  XOR U3591 ( .A(n3789), .B(n3790), .Z(n3780) );
  AND U3592 ( .A(n3791), .B(n3792), .Z(n3790) );
  XOR U3593 ( .A(n3789), .B(n3625), .Z(n3792) );
  XNOR U3594 ( .A(p_input[1644]), .B(n3793), .Z(n3625) );
  AND U3595 ( .A(n142), .B(n3794), .Z(n3793) );
  XOR U3596 ( .A(p_input[1660]), .B(p_input[1644]), .Z(n3794) );
  XNOR U3597 ( .A(n3622), .B(n3789), .Z(n3791) );
  XOR U3598 ( .A(n3795), .B(n3796), .Z(n3622) );
  AND U3599 ( .A(n140), .B(n3797), .Z(n3796) );
  XOR U3600 ( .A(p_input[1628]), .B(p_input[1612]), .Z(n3797) );
  XOR U3601 ( .A(n3798), .B(n3799), .Z(n3789) );
  AND U3602 ( .A(n3800), .B(n3801), .Z(n3799) );
  XOR U3603 ( .A(n3798), .B(n3637), .Z(n3801) );
  XNOR U3604 ( .A(p_input[1643]), .B(n3802), .Z(n3637) );
  AND U3605 ( .A(n142), .B(n3803), .Z(n3802) );
  XOR U3606 ( .A(p_input[1659]), .B(p_input[1643]), .Z(n3803) );
  XNOR U3607 ( .A(n3634), .B(n3798), .Z(n3800) );
  XOR U3608 ( .A(n3804), .B(n3805), .Z(n3634) );
  AND U3609 ( .A(n140), .B(n3806), .Z(n3805) );
  XOR U3610 ( .A(p_input[1627]), .B(p_input[1611]), .Z(n3806) );
  XOR U3611 ( .A(n3807), .B(n3808), .Z(n3798) );
  AND U3612 ( .A(n3809), .B(n3810), .Z(n3808) );
  XOR U3613 ( .A(n3807), .B(n3649), .Z(n3810) );
  XNOR U3614 ( .A(p_input[1642]), .B(n3811), .Z(n3649) );
  AND U3615 ( .A(n142), .B(n3812), .Z(n3811) );
  XOR U3616 ( .A(p_input[1658]), .B(p_input[1642]), .Z(n3812) );
  XNOR U3617 ( .A(n3646), .B(n3807), .Z(n3809) );
  XOR U3618 ( .A(n3813), .B(n3814), .Z(n3646) );
  AND U3619 ( .A(n140), .B(n3815), .Z(n3814) );
  XOR U3620 ( .A(p_input[1626]), .B(p_input[1610]), .Z(n3815) );
  XOR U3621 ( .A(n3816), .B(n3817), .Z(n3807) );
  AND U3622 ( .A(n3818), .B(n3819), .Z(n3817) );
  XOR U3623 ( .A(n3816), .B(n3661), .Z(n3819) );
  XNOR U3624 ( .A(p_input[1641]), .B(n3820), .Z(n3661) );
  AND U3625 ( .A(n142), .B(n3821), .Z(n3820) );
  XOR U3626 ( .A(p_input[1657]), .B(p_input[1641]), .Z(n3821) );
  XNOR U3627 ( .A(n3658), .B(n3816), .Z(n3818) );
  XOR U3628 ( .A(n3822), .B(n3823), .Z(n3658) );
  AND U3629 ( .A(n140), .B(n3824), .Z(n3823) );
  XOR U3630 ( .A(p_input[1625]), .B(p_input[1609]), .Z(n3824) );
  XOR U3631 ( .A(n3825), .B(n3826), .Z(n3816) );
  AND U3632 ( .A(n3827), .B(n3828), .Z(n3826) );
  XOR U3633 ( .A(n3825), .B(n3673), .Z(n3828) );
  XNOR U3634 ( .A(p_input[1640]), .B(n3829), .Z(n3673) );
  AND U3635 ( .A(n142), .B(n3830), .Z(n3829) );
  XOR U3636 ( .A(p_input[1656]), .B(p_input[1640]), .Z(n3830) );
  XNOR U3637 ( .A(n3670), .B(n3825), .Z(n3827) );
  XOR U3638 ( .A(n3831), .B(n3832), .Z(n3670) );
  AND U3639 ( .A(n140), .B(n3833), .Z(n3832) );
  XOR U3640 ( .A(p_input[1624]), .B(p_input[1608]), .Z(n3833) );
  XOR U3641 ( .A(n3834), .B(n3835), .Z(n3825) );
  AND U3642 ( .A(n3836), .B(n3837), .Z(n3835) );
  XOR U3643 ( .A(n3834), .B(n3685), .Z(n3837) );
  XNOR U3644 ( .A(p_input[1639]), .B(n3838), .Z(n3685) );
  AND U3645 ( .A(n142), .B(n3839), .Z(n3838) );
  XOR U3646 ( .A(p_input[1655]), .B(p_input[1639]), .Z(n3839) );
  XNOR U3647 ( .A(n3682), .B(n3834), .Z(n3836) );
  XOR U3648 ( .A(n3840), .B(n3841), .Z(n3682) );
  AND U3649 ( .A(n140), .B(n3842), .Z(n3841) );
  XOR U3650 ( .A(p_input[1623]), .B(p_input[1607]), .Z(n3842) );
  XOR U3651 ( .A(n3843), .B(n3844), .Z(n3834) );
  AND U3652 ( .A(n3845), .B(n3846), .Z(n3844) );
  XOR U3653 ( .A(n3843), .B(n3697), .Z(n3846) );
  XNOR U3654 ( .A(p_input[1638]), .B(n3847), .Z(n3697) );
  AND U3655 ( .A(n142), .B(n3848), .Z(n3847) );
  XOR U3656 ( .A(p_input[1654]), .B(p_input[1638]), .Z(n3848) );
  XNOR U3657 ( .A(n3694), .B(n3843), .Z(n3845) );
  XOR U3658 ( .A(n3849), .B(n3850), .Z(n3694) );
  AND U3659 ( .A(n140), .B(n3851), .Z(n3850) );
  XOR U3660 ( .A(p_input[1622]), .B(p_input[1606]), .Z(n3851) );
  XOR U3661 ( .A(n3852), .B(n3853), .Z(n3843) );
  AND U3662 ( .A(n3854), .B(n3855), .Z(n3853) );
  XOR U3663 ( .A(n3852), .B(n3709), .Z(n3855) );
  XNOR U3664 ( .A(p_input[1637]), .B(n3856), .Z(n3709) );
  AND U3665 ( .A(n142), .B(n3857), .Z(n3856) );
  XOR U3666 ( .A(p_input[1653]), .B(p_input[1637]), .Z(n3857) );
  XNOR U3667 ( .A(n3706), .B(n3852), .Z(n3854) );
  XOR U3668 ( .A(n3858), .B(n3859), .Z(n3706) );
  AND U3669 ( .A(n140), .B(n3860), .Z(n3859) );
  XOR U3670 ( .A(p_input[1621]), .B(p_input[1605]), .Z(n3860) );
  XOR U3671 ( .A(n3861), .B(n3862), .Z(n3852) );
  AND U3672 ( .A(n3863), .B(n3864), .Z(n3862) );
  XOR U3673 ( .A(n3861), .B(n3721), .Z(n3864) );
  XNOR U3674 ( .A(p_input[1636]), .B(n3865), .Z(n3721) );
  AND U3675 ( .A(n142), .B(n3866), .Z(n3865) );
  XOR U3676 ( .A(p_input[1652]), .B(p_input[1636]), .Z(n3866) );
  XNOR U3677 ( .A(n3718), .B(n3861), .Z(n3863) );
  XOR U3678 ( .A(n3867), .B(n3868), .Z(n3718) );
  AND U3679 ( .A(n140), .B(n3869), .Z(n3868) );
  XOR U3680 ( .A(p_input[1620]), .B(p_input[1604]), .Z(n3869) );
  XOR U3681 ( .A(n3870), .B(n3871), .Z(n3861) );
  AND U3682 ( .A(n3872), .B(n3873), .Z(n3871) );
  XOR U3683 ( .A(n3870), .B(n3733), .Z(n3873) );
  XNOR U3684 ( .A(p_input[1635]), .B(n3874), .Z(n3733) );
  AND U3685 ( .A(n142), .B(n3875), .Z(n3874) );
  XOR U3686 ( .A(p_input[1651]), .B(p_input[1635]), .Z(n3875) );
  XNOR U3687 ( .A(n3730), .B(n3870), .Z(n3872) );
  XOR U3688 ( .A(n3876), .B(n3877), .Z(n3730) );
  AND U3689 ( .A(n140), .B(n3878), .Z(n3877) );
  XOR U3690 ( .A(p_input[1619]), .B(p_input[1603]), .Z(n3878) );
  XOR U3691 ( .A(n3879), .B(n3880), .Z(n3870) );
  AND U3692 ( .A(n3881), .B(n3882), .Z(n3880) );
  XOR U3693 ( .A(n3745), .B(n3879), .Z(n3882) );
  XNOR U3694 ( .A(p_input[1634]), .B(n3883), .Z(n3745) );
  AND U3695 ( .A(n142), .B(n3884), .Z(n3883) );
  XOR U3696 ( .A(p_input[1650]), .B(p_input[1634]), .Z(n3884) );
  XNOR U3697 ( .A(n3879), .B(n3742), .Z(n3881) );
  XOR U3698 ( .A(n3885), .B(n3886), .Z(n3742) );
  AND U3699 ( .A(n140), .B(n3887), .Z(n3886) );
  XOR U3700 ( .A(p_input[1618]), .B(p_input[1602]), .Z(n3887) );
  XOR U3701 ( .A(n3888), .B(n3889), .Z(n3879) );
  AND U3702 ( .A(n3890), .B(n3891), .Z(n3889) );
  XNOR U3703 ( .A(n3892), .B(n3758), .Z(n3891) );
  XNOR U3704 ( .A(p_input[1633]), .B(n3893), .Z(n3758) );
  AND U3705 ( .A(n142), .B(n3894), .Z(n3893) );
  XNOR U3706 ( .A(p_input[1649]), .B(n3895), .Z(n3894) );
  IV U3707 ( .A(p_input[1633]), .Z(n3895) );
  XNOR U3708 ( .A(n3755), .B(n3888), .Z(n3890) );
  XNOR U3709 ( .A(p_input[1601]), .B(n3896), .Z(n3755) );
  AND U3710 ( .A(n140), .B(n3897), .Z(n3896) );
  XOR U3711 ( .A(p_input[1617]), .B(p_input[1601]), .Z(n3897) );
  IV U3712 ( .A(n3892), .Z(n3888) );
  AND U3713 ( .A(n3763), .B(n3766), .Z(n3892) );
  XOR U3714 ( .A(p_input[1632]), .B(n3898), .Z(n3766) );
  AND U3715 ( .A(n142), .B(n3899), .Z(n3898) );
  XOR U3716 ( .A(p_input[1648]), .B(p_input[1632]), .Z(n3899) );
  XOR U3717 ( .A(n3900), .B(n3901), .Z(n142) );
  AND U3718 ( .A(n3902), .B(n3903), .Z(n3901) );
  XNOR U3719 ( .A(p_input[1663]), .B(n3900), .Z(n3903) );
  XOR U3720 ( .A(n3900), .B(p_input[1647]), .Z(n3902) );
  XOR U3721 ( .A(n3904), .B(n3905), .Z(n3900) );
  AND U3722 ( .A(n3906), .B(n3907), .Z(n3905) );
  XNOR U3723 ( .A(p_input[1662]), .B(n3904), .Z(n3907) );
  XOR U3724 ( .A(n3904), .B(p_input[1646]), .Z(n3906) );
  XOR U3725 ( .A(n3908), .B(n3909), .Z(n3904) );
  AND U3726 ( .A(n3910), .B(n3911), .Z(n3909) );
  XNOR U3727 ( .A(p_input[1661]), .B(n3908), .Z(n3911) );
  XOR U3728 ( .A(n3908), .B(p_input[1645]), .Z(n3910) );
  XOR U3729 ( .A(n3912), .B(n3913), .Z(n3908) );
  AND U3730 ( .A(n3914), .B(n3915), .Z(n3913) );
  XNOR U3731 ( .A(p_input[1660]), .B(n3912), .Z(n3915) );
  XOR U3732 ( .A(n3912), .B(p_input[1644]), .Z(n3914) );
  XOR U3733 ( .A(n3916), .B(n3917), .Z(n3912) );
  AND U3734 ( .A(n3918), .B(n3919), .Z(n3917) );
  XNOR U3735 ( .A(p_input[1659]), .B(n3916), .Z(n3919) );
  XOR U3736 ( .A(n3916), .B(p_input[1643]), .Z(n3918) );
  XOR U3737 ( .A(n3920), .B(n3921), .Z(n3916) );
  AND U3738 ( .A(n3922), .B(n3923), .Z(n3921) );
  XNOR U3739 ( .A(p_input[1658]), .B(n3920), .Z(n3923) );
  XOR U3740 ( .A(n3920), .B(p_input[1642]), .Z(n3922) );
  XOR U3741 ( .A(n3924), .B(n3925), .Z(n3920) );
  AND U3742 ( .A(n3926), .B(n3927), .Z(n3925) );
  XNOR U3743 ( .A(p_input[1657]), .B(n3924), .Z(n3927) );
  XOR U3744 ( .A(n3924), .B(p_input[1641]), .Z(n3926) );
  XOR U3745 ( .A(n3928), .B(n3929), .Z(n3924) );
  AND U3746 ( .A(n3930), .B(n3931), .Z(n3929) );
  XNOR U3747 ( .A(p_input[1656]), .B(n3928), .Z(n3931) );
  XOR U3748 ( .A(n3928), .B(p_input[1640]), .Z(n3930) );
  XOR U3749 ( .A(n3932), .B(n3933), .Z(n3928) );
  AND U3750 ( .A(n3934), .B(n3935), .Z(n3933) );
  XNOR U3751 ( .A(p_input[1655]), .B(n3932), .Z(n3935) );
  XOR U3752 ( .A(n3932), .B(p_input[1639]), .Z(n3934) );
  XOR U3753 ( .A(n3936), .B(n3937), .Z(n3932) );
  AND U3754 ( .A(n3938), .B(n3939), .Z(n3937) );
  XNOR U3755 ( .A(p_input[1654]), .B(n3936), .Z(n3939) );
  XOR U3756 ( .A(n3936), .B(p_input[1638]), .Z(n3938) );
  XOR U3757 ( .A(n3940), .B(n3941), .Z(n3936) );
  AND U3758 ( .A(n3942), .B(n3943), .Z(n3941) );
  XNOR U3759 ( .A(p_input[1653]), .B(n3940), .Z(n3943) );
  XOR U3760 ( .A(n3940), .B(p_input[1637]), .Z(n3942) );
  XOR U3761 ( .A(n3944), .B(n3945), .Z(n3940) );
  AND U3762 ( .A(n3946), .B(n3947), .Z(n3945) );
  XNOR U3763 ( .A(p_input[1652]), .B(n3944), .Z(n3947) );
  XOR U3764 ( .A(n3944), .B(p_input[1636]), .Z(n3946) );
  XOR U3765 ( .A(n3948), .B(n3949), .Z(n3944) );
  AND U3766 ( .A(n3950), .B(n3951), .Z(n3949) );
  XNOR U3767 ( .A(p_input[1651]), .B(n3948), .Z(n3951) );
  XOR U3768 ( .A(n3948), .B(p_input[1635]), .Z(n3950) );
  XOR U3769 ( .A(n3952), .B(n3953), .Z(n3948) );
  AND U3770 ( .A(n3954), .B(n3955), .Z(n3953) );
  XNOR U3771 ( .A(p_input[1650]), .B(n3952), .Z(n3955) );
  XOR U3772 ( .A(n3952), .B(p_input[1634]), .Z(n3954) );
  XNOR U3773 ( .A(n3956), .B(n3957), .Z(n3952) );
  AND U3774 ( .A(n3958), .B(n3959), .Z(n3957) );
  XOR U3775 ( .A(p_input[1649]), .B(n3956), .Z(n3959) );
  XNOR U3776 ( .A(p_input[1633]), .B(n3956), .Z(n3958) );
  AND U3777 ( .A(p_input[1648]), .B(n3960), .Z(n3956) );
  IV U3778 ( .A(p_input[1632]), .Z(n3960) );
  XNOR U3779 ( .A(p_input[1600]), .B(n3961), .Z(n3763) );
  AND U3780 ( .A(n140), .B(n3962), .Z(n3961) );
  XOR U3781 ( .A(p_input[1616]), .B(p_input[1600]), .Z(n3962) );
  XOR U3782 ( .A(n3963), .B(n3964), .Z(n140) );
  AND U3783 ( .A(n3965), .B(n3966), .Z(n3964) );
  XNOR U3784 ( .A(p_input[1631]), .B(n3963), .Z(n3966) );
  XOR U3785 ( .A(n3963), .B(p_input[1615]), .Z(n3965) );
  XOR U3786 ( .A(n3967), .B(n3968), .Z(n3963) );
  AND U3787 ( .A(n3969), .B(n3970), .Z(n3968) );
  XNOR U3788 ( .A(p_input[1630]), .B(n3967), .Z(n3970) );
  XNOR U3789 ( .A(n3967), .B(n3777), .Z(n3969) );
  IV U3790 ( .A(p_input[1614]), .Z(n3777) );
  XOR U3791 ( .A(n3971), .B(n3972), .Z(n3967) );
  AND U3792 ( .A(n3973), .B(n3974), .Z(n3972) );
  XNOR U3793 ( .A(p_input[1629]), .B(n3971), .Z(n3974) );
  XNOR U3794 ( .A(n3971), .B(n3786), .Z(n3973) );
  IV U3795 ( .A(p_input[1613]), .Z(n3786) );
  XOR U3796 ( .A(n3975), .B(n3976), .Z(n3971) );
  AND U3797 ( .A(n3977), .B(n3978), .Z(n3976) );
  XNOR U3798 ( .A(p_input[1628]), .B(n3975), .Z(n3978) );
  XNOR U3799 ( .A(n3975), .B(n3795), .Z(n3977) );
  IV U3800 ( .A(p_input[1612]), .Z(n3795) );
  XOR U3801 ( .A(n3979), .B(n3980), .Z(n3975) );
  AND U3802 ( .A(n3981), .B(n3982), .Z(n3980) );
  XNOR U3803 ( .A(p_input[1627]), .B(n3979), .Z(n3982) );
  XNOR U3804 ( .A(n3979), .B(n3804), .Z(n3981) );
  IV U3805 ( .A(p_input[1611]), .Z(n3804) );
  XOR U3806 ( .A(n3983), .B(n3984), .Z(n3979) );
  AND U3807 ( .A(n3985), .B(n3986), .Z(n3984) );
  XNOR U3808 ( .A(p_input[1626]), .B(n3983), .Z(n3986) );
  XNOR U3809 ( .A(n3983), .B(n3813), .Z(n3985) );
  IV U3810 ( .A(p_input[1610]), .Z(n3813) );
  XOR U3811 ( .A(n3987), .B(n3988), .Z(n3983) );
  AND U3812 ( .A(n3989), .B(n3990), .Z(n3988) );
  XNOR U3813 ( .A(p_input[1625]), .B(n3987), .Z(n3990) );
  XNOR U3814 ( .A(n3987), .B(n3822), .Z(n3989) );
  IV U3815 ( .A(p_input[1609]), .Z(n3822) );
  XOR U3816 ( .A(n3991), .B(n3992), .Z(n3987) );
  AND U3817 ( .A(n3993), .B(n3994), .Z(n3992) );
  XNOR U3818 ( .A(p_input[1624]), .B(n3991), .Z(n3994) );
  XNOR U3819 ( .A(n3991), .B(n3831), .Z(n3993) );
  IV U3820 ( .A(p_input[1608]), .Z(n3831) );
  XOR U3821 ( .A(n3995), .B(n3996), .Z(n3991) );
  AND U3822 ( .A(n3997), .B(n3998), .Z(n3996) );
  XNOR U3823 ( .A(p_input[1623]), .B(n3995), .Z(n3998) );
  XNOR U3824 ( .A(n3995), .B(n3840), .Z(n3997) );
  IV U3825 ( .A(p_input[1607]), .Z(n3840) );
  XOR U3826 ( .A(n3999), .B(n4000), .Z(n3995) );
  AND U3827 ( .A(n4001), .B(n4002), .Z(n4000) );
  XNOR U3828 ( .A(p_input[1622]), .B(n3999), .Z(n4002) );
  XNOR U3829 ( .A(n3999), .B(n3849), .Z(n4001) );
  IV U3830 ( .A(p_input[1606]), .Z(n3849) );
  XOR U3831 ( .A(n4003), .B(n4004), .Z(n3999) );
  AND U3832 ( .A(n4005), .B(n4006), .Z(n4004) );
  XNOR U3833 ( .A(p_input[1621]), .B(n4003), .Z(n4006) );
  XNOR U3834 ( .A(n4003), .B(n3858), .Z(n4005) );
  IV U3835 ( .A(p_input[1605]), .Z(n3858) );
  XOR U3836 ( .A(n4007), .B(n4008), .Z(n4003) );
  AND U3837 ( .A(n4009), .B(n4010), .Z(n4008) );
  XNOR U3838 ( .A(p_input[1620]), .B(n4007), .Z(n4010) );
  XNOR U3839 ( .A(n4007), .B(n3867), .Z(n4009) );
  IV U3840 ( .A(p_input[1604]), .Z(n3867) );
  XOR U3841 ( .A(n4011), .B(n4012), .Z(n4007) );
  AND U3842 ( .A(n4013), .B(n4014), .Z(n4012) );
  XNOR U3843 ( .A(p_input[1619]), .B(n4011), .Z(n4014) );
  XNOR U3844 ( .A(n4011), .B(n3876), .Z(n4013) );
  IV U3845 ( .A(p_input[1603]), .Z(n3876) );
  XOR U3846 ( .A(n4015), .B(n4016), .Z(n4011) );
  AND U3847 ( .A(n4017), .B(n4018), .Z(n4016) );
  XNOR U3848 ( .A(p_input[1618]), .B(n4015), .Z(n4018) );
  XNOR U3849 ( .A(n4015), .B(n3885), .Z(n4017) );
  IV U3850 ( .A(p_input[1602]), .Z(n3885) );
  XNOR U3851 ( .A(n4019), .B(n4020), .Z(n4015) );
  AND U3852 ( .A(n4021), .B(n4022), .Z(n4020) );
  XOR U3853 ( .A(p_input[1617]), .B(n4019), .Z(n4022) );
  XNOR U3854 ( .A(p_input[1601]), .B(n4019), .Z(n4021) );
  AND U3855 ( .A(p_input[1616]), .B(n4023), .Z(n4019) );
  IV U3856 ( .A(p_input[1600]), .Z(n4023) );
  XOR U3857 ( .A(n4024), .B(n4025), .Z(n3582) );
  AND U3858 ( .A(n239), .B(n4026), .Z(n4025) );
  XNOR U3859 ( .A(n4027), .B(n4024), .Z(n4026) );
  XOR U3860 ( .A(n4028), .B(n4029), .Z(n239) );
  AND U3861 ( .A(n4030), .B(n4031), .Z(n4029) );
  XNOR U3862 ( .A(n3593), .B(n4028), .Z(n4031) );
  AND U3863 ( .A(p_input[1599]), .B(p_input[1583]), .Z(n3593) );
  XOR U3864 ( .A(n4028), .B(n3592), .Z(n4030) );
  AND U3865 ( .A(p_input[1551]), .B(p_input[1567]), .Z(n3592) );
  XOR U3866 ( .A(n4032), .B(n4033), .Z(n4028) );
  AND U3867 ( .A(n4034), .B(n4035), .Z(n4033) );
  XOR U3868 ( .A(n4032), .B(n3605), .Z(n4035) );
  XNOR U3869 ( .A(p_input[1582]), .B(n4036), .Z(n3605) );
  AND U3870 ( .A(n146), .B(n4037), .Z(n4036) );
  XOR U3871 ( .A(p_input[1598]), .B(p_input[1582]), .Z(n4037) );
  XNOR U3872 ( .A(n3602), .B(n4032), .Z(n4034) );
  XOR U3873 ( .A(n4038), .B(n4039), .Z(n3602) );
  AND U3874 ( .A(n143), .B(n4040), .Z(n4039) );
  XOR U3875 ( .A(p_input[1566]), .B(p_input[1550]), .Z(n4040) );
  XOR U3876 ( .A(n4041), .B(n4042), .Z(n4032) );
  AND U3877 ( .A(n4043), .B(n4044), .Z(n4042) );
  XOR U3878 ( .A(n4041), .B(n3617), .Z(n4044) );
  XNOR U3879 ( .A(p_input[1581]), .B(n4045), .Z(n3617) );
  AND U3880 ( .A(n146), .B(n4046), .Z(n4045) );
  XOR U3881 ( .A(p_input[1597]), .B(p_input[1581]), .Z(n4046) );
  XNOR U3882 ( .A(n3614), .B(n4041), .Z(n4043) );
  XOR U3883 ( .A(n4047), .B(n4048), .Z(n3614) );
  AND U3884 ( .A(n143), .B(n4049), .Z(n4048) );
  XOR U3885 ( .A(p_input[1565]), .B(p_input[1549]), .Z(n4049) );
  XOR U3886 ( .A(n4050), .B(n4051), .Z(n4041) );
  AND U3887 ( .A(n4052), .B(n4053), .Z(n4051) );
  XOR U3888 ( .A(n4050), .B(n3629), .Z(n4053) );
  XNOR U3889 ( .A(p_input[1580]), .B(n4054), .Z(n3629) );
  AND U3890 ( .A(n146), .B(n4055), .Z(n4054) );
  XOR U3891 ( .A(p_input[1596]), .B(p_input[1580]), .Z(n4055) );
  XNOR U3892 ( .A(n3626), .B(n4050), .Z(n4052) );
  XOR U3893 ( .A(n4056), .B(n4057), .Z(n3626) );
  AND U3894 ( .A(n143), .B(n4058), .Z(n4057) );
  XOR U3895 ( .A(p_input[1564]), .B(p_input[1548]), .Z(n4058) );
  XOR U3896 ( .A(n4059), .B(n4060), .Z(n4050) );
  AND U3897 ( .A(n4061), .B(n4062), .Z(n4060) );
  XOR U3898 ( .A(n4059), .B(n3641), .Z(n4062) );
  XNOR U3899 ( .A(p_input[1579]), .B(n4063), .Z(n3641) );
  AND U3900 ( .A(n146), .B(n4064), .Z(n4063) );
  XOR U3901 ( .A(p_input[1595]), .B(p_input[1579]), .Z(n4064) );
  XNOR U3902 ( .A(n3638), .B(n4059), .Z(n4061) );
  XOR U3903 ( .A(n4065), .B(n4066), .Z(n3638) );
  AND U3904 ( .A(n143), .B(n4067), .Z(n4066) );
  XOR U3905 ( .A(p_input[1563]), .B(p_input[1547]), .Z(n4067) );
  XOR U3906 ( .A(n4068), .B(n4069), .Z(n4059) );
  AND U3907 ( .A(n4070), .B(n4071), .Z(n4069) );
  XOR U3908 ( .A(n4068), .B(n3653), .Z(n4071) );
  XNOR U3909 ( .A(p_input[1578]), .B(n4072), .Z(n3653) );
  AND U3910 ( .A(n146), .B(n4073), .Z(n4072) );
  XOR U3911 ( .A(p_input[1594]), .B(p_input[1578]), .Z(n4073) );
  XNOR U3912 ( .A(n3650), .B(n4068), .Z(n4070) );
  XOR U3913 ( .A(n4074), .B(n4075), .Z(n3650) );
  AND U3914 ( .A(n143), .B(n4076), .Z(n4075) );
  XOR U3915 ( .A(p_input[1562]), .B(p_input[1546]), .Z(n4076) );
  XOR U3916 ( .A(n4077), .B(n4078), .Z(n4068) );
  AND U3917 ( .A(n4079), .B(n4080), .Z(n4078) );
  XOR U3918 ( .A(n4077), .B(n3665), .Z(n4080) );
  XNOR U3919 ( .A(p_input[1577]), .B(n4081), .Z(n3665) );
  AND U3920 ( .A(n146), .B(n4082), .Z(n4081) );
  XOR U3921 ( .A(p_input[1593]), .B(p_input[1577]), .Z(n4082) );
  XNOR U3922 ( .A(n3662), .B(n4077), .Z(n4079) );
  XOR U3923 ( .A(n4083), .B(n4084), .Z(n3662) );
  AND U3924 ( .A(n143), .B(n4085), .Z(n4084) );
  XOR U3925 ( .A(p_input[1561]), .B(p_input[1545]), .Z(n4085) );
  XOR U3926 ( .A(n4086), .B(n4087), .Z(n4077) );
  AND U3927 ( .A(n4088), .B(n4089), .Z(n4087) );
  XOR U3928 ( .A(n4086), .B(n3677), .Z(n4089) );
  XNOR U3929 ( .A(p_input[1576]), .B(n4090), .Z(n3677) );
  AND U3930 ( .A(n146), .B(n4091), .Z(n4090) );
  XOR U3931 ( .A(p_input[1592]), .B(p_input[1576]), .Z(n4091) );
  XNOR U3932 ( .A(n3674), .B(n4086), .Z(n4088) );
  XOR U3933 ( .A(n4092), .B(n4093), .Z(n3674) );
  AND U3934 ( .A(n143), .B(n4094), .Z(n4093) );
  XOR U3935 ( .A(p_input[1560]), .B(p_input[1544]), .Z(n4094) );
  XOR U3936 ( .A(n4095), .B(n4096), .Z(n4086) );
  AND U3937 ( .A(n4097), .B(n4098), .Z(n4096) );
  XOR U3938 ( .A(n4095), .B(n3689), .Z(n4098) );
  XNOR U3939 ( .A(p_input[1575]), .B(n4099), .Z(n3689) );
  AND U3940 ( .A(n146), .B(n4100), .Z(n4099) );
  XOR U3941 ( .A(p_input[1591]), .B(p_input[1575]), .Z(n4100) );
  XNOR U3942 ( .A(n3686), .B(n4095), .Z(n4097) );
  XOR U3943 ( .A(n4101), .B(n4102), .Z(n3686) );
  AND U3944 ( .A(n143), .B(n4103), .Z(n4102) );
  XOR U3945 ( .A(p_input[1559]), .B(p_input[1543]), .Z(n4103) );
  XOR U3946 ( .A(n4104), .B(n4105), .Z(n4095) );
  AND U3947 ( .A(n4106), .B(n4107), .Z(n4105) );
  XOR U3948 ( .A(n4104), .B(n3701), .Z(n4107) );
  XNOR U3949 ( .A(p_input[1574]), .B(n4108), .Z(n3701) );
  AND U3950 ( .A(n146), .B(n4109), .Z(n4108) );
  XOR U3951 ( .A(p_input[1590]), .B(p_input[1574]), .Z(n4109) );
  XNOR U3952 ( .A(n3698), .B(n4104), .Z(n4106) );
  XOR U3953 ( .A(n4110), .B(n4111), .Z(n3698) );
  AND U3954 ( .A(n143), .B(n4112), .Z(n4111) );
  XOR U3955 ( .A(p_input[1558]), .B(p_input[1542]), .Z(n4112) );
  XOR U3956 ( .A(n4113), .B(n4114), .Z(n4104) );
  AND U3957 ( .A(n4115), .B(n4116), .Z(n4114) );
  XOR U3958 ( .A(n4113), .B(n3713), .Z(n4116) );
  XNOR U3959 ( .A(p_input[1573]), .B(n4117), .Z(n3713) );
  AND U3960 ( .A(n146), .B(n4118), .Z(n4117) );
  XOR U3961 ( .A(p_input[1589]), .B(p_input[1573]), .Z(n4118) );
  XNOR U3962 ( .A(n3710), .B(n4113), .Z(n4115) );
  XOR U3963 ( .A(n4119), .B(n4120), .Z(n3710) );
  AND U3964 ( .A(n143), .B(n4121), .Z(n4120) );
  XOR U3965 ( .A(p_input[1557]), .B(p_input[1541]), .Z(n4121) );
  XOR U3966 ( .A(n4122), .B(n4123), .Z(n4113) );
  AND U3967 ( .A(n4124), .B(n4125), .Z(n4123) );
  XOR U3968 ( .A(n4122), .B(n3725), .Z(n4125) );
  XNOR U3969 ( .A(p_input[1572]), .B(n4126), .Z(n3725) );
  AND U3970 ( .A(n146), .B(n4127), .Z(n4126) );
  XOR U3971 ( .A(p_input[1588]), .B(p_input[1572]), .Z(n4127) );
  XNOR U3972 ( .A(n3722), .B(n4122), .Z(n4124) );
  XOR U3973 ( .A(n4128), .B(n4129), .Z(n3722) );
  AND U3974 ( .A(n143), .B(n4130), .Z(n4129) );
  XOR U3975 ( .A(p_input[1556]), .B(p_input[1540]), .Z(n4130) );
  XOR U3976 ( .A(n4131), .B(n4132), .Z(n4122) );
  AND U3977 ( .A(n4133), .B(n4134), .Z(n4132) );
  XOR U3978 ( .A(n4131), .B(n3737), .Z(n4134) );
  XNOR U3979 ( .A(p_input[1571]), .B(n4135), .Z(n3737) );
  AND U3980 ( .A(n146), .B(n4136), .Z(n4135) );
  XOR U3981 ( .A(p_input[1587]), .B(p_input[1571]), .Z(n4136) );
  XNOR U3982 ( .A(n3734), .B(n4131), .Z(n4133) );
  XOR U3983 ( .A(n4137), .B(n4138), .Z(n3734) );
  AND U3984 ( .A(n143), .B(n4139), .Z(n4138) );
  XOR U3985 ( .A(p_input[1555]), .B(p_input[1539]), .Z(n4139) );
  XOR U3986 ( .A(n4140), .B(n4141), .Z(n4131) );
  AND U3987 ( .A(n4142), .B(n4143), .Z(n4141) );
  XOR U3988 ( .A(n3749), .B(n4140), .Z(n4143) );
  XNOR U3989 ( .A(p_input[1570]), .B(n4144), .Z(n3749) );
  AND U3990 ( .A(n146), .B(n4145), .Z(n4144) );
  XOR U3991 ( .A(p_input[1586]), .B(p_input[1570]), .Z(n4145) );
  XNOR U3992 ( .A(n4140), .B(n3746), .Z(n4142) );
  XOR U3993 ( .A(n4146), .B(n4147), .Z(n3746) );
  AND U3994 ( .A(n143), .B(n4148), .Z(n4147) );
  XOR U3995 ( .A(p_input[1554]), .B(p_input[1538]), .Z(n4148) );
  XOR U3996 ( .A(n4149), .B(n4150), .Z(n4140) );
  AND U3997 ( .A(n4151), .B(n4152), .Z(n4150) );
  XNOR U3998 ( .A(n4153), .B(n3762), .Z(n4152) );
  XNOR U3999 ( .A(p_input[1569]), .B(n4154), .Z(n3762) );
  AND U4000 ( .A(n146), .B(n4155), .Z(n4154) );
  XNOR U4001 ( .A(p_input[1585]), .B(n4156), .Z(n4155) );
  IV U4002 ( .A(p_input[1569]), .Z(n4156) );
  XNOR U4003 ( .A(n3759), .B(n4149), .Z(n4151) );
  XNOR U4004 ( .A(p_input[1537]), .B(n4157), .Z(n3759) );
  AND U4005 ( .A(n143), .B(n4158), .Z(n4157) );
  XOR U4006 ( .A(p_input[1553]), .B(p_input[1537]), .Z(n4158) );
  IV U4007 ( .A(n4153), .Z(n4149) );
  AND U4008 ( .A(n4024), .B(n4027), .Z(n4153) );
  XOR U4009 ( .A(p_input[1568]), .B(n4159), .Z(n4027) );
  AND U4010 ( .A(n146), .B(n4160), .Z(n4159) );
  XOR U4011 ( .A(p_input[1584]), .B(p_input[1568]), .Z(n4160) );
  XOR U4012 ( .A(n4161), .B(n4162), .Z(n146) );
  AND U4013 ( .A(n4163), .B(n4164), .Z(n4162) );
  XNOR U4014 ( .A(p_input[1599]), .B(n4161), .Z(n4164) );
  XOR U4015 ( .A(n4161), .B(p_input[1583]), .Z(n4163) );
  XOR U4016 ( .A(n4165), .B(n4166), .Z(n4161) );
  AND U4017 ( .A(n4167), .B(n4168), .Z(n4166) );
  XNOR U4018 ( .A(p_input[1598]), .B(n4165), .Z(n4168) );
  XOR U4019 ( .A(n4165), .B(p_input[1582]), .Z(n4167) );
  XOR U4020 ( .A(n4169), .B(n4170), .Z(n4165) );
  AND U4021 ( .A(n4171), .B(n4172), .Z(n4170) );
  XNOR U4022 ( .A(p_input[1597]), .B(n4169), .Z(n4172) );
  XOR U4023 ( .A(n4169), .B(p_input[1581]), .Z(n4171) );
  XOR U4024 ( .A(n4173), .B(n4174), .Z(n4169) );
  AND U4025 ( .A(n4175), .B(n4176), .Z(n4174) );
  XNOR U4026 ( .A(p_input[1596]), .B(n4173), .Z(n4176) );
  XOR U4027 ( .A(n4173), .B(p_input[1580]), .Z(n4175) );
  XOR U4028 ( .A(n4177), .B(n4178), .Z(n4173) );
  AND U4029 ( .A(n4179), .B(n4180), .Z(n4178) );
  XNOR U4030 ( .A(p_input[1595]), .B(n4177), .Z(n4180) );
  XOR U4031 ( .A(n4177), .B(p_input[1579]), .Z(n4179) );
  XOR U4032 ( .A(n4181), .B(n4182), .Z(n4177) );
  AND U4033 ( .A(n4183), .B(n4184), .Z(n4182) );
  XNOR U4034 ( .A(p_input[1594]), .B(n4181), .Z(n4184) );
  XOR U4035 ( .A(n4181), .B(p_input[1578]), .Z(n4183) );
  XOR U4036 ( .A(n4185), .B(n4186), .Z(n4181) );
  AND U4037 ( .A(n4187), .B(n4188), .Z(n4186) );
  XNOR U4038 ( .A(p_input[1593]), .B(n4185), .Z(n4188) );
  XOR U4039 ( .A(n4185), .B(p_input[1577]), .Z(n4187) );
  XOR U4040 ( .A(n4189), .B(n4190), .Z(n4185) );
  AND U4041 ( .A(n4191), .B(n4192), .Z(n4190) );
  XNOR U4042 ( .A(p_input[1592]), .B(n4189), .Z(n4192) );
  XOR U4043 ( .A(n4189), .B(p_input[1576]), .Z(n4191) );
  XOR U4044 ( .A(n4193), .B(n4194), .Z(n4189) );
  AND U4045 ( .A(n4195), .B(n4196), .Z(n4194) );
  XNOR U4046 ( .A(p_input[1591]), .B(n4193), .Z(n4196) );
  XOR U4047 ( .A(n4193), .B(p_input[1575]), .Z(n4195) );
  XOR U4048 ( .A(n4197), .B(n4198), .Z(n4193) );
  AND U4049 ( .A(n4199), .B(n4200), .Z(n4198) );
  XNOR U4050 ( .A(p_input[1590]), .B(n4197), .Z(n4200) );
  XOR U4051 ( .A(n4197), .B(p_input[1574]), .Z(n4199) );
  XOR U4052 ( .A(n4201), .B(n4202), .Z(n4197) );
  AND U4053 ( .A(n4203), .B(n4204), .Z(n4202) );
  XNOR U4054 ( .A(p_input[1589]), .B(n4201), .Z(n4204) );
  XOR U4055 ( .A(n4201), .B(p_input[1573]), .Z(n4203) );
  XOR U4056 ( .A(n4205), .B(n4206), .Z(n4201) );
  AND U4057 ( .A(n4207), .B(n4208), .Z(n4206) );
  XNOR U4058 ( .A(p_input[1588]), .B(n4205), .Z(n4208) );
  XOR U4059 ( .A(n4205), .B(p_input[1572]), .Z(n4207) );
  XOR U4060 ( .A(n4209), .B(n4210), .Z(n4205) );
  AND U4061 ( .A(n4211), .B(n4212), .Z(n4210) );
  XNOR U4062 ( .A(p_input[1587]), .B(n4209), .Z(n4212) );
  XOR U4063 ( .A(n4209), .B(p_input[1571]), .Z(n4211) );
  XOR U4064 ( .A(n4213), .B(n4214), .Z(n4209) );
  AND U4065 ( .A(n4215), .B(n4216), .Z(n4214) );
  XNOR U4066 ( .A(p_input[1586]), .B(n4213), .Z(n4216) );
  XOR U4067 ( .A(n4213), .B(p_input[1570]), .Z(n4215) );
  XNOR U4068 ( .A(n4217), .B(n4218), .Z(n4213) );
  AND U4069 ( .A(n4219), .B(n4220), .Z(n4218) );
  XOR U4070 ( .A(p_input[1585]), .B(n4217), .Z(n4220) );
  XNOR U4071 ( .A(p_input[1569]), .B(n4217), .Z(n4219) );
  AND U4072 ( .A(p_input[1584]), .B(n4221), .Z(n4217) );
  IV U4073 ( .A(p_input[1568]), .Z(n4221) );
  XNOR U4074 ( .A(p_input[1536]), .B(n4222), .Z(n4024) );
  AND U4075 ( .A(n143), .B(n4223), .Z(n4222) );
  XOR U4076 ( .A(p_input[1552]), .B(p_input[1536]), .Z(n4223) );
  XOR U4077 ( .A(n4224), .B(n4225), .Z(n143) );
  AND U4078 ( .A(n4226), .B(n4227), .Z(n4225) );
  XNOR U4079 ( .A(p_input[1567]), .B(n4224), .Z(n4227) );
  XOR U4080 ( .A(n4224), .B(p_input[1551]), .Z(n4226) );
  XOR U4081 ( .A(n4228), .B(n4229), .Z(n4224) );
  AND U4082 ( .A(n4230), .B(n4231), .Z(n4229) );
  XNOR U4083 ( .A(p_input[1566]), .B(n4228), .Z(n4231) );
  XNOR U4084 ( .A(n4228), .B(n4038), .Z(n4230) );
  IV U4085 ( .A(p_input[1550]), .Z(n4038) );
  XOR U4086 ( .A(n4232), .B(n4233), .Z(n4228) );
  AND U4087 ( .A(n4234), .B(n4235), .Z(n4233) );
  XNOR U4088 ( .A(p_input[1565]), .B(n4232), .Z(n4235) );
  XNOR U4089 ( .A(n4232), .B(n4047), .Z(n4234) );
  IV U4090 ( .A(p_input[1549]), .Z(n4047) );
  XOR U4091 ( .A(n4236), .B(n4237), .Z(n4232) );
  AND U4092 ( .A(n4238), .B(n4239), .Z(n4237) );
  XNOR U4093 ( .A(p_input[1564]), .B(n4236), .Z(n4239) );
  XNOR U4094 ( .A(n4236), .B(n4056), .Z(n4238) );
  IV U4095 ( .A(p_input[1548]), .Z(n4056) );
  XOR U4096 ( .A(n4240), .B(n4241), .Z(n4236) );
  AND U4097 ( .A(n4242), .B(n4243), .Z(n4241) );
  XNOR U4098 ( .A(p_input[1563]), .B(n4240), .Z(n4243) );
  XNOR U4099 ( .A(n4240), .B(n4065), .Z(n4242) );
  IV U4100 ( .A(p_input[1547]), .Z(n4065) );
  XOR U4101 ( .A(n4244), .B(n4245), .Z(n4240) );
  AND U4102 ( .A(n4246), .B(n4247), .Z(n4245) );
  XNOR U4103 ( .A(p_input[1562]), .B(n4244), .Z(n4247) );
  XNOR U4104 ( .A(n4244), .B(n4074), .Z(n4246) );
  IV U4105 ( .A(p_input[1546]), .Z(n4074) );
  XOR U4106 ( .A(n4248), .B(n4249), .Z(n4244) );
  AND U4107 ( .A(n4250), .B(n4251), .Z(n4249) );
  XNOR U4108 ( .A(p_input[1561]), .B(n4248), .Z(n4251) );
  XNOR U4109 ( .A(n4248), .B(n4083), .Z(n4250) );
  IV U4110 ( .A(p_input[1545]), .Z(n4083) );
  XOR U4111 ( .A(n4252), .B(n4253), .Z(n4248) );
  AND U4112 ( .A(n4254), .B(n4255), .Z(n4253) );
  XNOR U4113 ( .A(p_input[1560]), .B(n4252), .Z(n4255) );
  XNOR U4114 ( .A(n4252), .B(n4092), .Z(n4254) );
  IV U4115 ( .A(p_input[1544]), .Z(n4092) );
  XOR U4116 ( .A(n4256), .B(n4257), .Z(n4252) );
  AND U4117 ( .A(n4258), .B(n4259), .Z(n4257) );
  XNOR U4118 ( .A(p_input[1559]), .B(n4256), .Z(n4259) );
  XNOR U4119 ( .A(n4256), .B(n4101), .Z(n4258) );
  IV U4120 ( .A(p_input[1543]), .Z(n4101) );
  XOR U4121 ( .A(n4260), .B(n4261), .Z(n4256) );
  AND U4122 ( .A(n4262), .B(n4263), .Z(n4261) );
  XNOR U4123 ( .A(p_input[1558]), .B(n4260), .Z(n4263) );
  XNOR U4124 ( .A(n4260), .B(n4110), .Z(n4262) );
  IV U4125 ( .A(p_input[1542]), .Z(n4110) );
  XOR U4126 ( .A(n4264), .B(n4265), .Z(n4260) );
  AND U4127 ( .A(n4266), .B(n4267), .Z(n4265) );
  XNOR U4128 ( .A(p_input[1557]), .B(n4264), .Z(n4267) );
  XNOR U4129 ( .A(n4264), .B(n4119), .Z(n4266) );
  IV U4130 ( .A(p_input[1541]), .Z(n4119) );
  XOR U4131 ( .A(n4268), .B(n4269), .Z(n4264) );
  AND U4132 ( .A(n4270), .B(n4271), .Z(n4269) );
  XNOR U4133 ( .A(p_input[1556]), .B(n4268), .Z(n4271) );
  XNOR U4134 ( .A(n4268), .B(n4128), .Z(n4270) );
  IV U4135 ( .A(p_input[1540]), .Z(n4128) );
  XOR U4136 ( .A(n4272), .B(n4273), .Z(n4268) );
  AND U4137 ( .A(n4274), .B(n4275), .Z(n4273) );
  XNOR U4138 ( .A(p_input[1555]), .B(n4272), .Z(n4275) );
  XNOR U4139 ( .A(n4272), .B(n4137), .Z(n4274) );
  IV U4140 ( .A(p_input[1539]), .Z(n4137) );
  XOR U4141 ( .A(n4276), .B(n4277), .Z(n4272) );
  AND U4142 ( .A(n4278), .B(n4279), .Z(n4277) );
  XNOR U4143 ( .A(p_input[1554]), .B(n4276), .Z(n4279) );
  XNOR U4144 ( .A(n4276), .B(n4146), .Z(n4278) );
  IV U4145 ( .A(p_input[1538]), .Z(n4146) );
  XNOR U4146 ( .A(n4280), .B(n4281), .Z(n4276) );
  AND U4147 ( .A(n4282), .B(n4283), .Z(n4281) );
  XOR U4148 ( .A(p_input[1553]), .B(n4280), .Z(n4283) );
  XNOR U4149 ( .A(p_input[1537]), .B(n4280), .Z(n4282) );
  AND U4150 ( .A(p_input[1552]), .B(n4284), .Z(n4280) );
  IV U4151 ( .A(p_input[1536]), .Z(n4284) );
  XOR U4152 ( .A(n4285), .B(n4286), .Z(n739) );
  AND U4153 ( .A(n536), .B(n4287), .Z(n4286) );
  XNOR U4154 ( .A(n4288), .B(n4285), .Z(n4287) );
  XOR U4155 ( .A(n4289), .B(n4290), .Z(n536) );
  AND U4156 ( .A(n4291), .B(n4292), .Z(n4290) );
  XOR U4157 ( .A(n4289), .B(n754), .Z(n4292) );
  XNOR U4158 ( .A(n4293), .B(n4294), .Z(n754) );
  AND U4159 ( .A(n4295), .B(n502), .Z(n4294) );
  AND U4160 ( .A(n4293), .B(n4296), .Z(n4295) );
  XNOR U4161 ( .A(n751), .B(n4289), .Z(n4291) );
  XOR U4162 ( .A(n4297), .B(n4298), .Z(n751) );
  AND U4163 ( .A(n4299), .B(n499), .Z(n4298) );
  NOR U4164 ( .A(n4297), .B(n4300), .Z(n4299) );
  XOR U4165 ( .A(n4301), .B(n4302), .Z(n4289) );
  AND U4166 ( .A(n4303), .B(n4304), .Z(n4302) );
  XOR U4167 ( .A(n4301), .B(n766), .Z(n4304) );
  XOR U4168 ( .A(n4305), .B(n4306), .Z(n766) );
  AND U4169 ( .A(n502), .B(n4307), .Z(n4306) );
  XOR U4170 ( .A(n4308), .B(n4305), .Z(n4307) );
  XNOR U4171 ( .A(n763), .B(n4301), .Z(n4303) );
  XOR U4172 ( .A(n4309), .B(n4310), .Z(n763) );
  AND U4173 ( .A(n499), .B(n4311), .Z(n4310) );
  XOR U4174 ( .A(n4312), .B(n4309), .Z(n4311) );
  XOR U4175 ( .A(n4313), .B(n4314), .Z(n4301) );
  AND U4176 ( .A(n4315), .B(n4316), .Z(n4314) );
  XOR U4177 ( .A(n4313), .B(n778), .Z(n4316) );
  XOR U4178 ( .A(n4317), .B(n4318), .Z(n778) );
  AND U4179 ( .A(n502), .B(n4319), .Z(n4318) );
  XOR U4180 ( .A(n4320), .B(n4317), .Z(n4319) );
  XNOR U4181 ( .A(n775), .B(n4313), .Z(n4315) );
  XOR U4182 ( .A(n4321), .B(n4322), .Z(n775) );
  AND U4183 ( .A(n499), .B(n4323), .Z(n4322) );
  XOR U4184 ( .A(n4324), .B(n4321), .Z(n4323) );
  XOR U4185 ( .A(n4325), .B(n4326), .Z(n4313) );
  AND U4186 ( .A(n4327), .B(n4328), .Z(n4326) );
  XOR U4187 ( .A(n4325), .B(n790), .Z(n4328) );
  XOR U4188 ( .A(n4329), .B(n4330), .Z(n790) );
  AND U4189 ( .A(n502), .B(n4331), .Z(n4330) );
  XOR U4190 ( .A(n4332), .B(n4329), .Z(n4331) );
  XNOR U4191 ( .A(n787), .B(n4325), .Z(n4327) );
  XOR U4192 ( .A(n4333), .B(n4334), .Z(n787) );
  AND U4193 ( .A(n499), .B(n4335), .Z(n4334) );
  XOR U4194 ( .A(n4336), .B(n4333), .Z(n4335) );
  XOR U4195 ( .A(n4337), .B(n4338), .Z(n4325) );
  AND U4196 ( .A(n4339), .B(n4340), .Z(n4338) );
  XOR U4197 ( .A(n4337), .B(n802), .Z(n4340) );
  XOR U4198 ( .A(n4341), .B(n4342), .Z(n802) );
  AND U4199 ( .A(n502), .B(n4343), .Z(n4342) );
  XOR U4200 ( .A(n4344), .B(n4341), .Z(n4343) );
  XNOR U4201 ( .A(n799), .B(n4337), .Z(n4339) );
  XOR U4202 ( .A(n4345), .B(n4346), .Z(n799) );
  AND U4203 ( .A(n499), .B(n4347), .Z(n4346) );
  XOR U4204 ( .A(n4348), .B(n4345), .Z(n4347) );
  XOR U4205 ( .A(n4349), .B(n4350), .Z(n4337) );
  AND U4206 ( .A(n4351), .B(n4352), .Z(n4350) );
  XOR U4207 ( .A(n4349), .B(n814), .Z(n4352) );
  XOR U4208 ( .A(n4353), .B(n4354), .Z(n814) );
  AND U4209 ( .A(n502), .B(n4355), .Z(n4354) );
  XOR U4210 ( .A(n4356), .B(n4353), .Z(n4355) );
  XNOR U4211 ( .A(n811), .B(n4349), .Z(n4351) );
  XOR U4212 ( .A(n4357), .B(n4358), .Z(n811) );
  AND U4213 ( .A(n499), .B(n4359), .Z(n4358) );
  XOR U4214 ( .A(n4360), .B(n4357), .Z(n4359) );
  XOR U4215 ( .A(n4361), .B(n4362), .Z(n4349) );
  AND U4216 ( .A(n4363), .B(n4364), .Z(n4362) );
  XOR U4217 ( .A(n4361), .B(n826), .Z(n4364) );
  XOR U4218 ( .A(n4365), .B(n4366), .Z(n826) );
  AND U4219 ( .A(n502), .B(n4367), .Z(n4366) );
  XOR U4220 ( .A(n4368), .B(n4365), .Z(n4367) );
  XNOR U4221 ( .A(n823), .B(n4361), .Z(n4363) );
  XOR U4222 ( .A(n4369), .B(n4370), .Z(n823) );
  AND U4223 ( .A(n499), .B(n4371), .Z(n4370) );
  XOR U4224 ( .A(n4372), .B(n4369), .Z(n4371) );
  XOR U4225 ( .A(n4373), .B(n4374), .Z(n4361) );
  AND U4226 ( .A(n4375), .B(n4376), .Z(n4374) );
  XOR U4227 ( .A(n4373), .B(n838), .Z(n4376) );
  XOR U4228 ( .A(n4377), .B(n4378), .Z(n838) );
  AND U4229 ( .A(n502), .B(n4379), .Z(n4378) );
  XOR U4230 ( .A(n4380), .B(n4377), .Z(n4379) );
  XNOR U4231 ( .A(n835), .B(n4373), .Z(n4375) );
  XOR U4232 ( .A(n4381), .B(n4382), .Z(n835) );
  AND U4233 ( .A(n499), .B(n4383), .Z(n4382) );
  XOR U4234 ( .A(n4384), .B(n4381), .Z(n4383) );
  XOR U4235 ( .A(n4385), .B(n4386), .Z(n4373) );
  AND U4236 ( .A(n4387), .B(n4388), .Z(n4386) );
  XOR U4237 ( .A(n4385), .B(n850), .Z(n4388) );
  XOR U4238 ( .A(n4389), .B(n4390), .Z(n850) );
  AND U4239 ( .A(n502), .B(n4391), .Z(n4390) );
  XOR U4240 ( .A(n4392), .B(n4389), .Z(n4391) );
  XNOR U4241 ( .A(n847), .B(n4385), .Z(n4387) );
  XOR U4242 ( .A(n4393), .B(n4394), .Z(n847) );
  AND U4243 ( .A(n499), .B(n4395), .Z(n4394) );
  XOR U4244 ( .A(n4396), .B(n4393), .Z(n4395) );
  XOR U4245 ( .A(n4397), .B(n4398), .Z(n4385) );
  AND U4246 ( .A(n4399), .B(n4400), .Z(n4398) );
  XOR U4247 ( .A(n4397), .B(n862), .Z(n4400) );
  XOR U4248 ( .A(n4401), .B(n4402), .Z(n862) );
  AND U4249 ( .A(n502), .B(n4403), .Z(n4402) );
  XOR U4250 ( .A(n4404), .B(n4401), .Z(n4403) );
  XNOR U4251 ( .A(n859), .B(n4397), .Z(n4399) );
  XOR U4252 ( .A(n4405), .B(n4406), .Z(n859) );
  AND U4253 ( .A(n499), .B(n4407), .Z(n4406) );
  XOR U4254 ( .A(n4408), .B(n4405), .Z(n4407) );
  XOR U4255 ( .A(n4409), .B(n4410), .Z(n4397) );
  AND U4256 ( .A(n4411), .B(n4412), .Z(n4410) );
  XOR U4257 ( .A(n4409), .B(n874), .Z(n4412) );
  XOR U4258 ( .A(n4413), .B(n4414), .Z(n874) );
  AND U4259 ( .A(n502), .B(n4415), .Z(n4414) );
  XOR U4260 ( .A(n4416), .B(n4413), .Z(n4415) );
  XNOR U4261 ( .A(n871), .B(n4409), .Z(n4411) );
  XOR U4262 ( .A(n4417), .B(n4418), .Z(n871) );
  AND U4263 ( .A(n499), .B(n4419), .Z(n4418) );
  XOR U4264 ( .A(n4420), .B(n4417), .Z(n4419) );
  XOR U4265 ( .A(n4421), .B(n4422), .Z(n4409) );
  AND U4266 ( .A(n4423), .B(n4424), .Z(n4422) );
  XOR U4267 ( .A(n4421), .B(n886), .Z(n4424) );
  XOR U4268 ( .A(n4425), .B(n4426), .Z(n886) );
  AND U4269 ( .A(n502), .B(n4427), .Z(n4426) );
  XOR U4270 ( .A(n4428), .B(n4425), .Z(n4427) );
  XNOR U4271 ( .A(n883), .B(n4421), .Z(n4423) );
  XOR U4272 ( .A(n4429), .B(n4430), .Z(n883) );
  AND U4273 ( .A(n499), .B(n4431), .Z(n4430) );
  XOR U4274 ( .A(n4432), .B(n4429), .Z(n4431) );
  XOR U4275 ( .A(n4433), .B(n4434), .Z(n4421) );
  AND U4276 ( .A(n4435), .B(n4436), .Z(n4434) );
  XOR U4277 ( .A(n4433), .B(n898), .Z(n4436) );
  XOR U4278 ( .A(n4437), .B(n4438), .Z(n898) );
  AND U4279 ( .A(n502), .B(n4439), .Z(n4438) );
  XOR U4280 ( .A(n4440), .B(n4437), .Z(n4439) );
  XNOR U4281 ( .A(n895), .B(n4433), .Z(n4435) );
  XOR U4282 ( .A(n4441), .B(n4442), .Z(n895) );
  AND U4283 ( .A(n499), .B(n4443), .Z(n4442) );
  XOR U4284 ( .A(n4444), .B(n4441), .Z(n4443) );
  XOR U4285 ( .A(n4445), .B(n4446), .Z(n4433) );
  AND U4286 ( .A(n4447), .B(n4448), .Z(n4446) );
  XOR U4287 ( .A(n910), .B(n4445), .Z(n4448) );
  XOR U4288 ( .A(n4449), .B(n4450), .Z(n910) );
  AND U4289 ( .A(n502), .B(n4451), .Z(n4450) );
  XOR U4290 ( .A(n4449), .B(n4452), .Z(n4451) );
  XNOR U4291 ( .A(n4445), .B(n907), .Z(n4447) );
  XOR U4292 ( .A(n4453), .B(n4454), .Z(n907) );
  AND U4293 ( .A(n499), .B(n4455), .Z(n4454) );
  XOR U4294 ( .A(n4453), .B(n4456), .Z(n4455) );
  XOR U4295 ( .A(n4457), .B(n4458), .Z(n4445) );
  AND U4296 ( .A(n4459), .B(n4460), .Z(n4458) );
  XNOR U4297 ( .A(n4461), .B(n923), .Z(n4460) );
  XOR U4298 ( .A(n4462), .B(n4463), .Z(n923) );
  AND U4299 ( .A(n502), .B(n4464), .Z(n4463) );
  XOR U4300 ( .A(n4465), .B(n4462), .Z(n4464) );
  XNOR U4301 ( .A(n920), .B(n4457), .Z(n4459) );
  XOR U4302 ( .A(n4466), .B(n4467), .Z(n920) );
  AND U4303 ( .A(n499), .B(n4468), .Z(n4467) );
  XOR U4304 ( .A(n4469), .B(n4466), .Z(n4468) );
  IV U4305 ( .A(n4461), .Z(n4457) );
  AND U4306 ( .A(n4285), .B(n4288), .Z(n4461) );
  XNOR U4307 ( .A(n4470), .B(n4471), .Z(n4288) );
  AND U4308 ( .A(n502), .B(n4472), .Z(n4471) );
  XNOR U4309 ( .A(n4473), .B(n4470), .Z(n4472) );
  XOR U4310 ( .A(n4474), .B(n4475), .Z(n502) );
  AND U4311 ( .A(n4476), .B(n4477), .Z(n4475) );
  XOR U4312 ( .A(n4296), .B(n4474), .Z(n4477) );
  IV U4313 ( .A(n4478), .Z(n4296) );
  AND U4314 ( .A(n4479), .B(n4480), .Z(n4478) );
  XOR U4315 ( .A(n4474), .B(n4293), .Z(n4476) );
  AND U4316 ( .A(n4481), .B(n4482), .Z(n4293) );
  XOR U4317 ( .A(n4483), .B(n4484), .Z(n4474) );
  AND U4318 ( .A(n4485), .B(n4486), .Z(n4484) );
  XOR U4319 ( .A(n4483), .B(n4308), .Z(n4486) );
  XOR U4320 ( .A(n4487), .B(n4488), .Z(n4308) );
  AND U4321 ( .A(n422), .B(n4489), .Z(n4488) );
  XOR U4322 ( .A(n4490), .B(n4487), .Z(n4489) );
  XNOR U4323 ( .A(n4305), .B(n4483), .Z(n4485) );
  XOR U4324 ( .A(n4491), .B(n4492), .Z(n4305) );
  AND U4325 ( .A(n420), .B(n4493), .Z(n4492) );
  XOR U4326 ( .A(n4494), .B(n4491), .Z(n4493) );
  XOR U4327 ( .A(n4495), .B(n4496), .Z(n4483) );
  AND U4328 ( .A(n4497), .B(n4498), .Z(n4496) );
  XOR U4329 ( .A(n4495), .B(n4320), .Z(n4498) );
  XOR U4330 ( .A(n4499), .B(n4500), .Z(n4320) );
  AND U4331 ( .A(n422), .B(n4501), .Z(n4500) );
  XOR U4332 ( .A(n4502), .B(n4499), .Z(n4501) );
  XNOR U4333 ( .A(n4317), .B(n4495), .Z(n4497) );
  XOR U4334 ( .A(n4503), .B(n4504), .Z(n4317) );
  AND U4335 ( .A(n420), .B(n4505), .Z(n4504) );
  XOR U4336 ( .A(n4506), .B(n4503), .Z(n4505) );
  XOR U4337 ( .A(n4507), .B(n4508), .Z(n4495) );
  AND U4338 ( .A(n4509), .B(n4510), .Z(n4508) );
  XOR U4339 ( .A(n4507), .B(n4332), .Z(n4510) );
  XOR U4340 ( .A(n4511), .B(n4512), .Z(n4332) );
  AND U4341 ( .A(n422), .B(n4513), .Z(n4512) );
  XOR U4342 ( .A(n4514), .B(n4511), .Z(n4513) );
  XNOR U4343 ( .A(n4329), .B(n4507), .Z(n4509) );
  XOR U4344 ( .A(n4515), .B(n4516), .Z(n4329) );
  AND U4345 ( .A(n420), .B(n4517), .Z(n4516) );
  XOR U4346 ( .A(n4518), .B(n4515), .Z(n4517) );
  XOR U4347 ( .A(n4519), .B(n4520), .Z(n4507) );
  AND U4348 ( .A(n4521), .B(n4522), .Z(n4520) );
  XOR U4349 ( .A(n4519), .B(n4344), .Z(n4522) );
  XOR U4350 ( .A(n4523), .B(n4524), .Z(n4344) );
  AND U4351 ( .A(n422), .B(n4525), .Z(n4524) );
  XOR U4352 ( .A(n4526), .B(n4523), .Z(n4525) );
  XNOR U4353 ( .A(n4341), .B(n4519), .Z(n4521) );
  XOR U4354 ( .A(n4527), .B(n4528), .Z(n4341) );
  AND U4355 ( .A(n420), .B(n4529), .Z(n4528) );
  XOR U4356 ( .A(n4530), .B(n4527), .Z(n4529) );
  XOR U4357 ( .A(n4531), .B(n4532), .Z(n4519) );
  AND U4358 ( .A(n4533), .B(n4534), .Z(n4532) );
  XOR U4359 ( .A(n4531), .B(n4356), .Z(n4534) );
  XOR U4360 ( .A(n4535), .B(n4536), .Z(n4356) );
  AND U4361 ( .A(n422), .B(n4537), .Z(n4536) );
  XOR U4362 ( .A(n4538), .B(n4535), .Z(n4537) );
  XNOR U4363 ( .A(n4353), .B(n4531), .Z(n4533) );
  XOR U4364 ( .A(n4539), .B(n4540), .Z(n4353) );
  AND U4365 ( .A(n420), .B(n4541), .Z(n4540) );
  XOR U4366 ( .A(n4542), .B(n4539), .Z(n4541) );
  XOR U4367 ( .A(n4543), .B(n4544), .Z(n4531) );
  AND U4368 ( .A(n4545), .B(n4546), .Z(n4544) );
  XOR U4369 ( .A(n4543), .B(n4368), .Z(n4546) );
  XOR U4370 ( .A(n4547), .B(n4548), .Z(n4368) );
  AND U4371 ( .A(n422), .B(n4549), .Z(n4548) );
  XOR U4372 ( .A(n4550), .B(n4547), .Z(n4549) );
  XNOR U4373 ( .A(n4365), .B(n4543), .Z(n4545) );
  XOR U4374 ( .A(n4551), .B(n4552), .Z(n4365) );
  AND U4375 ( .A(n420), .B(n4553), .Z(n4552) );
  XOR U4376 ( .A(n4554), .B(n4551), .Z(n4553) );
  XOR U4377 ( .A(n4555), .B(n4556), .Z(n4543) );
  AND U4378 ( .A(n4557), .B(n4558), .Z(n4556) );
  XOR U4379 ( .A(n4555), .B(n4380), .Z(n4558) );
  XOR U4380 ( .A(n4559), .B(n4560), .Z(n4380) );
  AND U4381 ( .A(n422), .B(n4561), .Z(n4560) );
  XOR U4382 ( .A(n4562), .B(n4559), .Z(n4561) );
  XNOR U4383 ( .A(n4377), .B(n4555), .Z(n4557) );
  XOR U4384 ( .A(n4563), .B(n4564), .Z(n4377) );
  AND U4385 ( .A(n420), .B(n4565), .Z(n4564) );
  XOR U4386 ( .A(n4566), .B(n4563), .Z(n4565) );
  XOR U4387 ( .A(n4567), .B(n4568), .Z(n4555) );
  AND U4388 ( .A(n4569), .B(n4570), .Z(n4568) );
  XOR U4389 ( .A(n4567), .B(n4392), .Z(n4570) );
  XOR U4390 ( .A(n4571), .B(n4572), .Z(n4392) );
  AND U4391 ( .A(n422), .B(n4573), .Z(n4572) );
  XOR U4392 ( .A(n4574), .B(n4571), .Z(n4573) );
  XNOR U4393 ( .A(n4389), .B(n4567), .Z(n4569) );
  XOR U4394 ( .A(n4575), .B(n4576), .Z(n4389) );
  AND U4395 ( .A(n420), .B(n4577), .Z(n4576) );
  XOR U4396 ( .A(n4578), .B(n4575), .Z(n4577) );
  XOR U4397 ( .A(n4579), .B(n4580), .Z(n4567) );
  AND U4398 ( .A(n4581), .B(n4582), .Z(n4580) );
  XOR U4399 ( .A(n4579), .B(n4404), .Z(n4582) );
  XOR U4400 ( .A(n4583), .B(n4584), .Z(n4404) );
  AND U4401 ( .A(n422), .B(n4585), .Z(n4584) );
  XOR U4402 ( .A(n4586), .B(n4583), .Z(n4585) );
  XNOR U4403 ( .A(n4401), .B(n4579), .Z(n4581) );
  XOR U4404 ( .A(n4587), .B(n4588), .Z(n4401) );
  AND U4405 ( .A(n420), .B(n4589), .Z(n4588) );
  XOR U4406 ( .A(n4590), .B(n4587), .Z(n4589) );
  XOR U4407 ( .A(n4591), .B(n4592), .Z(n4579) );
  AND U4408 ( .A(n4593), .B(n4594), .Z(n4592) );
  XOR U4409 ( .A(n4591), .B(n4416), .Z(n4594) );
  XOR U4410 ( .A(n4595), .B(n4596), .Z(n4416) );
  AND U4411 ( .A(n422), .B(n4597), .Z(n4596) );
  XOR U4412 ( .A(n4598), .B(n4595), .Z(n4597) );
  XNOR U4413 ( .A(n4413), .B(n4591), .Z(n4593) );
  XOR U4414 ( .A(n4599), .B(n4600), .Z(n4413) );
  AND U4415 ( .A(n420), .B(n4601), .Z(n4600) );
  XOR U4416 ( .A(n4602), .B(n4599), .Z(n4601) );
  XOR U4417 ( .A(n4603), .B(n4604), .Z(n4591) );
  AND U4418 ( .A(n4605), .B(n4606), .Z(n4604) );
  XOR U4419 ( .A(n4603), .B(n4428), .Z(n4606) );
  XOR U4420 ( .A(n4607), .B(n4608), .Z(n4428) );
  AND U4421 ( .A(n422), .B(n4609), .Z(n4608) );
  XOR U4422 ( .A(n4610), .B(n4607), .Z(n4609) );
  XNOR U4423 ( .A(n4425), .B(n4603), .Z(n4605) );
  XOR U4424 ( .A(n4611), .B(n4612), .Z(n4425) );
  AND U4425 ( .A(n420), .B(n4613), .Z(n4612) );
  XOR U4426 ( .A(n4614), .B(n4611), .Z(n4613) );
  XOR U4427 ( .A(n4615), .B(n4616), .Z(n4603) );
  AND U4428 ( .A(n4617), .B(n4618), .Z(n4616) );
  XOR U4429 ( .A(n4615), .B(n4440), .Z(n4618) );
  XOR U4430 ( .A(n4619), .B(n4620), .Z(n4440) );
  AND U4431 ( .A(n422), .B(n4621), .Z(n4620) );
  XOR U4432 ( .A(n4622), .B(n4619), .Z(n4621) );
  XNOR U4433 ( .A(n4437), .B(n4615), .Z(n4617) );
  XOR U4434 ( .A(n4623), .B(n4624), .Z(n4437) );
  AND U4435 ( .A(n420), .B(n4625), .Z(n4624) );
  XOR U4436 ( .A(n4626), .B(n4623), .Z(n4625) );
  XOR U4437 ( .A(n4627), .B(n4628), .Z(n4615) );
  AND U4438 ( .A(n4629), .B(n4630), .Z(n4628) );
  XOR U4439 ( .A(n4452), .B(n4627), .Z(n4630) );
  XOR U4440 ( .A(n4631), .B(n4632), .Z(n4452) );
  AND U4441 ( .A(n422), .B(n4633), .Z(n4632) );
  XOR U4442 ( .A(n4631), .B(n4634), .Z(n4633) );
  XNOR U4443 ( .A(n4627), .B(n4449), .Z(n4629) );
  XOR U4444 ( .A(n4635), .B(n4636), .Z(n4449) );
  AND U4445 ( .A(n420), .B(n4637), .Z(n4636) );
  XOR U4446 ( .A(n4635), .B(n4638), .Z(n4637) );
  XOR U4447 ( .A(n4639), .B(n4640), .Z(n4627) );
  AND U4448 ( .A(n4641), .B(n4642), .Z(n4640) );
  XNOR U4449 ( .A(n4643), .B(n4465), .Z(n4642) );
  XOR U4450 ( .A(n4644), .B(n4645), .Z(n4465) );
  AND U4451 ( .A(n422), .B(n4646), .Z(n4645) );
  XOR U4452 ( .A(n4647), .B(n4644), .Z(n4646) );
  XNOR U4453 ( .A(n4462), .B(n4639), .Z(n4641) );
  XOR U4454 ( .A(n4648), .B(n4649), .Z(n4462) );
  AND U4455 ( .A(n420), .B(n4650), .Z(n4649) );
  XOR U4456 ( .A(n4651), .B(n4648), .Z(n4650) );
  IV U4457 ( .A(n4643), .Z(n4639) );
  AND U4458 ( .A(n4470), .B(n4473), .Z(n4643) );
  XNOR U4459 ( .A(n4652), .B(n4653), .Z(n4473) );
  AND U4460 ( .A(n422), .B(n4654), .Z(n4653) );
  XNOR U4461 ( .A(n4655), .B(n4652), .Z(n4654) );
  XOR U4462 ( .A(n4656), .B(n4657), .Z(n422) );
  AND U4463 ( .A(n4658), .B(n4659), .Z(n4657) );
  XNOR U4464 ( .A(n4479), .B(n4656), .Z(n4659) );
  AND U4465 ( .A(n4660), .B(n4661), .Z(n4479) );
  XOR U4466 ( .A(n4656), .B(n4480), .Z(n4658) );
  AND U4467 ( .A(n4662), .B(n4663), .Z(n4480) );
  XOR U4468 ( .A(n4664), .B(n4665), .Z(n4656) );
  AND U4469 ( .A(n4666), .B(n4667), .Z(n4665) );
  XOR U4470 ( .A(n4664), .B(n4490), .Z(n4667) );
  XOR U4471 ( .A(n4668), .B(n4669), .Z(n4490) );
  AND U4472 ( .A(n254), .B(n4670), .Z(n4669) );
  XOR U4473 ( .A(n4671), .B(n4668), .Z(n4670) );
  XNOR U4474 ( .A(n4487), .B(n4664), .Z(n4666) );
  XOR U4475 ( .A(n4672), .B(n4673), .Z(n4487) );
  AND U4476 ( .A(n252), .B(n4674), .Z(n4673) );
  XOR U4477 ( .A(n4675), .B(n4672), .Z(n4674) );
  XOR U4478 ( .A(n4676), .B(n4677), .Z(n4664) );
  AND U4479 ( .A(n4678), .B(n4679), .Z(n4677) );
  XOR U4480 ( .A(n4676), .B(n4502), .Z(n4679) );
  XOR U4481 ( .A(n4680), .B(n4681), .Z(n4502) );
  AND U4482 ( .A(n254), .B(n4682), .Z(n4681) );
  XOR U4483 ( .A(n4683), .B(n4680), .Z(n4682) );
  XNOR U4484 ( .A(n4499), .B(n4676), .Z(n4678) );
  XOR U4485 ( .A(n4684), .B(n4685), .Z(n4499) );
  AND U4486 ( .A(n252), .B(n4686), .Z(n4685) );
  XOR U4487 ( .A(n4687), .B(n4684), .Z(n4686) );
  XOR U4488 ( .A(n4688), .B(n4689), .Z(n4676) );
  AND U4489 ( .A(n4690), .B(n4691), .Z(n4689) );
  XOR U4490 ( .A(n4688), .B(n4514), .Z(n4691) );
  XOR U4491 ( .A(n4692), .B(n4693), .Z(n4514) );
  AND U4492 ( .A(n254), .B(n4694), .Z(n4693) );
  XOR U4493 ( .A(n4695), .B(n4692), .Z(n4694) );
  XNOR U4494 ( .A(n4511), .B(n4688), .Z(n4690) );
  XOR U4495 ( .A(n4696), .B(n4697), .Z(n4511) );
  AND U4496 ( .A(n252), .B(n4698), .Z(n4697) );
  XOR U4497 ( .A(n4699), .B(n4696), .Z(n4698) );
  XOR U4498 ( .A(n4700), .B(n4701), .Z(n4688) );
  AND U4499 ( .A(n4702), .B(n4703), .Z(n4701) );
  XOR U4500 ( .A(n4700), .B(n4526), .Z(n4703) );
  XOR U4501 ( .A(n4704), .B(n4705), .Z(n4526) );
  AND U4502 ( .A(n254), .B(n4706), .Z(n4705) );
  XOR U4503 ( .A(n4707), .B(n4704), .Z(n4706) );
  XNOR U4504 ( .A(n4523), .B(n4700), .Z(n4702) );
  XOR U4505 ( .A(n4708), .B(n4709), .Z(n4523) );
  AND U4506 ( .A(n252), .B(n4710), .Z(n4709) );
  XOR U4507 ( .A(n4711), .B(n4708), .Z(n4710) );
  XOR U4508 ( .A(n4712), .B(n4713), .Z(n4700) );
  AND U4509 ( .A(n4714), .B(n4715), .Z(n4713) );
  XOR U4510 ( .A(n4712), .B(n4538), .Z(n4715) );
  XOR U4511 ( .A(n4716), .B(n4717), .Z(n4538) );
  AND U4512 ( .A(n254), .B(n4718), .Z(n4717) );
  XOR U4513 ( .A(n4719), .B(n4716), .Z(n4718) );
  XNOR U4514 ( .A(n4535), .B(n4712), .Z(n4714) );
  XOR U4515 ( .A(n4720), .B(n4721), .Z(n4535) );
  AND U4516 ( .A(n252), .B(n4722), .Z(n4721) );
  XOR U4517 ( .A(n4723), .B(n4720), .Z(n4722) );
  XOR U4518 ( .A(n4724), .B(n4725), .Z(n4712) );
  AND U4519 ( .A(n4726), .B(n4727), .Z(n4725) );
  XOR U4520 ( .A(n4724), .B(n4550), .Z(n4727) );
  XOR U4521 ( .A(n4728), .B(n4729), .Z(n4550) );
  AND U4522 ( .A(n254), .B(n4730), .Z(n4729) );
  XOR U4523 ( .A(n4731), .B(n4728), .Z(n4730) );
  XNOR U4524 ( .A(n4547), .B(n4724), .Z(n4726) );
  XOR U4525 ( .A(n4732), .B(n4733), .Z(n4547) );
  AND U4526 ( .A(n252), .B(n4734), .Z(n4733) );
  XOR U4527 ( .A(n4735), .B(n4732), .Z(n4734) );
  XOR U4528 ( .A(n4736), .B(n4737), .Z(n4724) );
  AND U4529 ( .A(n4738), .B(n4739), .Z(n4737) );
  XOR U4530 ( .A(n4736), .B(n4562), .Z(n4739) );
  XOR U4531 ( .A(n4740), .B(n4741), .Z(n4562) );
  AND U4532 ( .A(n254), .B(n4742), .Z(n4741) );
  XOR U4533 ( .A(n4743), .B(n4740), .Z(n4742) );
  XNOR U4534 ( .A(n4559), .B(n4736), .Z(n4738) );
  XOR U4535 ( .A(n4744), .B(n4745), .Z(n4559) );
  AND U4536 ( .A(n252), .B(n4746), .Z(n4745) );
  XOR U4537 ( .A(n4747), .B(n4744), .Z(n4746) );
  XOR U4538 ( .A(n4748), .B(n4749), .Z(n4736) );
  AND U4539 ( .A(n4750), .B(n4751), .Z(n4749) );
  XOR U4540 ( .A(n4748), .B(n4574), .Z(n4751) );
  XOR U4541 ( .A(n4752), .B(n4753), .Z(n4574) );
  AND U4542 ( .A(n254), .B(n4754), .Z(n4753) );
  XOR U4543 ( .A(n4755), .B(n4752), .Z(n4754) );
  XNOR U4544 ( .A(n4571), .B(n4748), .Z(n4750) );
  XOR U4545 ( .A(n4756), .B(n4757), .Z(n4571) );
  AND U4546 ( .A(n252), .B(n4758), .Z(n4757) );
  XOR U4547 ( .A(n4759), .B(n4756), .Z(n4758) );
  XOR U4548 ( .A(n4760), .B(n4761), .Z(n4748) );
  AND U4549 ( .A(n4762), .B(n4763), .Z(n4761) );
  XOR U4550 ( .A(n4760), .B(n4586), .Z(n4763) );
  XOR U4551 ( .A(n4764), .B(n4765), .Z(n4586) );
  AND U4552 ( .A(n254), .B(n4766), .Z(n4765) );
  XOR U4553 ( .A(n4767), .B(n4764), .Z(n4766) );
  XNOR U4554 ( .A(n4583), .B(n4760), .Z(n4762) );
  XOR U4555 ( .A(n4768), .B(n4769), .Z(n4583) );
  AND U4556 ( .A(n252), .B(n4770), .Z(n4769) );
  XOR U4557 ( .A(n4771), .B(n4768), .Z(n4770) );
  XOR U4558 ( .A(n4772), .B(n4773), .Z(n4760) );
  AND U4559 ( .A(n4774), .B(n4775), .Z(n4773) );
  XOR U4560 ( .A(n4772), .B(n4598), .Z(n4775) );
  XOR U4561 ( .A(n4776), .B(n4777), .Z(n4598) );
  AND U4562 ( .A(n254), .B(n4778), .Z(n4777) );
  XOR U4563 ( .A(n4779), .B(n4776), .Z(n4778) );
  XNOR U4564 ( .A(n4595), .B(n4772), .Z(n4774) );
  XOR U4565 ( .A(n4780), .B(n4781), .Z(n4595) );
  AND U4566 ( .A(n252), .B(n4782), .Z(n4781) );
  XOR U4567 ( .A(n4783), .B(n4780), .Z(n4782) );
  XOR U4568 ( .A(n4784), .B(n4785), .Z(n4772) );
  AND U4569 ( .A(n4786), .B(n4787), .Z(n4785) );
  XOR U4570 ( .A(n4784), .B(n4610), .Z(n4787) );
  XOR U4571 ( .A(n4788), .B(n4789), .Z(n4610) );
  AND U4572 ( .A(n254), .B(n4790), .Z(n4789) );
  XOR U4573 ( .A(n4791), .B(n4788), .Z(n4790) );
  XNOR U4574 ( .A(n4607), .B(n4784), .Z(n4786) );
  XOR U4575 ( .A(n4792), .B(n4793), .Z(n4607) );
  AND U4576 ( .A(n252), .B(n4794), .Z(n4793) );
  XOR U4577 ( .A(n4795), .B(n4792), .Z(n4794) );
  XOR U4578 ( .A(n4796), .B(n4797), .Z(n4784) );
  AND U4579 ( .A(n4798), .B(n4799), .Z(n4797) );
  XOR U4580 ( .A(n4796), .B(n4622), .Z(n4799) );
  XOR U4581 ( .A(n4800), .B(n4801), .Z(n4622) );
  AND U4582 ( .A(n254), .B(n4802), .Z(n4801) );
  XOR U4583 ( .A(n4803), .B(n4800), .Z(n4802) );
  XNOR U4584 ( .A(n4619), .B(n4796), .Z(n4798) );
  XOR U4585 ( .A(n4804), .B(n4805), .Z(n4619) );
  AND U4586 ( .A(n252), .B(n4806), .Z(n4805) );
  XOR U4587 ( .A(n4807), .B(n4804), .Z(n4806) );
  XOR U4588 ( .A(n4808), .B(n4809), .Z(n4796) );
  AND U4589 ( .A(n4810), .B(n4811), .Z(n4809) );
  XOR U4590 ( .A(n4634), .B(n4808), .Z(n4811) );
  XOR U4591 ( .A(n4812), .B(n4813), .Z(n4634) );
  AND U4592 ( .A(n254), .B(n4814), .Z(n4813) );
  XOR U4593 ( .A(n4812), .B(n4815), .Z(n4814) );
  XNOR U4594 ( .A(n4808), .B(n4631), .Z(n4810) );
  XOR U4595 ( .A(n4816), .B(n4817), .Z(n4631) );
  AND U4596 ( .A(n252), .B(n4818), .Z(n4817) );
  XOR U4597 ( .A(n4816), .B(n4819), .Z(n4818) );
  XOR U4598 ( .A(n4820), .B(n4821), .Z(n4808) );
  AND U4599 ( .A(n4822), .B(n4823), .Z(n4821) );
  XNOR U4600 ( .A(n4824), .B(n4647), .Z(n4823) );
  XOR U4601 ( .A(n4825), .B(n4826), .Z(n4647) );
  AND U4602 ( .A(n254), .B(n4827), .Z(n4826) );
  XOR U4603 ( .A(n4828), .B(n4825), .Z(n4827) );
  XNOR U4604 ( .A(n4644), .B(n4820), .Z(n4822) );
  XOR U4605 ( .A(n4829), .B(n4830), .Z(n4644) );
  AND U4606 ( .A(n252), .B(n4831), .Z(n4830) );
  XOR U4607 ( .A(n4832), .B(n4829), .Z(n4831) );
  IV U4608 ( .A(n4824), .Z(n4820) );
  AND U4609 ( .A(n4652), .B(n4655), .Z(n4824) );
  XNOR U4610 ( .A(n4833), .B(n4834), .Z(n4655) );
  AND U4611 ( .A(n254), .B(n4835), .Z(n4834) );
  XNOR U4612 ( .A(n4836), .B(n4833), .Z(n4835) );
  XOR U4613 ( .A(n4837), .B(n4838), .Z(n254) );
  AND U4614 ( .A(n4839), .B(n4840), .Z(n4838) );
  XNOR U4615 ( .A(n4660), .B(n4837), .Z(n4840) );
  AND U4616 ( .A(p_input[1535]), .B(p_input[1519]), .Z(n4660) );
  XOR U4617 ( .A(n4837), .B(n4661), .Z(n4839) );
  AND U4618 ( .A(p_input[1503]), .B(p_input[1487]), .Z(n4661) );
  XOR U4619 ( .A(n4841), .B(n4842), .Z(n4837) );
  AND U4620 ( .A(n4843), .B(n4844), .Z(n4842) );
  XOR U4621 ( .A(n4841), .B(n4671), .Z(n4844) );
  XNOR U4622 ( .A(p_input[1518]), .B(n4845), .Z(n4671) );
  AND U4623 ( .A(n162), .B(n4846), .Z(n4845) );
  XOR U4624 ( .A(p_input[1534]), .B(p_input[1518]), .Z(n4846) );
  XNOR U4625 ( .A(n4668), .B(n4841), .Z(n4843) );
  XOR U4626 ( .A(n4847), .B(n4848), .Z(n4668) );
  AND U4627 ( .A(n160), .B(n4849), .Z(n4848) );
  XOR U4628 ( .A(p_input[1502]), .B(p_input[1486]), .Z(n4849) );
  XOR U4629 ( .A(n4850), .B(n4851), .Z(n4841) );
  AND U4630 ( .A(n4852), .B(n4853), .Z(n4851) );
  XOR U4631 ( .A(n4850), .B(n4683), .Z(n4853) );
  XNOR U4632 ( .A(p_input[1517]), .B(n4854), .Z(n4683) );
  AND U4633 ( .A(n162), .B(n4855), .Z(n4854) );
  XOR U4634 ( .A(p_input[1533]), .B(p_input[1517]), .Z(n4855) );
  XNOR U4635 ( .A(n4680), .B(n4850), .Z(n4852) );
  XOR U4636 ( .A(n4856), .B(n4857), .Z(n4680) );
  AND U4637 ( .A(n160), .B(n4858), .Z(n4857) );
  XOR U4638 ( .A(p_input[1501]), .B(p_input[1485]), .Z(n4858) );
  XOR U4639 ( .A(n4859), .B(n4860), .Z(n4850) );
  AND U4640 ( .A(n4861), .B(n4862), .Z(n4860) );
  XOR U4641 ( .A(n4859), .B(n4695), .Z(n4862) );
  XNOR U4642 ( .A(p_input[1516]), .B(n4863), .Z(n4695) );
  AND U4643 ( .A(n162), .B(n4864), .Z(n4863) );
  XOR U4644 ( .A(p_input[1532]), .B(p_input[1516]), .Z(n4864) );
  XNOR U4645 ( .A(n4692), .B(n4859), .Z(n4861) );
  XOR U4646 ( .A(n4865), .B(n4866), .Z(n4692) );
  AND U4647 ( .A(n160), .B(n4867), .Z(n4866) );
  XOR U4648 ( .A(p_input[1500]), .B(p_input[1484]), .Z(n4867) );
  XOR U4649 ( .A(n4868), .B(n4869), .Z(n4859) );
  AND U4650 ( .A(n4870), .B(n4871), .Z(n4869) );
  XOR U4651 ( .A(n4868), .B(n4707), .Z(n4871) );
  XNOR U4652 ( .A(p_input[1515]), .B(n4872), .Z(n4707) );
  AND U4653 ( .A(n162), .B(n4873), .Z(n4872) );
  XOR U4654 ( .A(p_input[1531]), .B(p_input[1515]), .Z(n4873) );
  XNOR U4655 ( .A(n4704), .B(n4868), .Z(n4870) );
  XOR U4656 ( .A(n4874), .B(n4875), .Z(n4704) );
  AND U4657 ( .A(n160), .B(n4876), .Z(n4875) );
  XOR U4658 ( .A(p_input[1499]), .B(p_input[1483]), .Z(n4876) );
  XOR U4659 ( .A(n4877), .B(n4878), .Z(n4868) );
  AND U4660 ( .A(n4879), .B(n4880), .Z(n4878) );
  XOR U4661 ( .A(n4877), .B(n4719), .Z(n4880) );
  XNOR U4662 ( .A(p_input[1514]), .B(n4881), .Z(n4719) );
  AND U4663 ( .A(n162), .B(n4882), .Z(n4881) );
  XOR U4664 ( .A(p_input[1530]), .B(p_input[1514]), .Z(n4882) );
  XNOR U4665 ( .A(n4716), .B(n4877), .Z(n4879) );
  XOR U4666 ( .A(n4883), .B(n4884), .Z(n4716) );
  AND U4667 ( .A(n160), .B(n4885), .Z(n4884) );
  XOR U4668 ( .A(p_input[1498]), .B(p_input[1482]), .Z(n4885) );
  XOR U4669 ( .A(n4886), .B(n4887), .Z(n4877) );
  AND U4670 ( .A(n4888), .B(n4889), .Z(n4887) );
  XOR U4671 ( .A(n4886), .B(n4731), .Z(n4889) );
  XNOR U4672 ( .A(p_input[1513]), .B(n4890), .Z(n4731) );
  AND U4673 ( .A(n162), .B(n4891), .Z(n4890) );
  XOR U4674 ( .A(p_input[1529]), .B(p_input[1513]), .Z(n4891) );
  XNOR U4675 ( .A(n4728), .B(n4886), .Z(n4888) );
  XOR U4676 ( .A(n4892), .B(n4893), .Z(n4728) );
  AND U4677 ( .A(n160), .B(n4894), .Z(n4893) );
  XOR U4678 ( .A(p_input[1497]), .B(p_input[1481]), .Z(n4894) );
  XOR U4679 ( .A(n4895), .B(n4896), .Z(n4886) );
  AND U4680 ( .A(n4897), .B(n4898), .Z(n4896) );
  XOR U4681 ( .A(n4895), .B(n4743), .Z(n4898) );
  XNOR U4682 ( .A(p_input[1512]), .B(n4899), .Z(n4743) );
  AND U4683 ( .A(n162), .B(n4900), .Z(n4899) );
  XOR U4684 ( .A(p_input[1528]), .B(p_input[1512]), .Z(n4900) );
  XNOR U4685 ( .A(n4740), .B(n4895), .Z(n4897) );
  XOR U4686 ( .A(n4901), .B(n4902), .Z(n4740) );
  AND U4687 ( .A(n160), .B(n4903), .Z(n4902) );
  XOR U4688 ( .A(p_input[1496]), .B(p_input[1480]), .Z(n4903) );
  XOR U4689 ( .A(n4904), .B(n4905), .Z(n4895) );
  AND U4690 ( .A(n4906), .B(n4907), .Z(n4905) );
  XOR U4691 ( .A(n4904), .B(n4755), .Z(n4907) );
  XNOR U4692 ( .A(p_input[1511]), .B(n4908), .Z(n4755) );
  AND U4693 ( .A(n162), .B(n4909), .Z(n4908) );
  XOR U4694 ( .A(p_input[1527]), .B(p_input[1511]), .Z(n4909) );
  XNOR U4695 ( .A(n4752), .B(n4904), .Z(n4906) );
  XOR U4696 ( .A(n4910), .B(n4911), .Z(n4752) );
  AND U4697 ( .A(n160), .B(n4912), .Z(n4911) );
  XOR U4698 ( .A(p_input[1495]), .B(p_input[1479]), .Z(n4912) );
  XOR U4699 ( .A(n4913), .B(n4914), .Z(n4904) );
  AND U4700 ( .A(n4915), .B(n4916), .Z(n4914) );
  XOR U4701 ( .A(n4913), .B(n4767), .Z(n4916) );
  XNOR U4702 ( .A(p_input[1510]), .B(n4917), .Z(n4767) );
  AND U4703 ( .A(n162), .B(n4918), .Z(n4917) );
  XOR U4704 ( .A(p_input[1526]), .B(p_input[1510]), .Z(n4918) );
  XNOR U4705 ( .A(n4764), .B(n4913), .Z(n4915) );
  XOR U4706 ( .A(n4919), .B(n4920), .Z(n4764) );
  AND U4707 ( .A(n160), .B(n4921), .Z(n4920) );
  XOR U4708 ( .A(p_input[1494]), .B(p_input[1478]), .Z(n4921) );
  XOR U4709 ( .A(n4922), .B(n4923), .Z(n4913) );
  AND U4710 ( .A(n4924), .B(n4925), .Z(n4923) );
  XOR U4711 ( .A(n4922), .B(n4779), .Z(n4925) );
  XNOR U4712 ( .A(p_input[1509]), .B(n4926), .Z(n4779) );
  AND U4713 ( .A(n162), .B(n4927), .Z(n4926) );
  XOR U4714 ( .A(p_input[1525]), .B(p_input[1509]), .Z(n4927) );
  XNOR U4715 ( .A(n4776), .B(n4922), .Z(n4924) );
  XOR U4716 ( .A(n4928), .B(n4929), .Z(n4776) );
  AND U4717 ( .A(n160), .B(n4930), .Z(n4929) );
  XOR U4718 ( .A(p_input[1493]), .B(p_input[1477]), .Z(n4930) );
  XOR U4719 ( .A(n4931), .B(n4932), .Z(n4922) );
  AND U4720 ( .A(n4933), .B(n4934), .Z(n4932) );
  XOR U4721 ( .A(n4931), .B(n4791), .Z(n4934) );
  XNOR U4722 ( .A(p_input[1508]), .B(n4935), .Z(n4791) );
  AND U4723 ( .A(n162), .B(n4936), .Z(n4935) );
  XOR U4724 ( .A(p_input[1524]), .B(p_input[1508]), .Z(n4936) );
  XNOR U4725 ( .A(n4788), .B(n4931), .Z(n4933) );
  XOR U4726 ( .A(n4937), .B(n4938), .Z(n4788) );
  AND U4727 ( .A(n160), .B(n4939), .Z(n4938) );
  XOR U4728 ( .A(p_input[1492]), .B(p_input[1476]), .Z(n4939) );
  XOR U4729 ( .A(n4940), .B(n4941), .Z(n4931) );
  AND U4730 ( .A(n4942), .B(n4943), .Z(n4941) );
  XOR U4731 ( .A(n4940), .B(n4803), .Z(n4943) );
  XNOR U4732 ( .A(p_input[1507]), .B(n4944), .Z(n4803) );
  AND U4733 ( .A(n162), .B(n4945), .Z(n4944) );
  XOR U4734 ( .A(p_input[1523]), .B(p_input[1507]), .Z(n4945) );
  XNOR U4735 ( .A(n4800), .B(n4940), .Z(n4942) );
  XOR U4736 ( .A(n4946), .B(n4947), .Z(n4800) );
  AND U4737 ( .A(n160), .B(n4948), .Z(n4947) );
  XOR U4738 ( .A(p_input[1491]), .B(p_input[1475]), .Z(n4948) );
  XOR U4739 ( .A(n4949), .B(n4950), .Z(n4940) );
  AND U4740 ( .A(n4951), .B(n4952), .Z(n4950) );
  XOR U4741 ( .A(n4815), .B(n4949), .Z(n4952) );
  XNOR U4742 ( .A(p_input[1506]), .B(n4953), .Z(n4815) );
  AND U4743 ( .A(n162), .B(n4954), .Z(n4953) );
  XOR U4744 ( .A(p_input[1522]), .B(p_input[1506]), .Z(n4954) );
  XNOR U4745 ( .A(n4949), .B(n4812), .Z(n4951) );
  XOR U4746 ( .A(n4955), .B(n4956), .Z(n4812) );
  AND U4747 ( .A(n160), .B(n4957), .Z(n4956) );
  XOR U4748 ( .A(p_input[1490]), .B(p_input[1474]), .Z(n4957) );
  XOR U4749 ( .A(n4958), .B(n4959), .Z(n4949) );
  AND U4750 ( .A(n4960), .B(n4961), .Z(n4959) );
  XNOR U4751 ( .A(n4962), .B(n4828), .Z(n4961) );
  XNOR U4752 ( .A(p_input[1505]), .B(n4963), .Z(n4828) );
  AND U4753 ( .A(n162), .B(n4964), .Z(n4963) );
  XNOR U4754 ( .A(p_input[1521]), .B(n4965), .Z(n4964) );
  IV U4755 ( .A(p_input[1505]), .Z(n4965) );
  XNOR U4756 ( .A(n4825), .B(n4958), .Z(n4960) );
  XNOR U4757 ( .A(p_input[1473]), .B(n4966), .Z(n4825) );
  AND U4758 ( .A(n160), .B(n4967), .Z(n4966) );
  XOR U4759 ( .A(p_input[1489]), .B(p_input[1473]), .Z(n4967) );
  IV U4760 ( .A(n4962), .Z(n4958) );
  AND U4761 ( .A(n4833), .B(n4836), .Z(n4962) );
  XOR U4762 ( .A(p_input[1504]), .B(n4968), .Z(n4836) );
  AND U4763 ( .A(n162), .B(n4969), .Z(n4968) );
  XOR U4764 ( .A(p_input[1520]), .B(p_input[1504]), .Z(n4969) );
  XOR U4765 ( .A(n4970), .B(n4971), .Z(n162) );
  AND U4766 ( .A(n4972), .B(n4973), .Z(n4971) );
  XNOR U4767 ( .A(p_input[1535]), .B(n4970), .Z(n4973) );
  XOR U4768 ( .A(n4970), .B(p_input[1519]), .Z(n4972) );
  XOR U4769 ( .A(n4974), .B(n4975), .Z(n4970) );
  AND U4770 ( .A(n4976), .B(n4977), .Z(n4975) );
  XNOR U4771 ( .A(p_input[1534]), .B(n4974), .Z(n4977) );
  XOR U4772 ( .A(n4974), .B(p_input[1518]), .Z(n4976) );
  XOR U4773 ( .A(n4978), .B(n4979), .Z(n4974) );
  AND U4774 ( .A(n4980), .B(n4981), .Z(n4979) );
  XNOR U4775 ( .A(p_input[1533]), .B(n4978), .Z(n4981) );
  XOR U4776 ( .A(n4978), .B(p_input[1517]), .Z(n4980) );
  XOR U4777 ( .A(n4982), .B(n4983), .Z(n4978) );
  AND U4778 ( .A(n4984), .B(n4985), .Z(n4983) );
  XNOR U4779 ( .A(p_input[1532]), .B(n4982), .Z(n4985) );
  XOR U4780 ( .A(n4982), .B(p_input[1516]), .Z(n4984) );
  XOR U4781 ( .A(n4986), .B(n4987), .Z(n4982) );
  AND U4782 ( .A(n4988), .B(n4989), .Z(n4987) );
  XNOR U4783 ( .A(p_input[1531]), .B(n4986), .Z(n4989) );
  XOR U4784 ( .A(n4986), .B(p_input[1515]), .Z(n4988) );
  XOR U4785 ( .A(n4990), .B(n4991), .Z(n4986) );
  AND U4786 ( .A(n4992), .B(n4993), .Z(n4991) );
  XNOR U4787 ( .A(p_input[1530]), .B(n4990), .Z(n4993) );
  XOR U4788 ( .A(n4990), .B(p_input[1514]), .Z(n4992) );
  XOR U4789 ( .A(n4994), .B(n4995), .Z(n4990) );
  AND U4790 ( .A(n4996), .B(n4997), .Z(n4995) );
  XNOR U4791 ( .A(p_input[1529]), .B(n4994), .Z(n4997) );
  XOR U4792 ( .A(n4994), .B(p_input[1513]), .Z(n4996) );
  XOR U4793 ( .A(n4998), .B(n4999), .Z(n4994) );
  AND U4794 ( .A(n5000), .B(n5001), .Z(n4999) );
  XNOR U4795 ( .A(p_input[1528]), .B(n4998), .Z(n5001) );
  XOR U4796 ( .A(n4998), .B(p_input[1512]), .Z(n5000) );
  XOR U4797 ( .A(n5002), .B(n5003), .Z(n4998) );
  AND U4798 ( .A(n5004), .B(n5005), .Z(n5003) );
  XNOR U4799 ( .A(p_input[1527]), .B(n5002), .Z(n5005) );
  XOR U4800 ( .A(n5002), .B(p_input[1511]), .Z(n5004) );
  XOR U4801 ( .A(n5006), .B(n5007), .Z(n5002) );
  AND U4802 ( .A(n5008), .B(n5009), .Z(n5007) );
  XNOR U4803 ( .A(p_input[1526]), .B(n5006), .Z(n5009) );
  XOR U4804 ( .A(n5006), .B(p_input[1510]), .Z(n5008) );
  XOR U4805 ( .A(n5010), .B(n5011), .Z(n5006) );
  AND U4806 ( .A(n5012), .B(n5013), .Z(n5011) );
  XNOR U4807 ( .A(p_input[1525]), .B(n5010), .Z(n5013) );
  XOR U4808 ( .A(n5010), .B(p_input[1509]), .Z(n5012) );
  XOR U4809 ( .A(n5014), .B(n5015), .Z(n5010) );
  AND U4810 ( .A(n5016), .B(n5017), .Z(n5015) );
  XNOR U4811 ( .A(p_input[1524]), .B(n5014), .Z(n5017) );
  XOR U4812 ( .A(n5014), .B(p_input[1508]), .Z(n5016) );
  XOR U4813 ( .A(n5018), .B(n5019), .Z(n5014) );
  AND U4814 ( .A(n5020), .B(n5021), .Z(n5019) );
  XNOR U4815 ( .A(p_input[1523]), .B(n5018), .Z(n5021) );
  XOR U4816 ( .A(n5018), .B(p_input[1507]), .Z(n5020) );
  XOR U4817 ( .A(n5022), .B(n5023), .Z(n5018) );
  AND U4818 ( .A(n5024), .B(n5025), .Z(n5023) );
  XNOR U4819 ( .A(p_input[1522]), .B(n5022), .Z(n5025) );
  XOR U4820 ( .A(n5022), .B(p_input[1506]), .Z(n5024) );
  XNOR U4821 ( .A(n5026), .B(n5027), .Z(n5022) );
  AND U4822 ( .A(n5028), .B(n5029), .Z(n5027) );
  XOR U4823 ( .A(p_input[1521]), .B(n5026), .Z(n5029) );
  XNOR U4824 ( .A(p_input[1505]), .B(n5026), .Z(n5028) );
  AND U4825 ( .A(p_input[1520]), .B(n5030), .Z(n5026) );
  IV U4826 ( .A(p_input[1504]), .Z(n5030) );
  XNOR U4827 ( .A(p_input[1472]), .B(n5031), .Z(n4833) );
  AND U4828 ( .A(n160), .B(n5032), .Z(n5031) );
  XOR U4829 ( .A(p_input[1488]), .B(p_input[1472]), .Z(n5032) );
  XOR U4830 ( .A(n5033), .B(n5034), .Z(n160) );
  AND U4831 ( .A(n5035), .B(n5036), .Z(n5034) );
  XNOR U4832 ( .A(p_input[1503]), .B(n5033), .Z(n5036) );
  XOR U4833 ( .A(n5033), .B(p_input[1487]), .Z(n5035) );
  XOR U4834 ( .A(n5037), .B(n5038), .Z(n5033) );
  AND U4835 ( .A(n5039), .B(n5040), .Z(n5038) );
  XNOR U4836 ( .A(p_input[1502]), .B(n5037), .Z(n5040) );
  XNOR U4837 ( .A(n5037), .B(n4847), .Z(n5039) );
  IV U4838 ( .A(p_input[1486]), .Z(n4847) );
  XOR U4839 ( .A(n5041), .B(n5042), .Z(n5037) );
  AND U4840 ( .A(n5043), .B(n5044), .Z(n5042) );
  XNOR U4841 ( .A(p_input[1501]), .B(n5041), .Z(n5044) );
  XNOR U4842 ( .A(n5041), .B(n4856), .Z(n5043) );
  IV U4843 ( .A(p_input[1485]), .Z(n4856) );
  XOR U4844 ( .A(n5045), .B(n5046), .Z(n5041) );
  AND U4845 ( .A(n5047), .B(n5048), .Z(n5046) );
  XNOR U4846 ( .A(p_input[1500]), .B(n5045), .Z(n5048) );
  XNOR U4847 ( .A(n5045), .B(n4865), .Z(n5047) );
  IV U4848 ( .A(p_input[1484]), .Z(n4865) );
  XOR U4849 ( .A(n5049), .B(n5050), .Z(n5045) );
  AND U4850 ( .A(n5051), .B(n5052), .Z(n5050) );
  XNOR U4851 ( .A(p_input[1499]), .B(n5049), .Z(n5052) );
  XNOR U4852 ( .A(n5049), .B(n4874), .Z(n5051) );
  IV U4853 ( .A(p_input[1483]), .Z(n4874) );
  XOR U4854 ( .A(n5053), .B(n5054), .Z(n5049) );
  AND U4855 ( .A(n5055), .B(n5056), .Z(n5054) );
  XNOR U4856 ( .A(p_input[1498]), .B(n5053), .Z(n5056) );
  XNOR U4857 ( .A(n5053), .B(n4883), .Z(n5055) );
  IV U4858 ( .A(p_input[1482]), .Z(n4883) );
  XOR U4859 ( .A(n5057), .B(n5058), .Z(n5053) );
  AND U4860 ( .A(n5059), .B(n5060), .Z(n5058) );
  XNOR U4861 ( .A(p_input[1497]), .B(n5057), .Z(n5060) );
  XNOR U4862 ( .A(n5057), .B(n4892), .Z(n5059) );
  IV U4863 ( .A(p_input[1481]), .Z(n4892) );
  XOR U4864 ( .A(n5061), .B(n5062), .Z(n5057) );
  AND U4865 ( .A(n5063), .B(n5064), .Z(n5062) );
  XNOR U4866 ( .A(p_input[1496]), .B(n5061), .Z(n5064) );
  XNOR U4867 ( .A(n5061), .B(n4901), .Z(n5063) );
  IV U4868 ( .A(p_input[1480]), .Z(n4901) );
  XOR U4869 ( .A(n5065), .B(n5066), .Z(n5061) );
  AND U4870 ( .A(n5067), .B(n5068), .Z(n5066) );
  XNOR U4871 ( .A(p_input[1495]), .B(n5065), .Z(n5068) );
  XNOR U4872 ( .A(n5065), .B(n4910), .Z(n5067) );
  IV U4873 ( .A(p_input[1479]), .Z(n4910) );
  XOR U4874 ( .A(n5069), .B(n5070), .Z(n5065) );
  AND U4875 ( .A(n5071), .B(n5072), .Z(n5070) );
  XNOR U4876 ( .A(p_input[1494]), .B(n5069), .Z(n5072) );
  XNOR U4877 ( .A(n5069), .B(n4919), .Z(n5071) );
  IV U4878 ( .A(p_input[1478]), .Z(n4919) );
  XOR U4879 ( .A(n5073), .B(n5074), .Z(n5069) );
  AND U4880 ( .A(n5075), .B(n5076), .Z(n5074) );
  XNOR U4881 ( .A(p_input[1493]), .B(n5073), .Z(n5076) );
  XNOR U4882 ( .A(n5073), .B(n4928), .Z(n5075) );
  IV U4883 ( .A(p_input[1477]), .Z(n4928) );
  XOR U4884 ( .A(n5077), .B(n5078), .Z(n5073) );
  AND U4885 ( .A(n5079), .B(n5080), .Z(n5078) );
  XNOR U4886 ( .A(p_input[1492]), .B(n5077), .Z(n5080) );
  XNOR U4887 ( .A(n5077), .B(n4937), .Z(n5079) );
  IV U4888 ( .A(p_input[1476]), .Z(n4937) );
  XOR U4889 ( .A(n5081), .B(n5082), .Z(n5077) );
  AND U4890 ( .A(n5083), .B(n5084), .Z(n5082) );
  XNOR U4891 ( .A(p_input[1491]), .B(n5081), .Z(n5084) );
  XNOR U4892 ( .A(n5081), .B(n4946), .Z(n5083) );
  IV U4893 ( .A(p_input[1475]), .Z(n4946) );
  XOR U4894 ( .A(n5085), .B(n5086), .Z(n5081) );
  AND U4895 ( .A(n5087), .B(n5088), .Z(n5086) );
  XNOR U4896 ( .A(p_input[1490]), .B(n5085), .Z(n5088) );
  XNOR U4897 ( .A(n5085), .B(n4955), .Z(n5087) );
  IV U4898 ( .A(p_input[1474]), .Z(n4955) );
  XNOR U4899 ( .A(n5089), .B(n5090), .Z(n5085) );
  AND U4900 ( .A(n5091), .B(n5092), .Z(n5090) );
  XOR U4901 ( .A(p_input[1489]), .B(n5089), .Z(n5092) );
  XNOR U4902 ( .A(p_input[1473]), .B(n5089), .Z(n5091) );
  AND U4903 ( .A(p_input[1488]), .B(n5093), .Z(n5089) );
  IV U4904 ( .A(p_input[1472]), .Z(n5093) );
  XOR U4905 ( .A(n5094), .B(n5095), .Z(n4652) );
  AND U4906 ( .A(n252), .B(n5096), .Z(n5095) );
  XNOR U4907 ( .A(n5097), .B(n5094), .Z(n5096) );
  XOR U4908 ( .A(n5098), .B(n5099), .Z(n252) );
  AND U4909 ( .A(n5100), .B(n5101), .Z(n5099) );
  XNOR U4910 ( .A(n4662), .B(n5098), .Z(n5101) );
  AND U4911 ( .A(p_input[1471]), .B(p_input[1455]), .Z(n4662) );
  XOR U4912 ( .A(n5098), .B(n4663), .Z(n5100) );
  AND U4913 ( .A(p_input[1439]), .B(p_input[1423]), .Z(n4663) );
  XOR U4914 ( .A(n5102), .B(n5103), .Z(n5098) );
  AND U4915 ( .A(n5104), .B(n5105), .Z(n5103) );
  XOR U4916 ( .A(n5102), .B(n4675), .Z(n5105) );
  XNOR U4917 ( .A(p_input[1454]), .B(n5106), .Z(n4675) );
  AND U4918 ( .A(n166), .B(n5107), .Z(n5106) );
  XOR U4919 ( .A(p_input[1470]), .B(p_input[1454]), .Z(n5107) );
  XNOR U4920 ( .A(n4672), .B(n5102), .Z(n5104) );
  XOR U4921 ( .A(n5108), .B(n5109), .Z(n4672) );
  AND U4922 ( .A(n163), .B(n5110), .Z(n5109) );
  XOR U4923 ( .A(p_input[1438]), .B(p_input[1422]), .Z(n5110) );
  XOR U4924 ( .A(n5111), .B(n5112), .Z(n5102) );
  AND U4925 ( .A(n5113), .B(n5114), .Z(n5112) );
  XOR U4926 ( .A(n5111), .B(n4687), .Z(n5114) );
  XNOR U4927 ( .A(p_input[1453]), .B(n5115), .Z(n4687) );
  AND U4928 ( .A(n166), .B(n5116), .Z(n5115) );
  XOR U4929 ( .A(p_input[1469]), .B(p_input[1453]), .Z(n5116) );
  XNOR U4930 ( .A(n4684), .B(n5111), .Z(n5113) );
  XOR U4931 ( .A(n5117), .B(n5118), .Z(n4684) );
  AND U4932 ( .A(n163), .B(n5119), .Z(n5118) );
  XOR U4933 ( .A(p_input[1437]), .B(p_input[1421]), .Z(n5119) );
  XOR U4934 ( .A(n5120), .B(n5121), .Z(n5111) );
  AND U4935 ( .A(n5122), .B(n5123), .Z(n5121) );
  XOR U4936 ( .A(n5120), .B(n4699), .Z(n5123) );
  XNOR U4937 ( .A(p_input[1452]), .B(n5124), .Z(n4699) );
  AND U4938 ( .A(n166), .B(n5125), .Z(n5124) );
  XOR U4939 ( .A(p_input[1468]), .B(p_input[1452]), .Z(n5125) );
  XNOR U4940 ( .A(n4696), .B(n5120), .Z(n5122) );
  XOR U4941 ( .A(n5126), .B(n5127), .Z(n4696) );
  AND U4942 ( .A(n163), .B(n5128), .Z(n5127) );
  XOR U4943 ( .A(p_input[1436]), .B(p_input[1420]), .Z(n5128) );
  XOR U4944 ( .A(n5129), .B(n5130), .Z(n5120) );
  AND U4945 ( .A(n5131), .B(n5132), .Z(n5130) );
  XOR U4946 ( .A(n5129), .B(n4711), .Z(n5132) );
  XNOR U4947 ( .A(p_input[1451]), .B(n5133), .Z(n4711) );
  AND U4948 ( .A(n166), .B(n5134), .Z(n5133) );
  XOR U4949 ( .A(p_input[1467]), .B(p_input[1451]), .Z(n5134) );
  XNOR U4950 ( .A(n4708), .B(n5129), .Z(n5131) );
  XOR U4951 ( .A(n5135), .B(n5136), .Z(n4708) );
  AND U4952 ( .A(n163), .B(n5137), .Z(n5136) );
  XOR U4953 ( .A(p_input[1435]), .B(p_input[1419]), .Z(n5137) );
  XOR U4954 ( .A(n5138), .B(n5139), .Z(n5129) );
  AND U4955 ( .A(n5140), .B(n5141), .Z(n5139) );
  XOR U4956 ( .A(n5138), .B(n4723), .Z(n5141) );
  XNOR U4957 ( .A(p_input[1450]), .B(n5142), .Z(n4723) );
  AND U4958 ( .A(n166), .B(n5143), .Z(n5142) );
  XOR U4959 ( .A(p_input[1466]), .B(p_input[1450]), .Z(n5143) );
  XNOR U4960 ( .A(n4720), .B(n5138), .Z(n5140) );
  XOR U4961 ( .A(n5144), .B(n5145), .Z(n4720) );
  AND U4962 ( .A(n163), .B(n5146), .Z(n5145) );
  XOR U4963 ( .A(p_input[1434]), .B(p_input[1418]), .Z(n5146) );
  XOR U4964 ( .A(n5147), .B(n5148), .Z(n5138) );
  AND U4965 ( .A(n5149), .B(n5150), .Z(n5148) );
  XOR U4966 ( .A(n5147), .B(n4735), .Z(n5150) );
  XNOR U4967 ( .A(p_input[1449]), .B(n5151), .Z(n4735) );
  AND U4968 ( .A(n166), .B(n5152), .Z(n5151) );
  XOR U4969 ( .A(p_input[1465]), .B(p_input[1449]), .Z(n5152) );
  XNOR U4970 ( .A(n4732), .B(n5147), .Z(n5149) );
  XOR U4971 ( .A(n5153), .B(n5154), .Z(n4732) );
  AND U4972 ( .A(n163), .B(n5155), .Z(n5154) );
  XOR U4973 ( .A(p_input[1433]), .B(p_input[1417]), .Z(n5155) );
  XOR U4974 ( .A(n5156), .B(n5157), .Z(n5147) );
  AND U4975 ( .A(n5158), .B(n5159), .Z(n5157) );
  XOR U4976 ( .A(n5156), .B(n4747), .Z(n5159) );
  XNOR U4977 ( .A(p_input[1448]), .B(n5160), .Z(n4747) );
  AND U4978 ( .A(n166), .B(n5161), .Z(n5160) );
  XOR U4979 ( .A(p_input[1464]), .B(p_input[1448]), .Z(n5161) );
  XNOR U4980 ( .A(n4744), .B(n5156), .Z(n5158) );
  XOR U4981 ( .A(n5162), .B(n5163), .Z(n4744) );
  AND U4982 ( .A(n163), .B(n5164), .Z(n5163) );
  XOR U4983 ( .A(p_input[1432]), .B(p_input[1416]), .Z(n5164) );
  XOR U4984 ( .A(n5165), .B(n5166), .Z(n5156) );
  AND U4985 ( .A(n5167), .B(n5168), .Z(n5166) );
  XOR U4986 ( .A(n5165), .B(n4759), .Z(n5168) );
  XNOR U4987 ( .A(p_input[1447]), .B(n5169), .Z(n4759) );
  AND U4988 ( .A(n166), .B(n5170), .Z(n5169) );
  XOR U4989 ( .A(p_input[1463]), .B(p_input[1447]), .Z(n5170) );
  XNOR U4990 ( .A(n4756), .B(n5165), .Z(n5167) );
  XOR U4991 ( .A(n5171), .B(n5172), .Z(n4756) );
  AND U4992 ( .A(n163), .B(n5173), .Z(n5172) );
  XOR U4993 ( .A(p_input[1431]), .B(p_input[1415]), .Z(n5173) );
  XOR U4994 ( .A(n5174), .B(n5175), .Z(n5165) );
  AND U4995 ( .A(n5176), .B(n5177), .Z(n5175) );
  XOR U4996 ( .A(n5174), .B(n4771), .Z(n5177) );
  XNOR U4997 ( .A(p_input[1446]), .B(n5178), .Z(n4771) );
  AND U4998 ( .A(n166), .B(n5179), .Z(n5178) );
  XOR U4999 ( .A(p_input[1462]), .B(p_input[1446]), .Z(n5179) );
  XNOR U5000 ( .A(n4768), .B(n5174), .Z(n5176) );
  XOR U5001 ( .A(n5180), .B(n5181), .Z(n4768) );
  AND U5002 ( .A(n163), .B(n5182), .Z(n5181) );
  XOR U5003 ( .A(p_input[1430]), .B(p_input[1414]), .Z(n5182) );
  XOR U5004 ( .A(n5183), .B(n5184), .Z(n5174) );
  AND U5005 ( .A(n5185), .B(n5186), .Z(n5184) );
  XOR U5006 ( .A(n5183), .B(n4783), .Z(n5186) );
  XNOR U5007 ( .A(p_input[1445]), .B(n5187), .Z(n4783) );
  AND U5008 ( .A(n166), .B(n5188), .Z(n5187) );
  XOR U5009 ( .A(p_input[1461]), .B(p_input[1445]), .Z(n5188) );
  XNOR U5010 ( .A(n4780), .B(n5183), .Z(n5185) );
  XOR U5011 ( .A(n5189), .B(n5190), .Z(n4780) );
  AND U5012 ( .A(n163), .B(n5191), .Z(n5190) );
  XOR U5013 ( .A(p_input[1429]), .B(p_input[1413]), .Z(n5191) );
  XOR U5014 ( .A(n5192), .B(n5193), .Z(n5183) );
  AND U5015 ( .A(n5194), .B(n5195), .Z(n5193) );
  XOR U5016 ( .A(n5192), .B(n4795), .Z(n5195) );
  XNOR U5017 ( .A(p_input[1444]), .B(n5196), .Z(n4795) );
  AND U5018 ( .A(n166), .B(n5197), .Z(n5196) );
  XOR U5019 ( .A(p_input[1460]), .B(p_input[1444]), .Z(n5197) );
  XNOR U5020 ( .A(n4792), .B(n5192), .Z(n5194) );
  XOR U5021 ( .A(n5198), .B(n5199), .Z(n4792) );
  AND U5022 ( .A(n163), .B(n5200), .Z(n5199) );
  XOR U5023 ( .A(p_input[1428]), .B(p_input[1412]), .Z(n5200) );
  XOR U5024 ( .A(n5201), .B(n5202), .Z(n5192) );
  AND U5025 ( .A(n5203), .B(n5204), .Z(n5202) );
  XOR U5026 ( .A(n5201), .B(n4807), .Z(n5204) );
  XNOR U5027 ( .A(p_input[1443]), .B(n5205), .Z(n4807) );
  AND U5028 ( .A(n166), .B(n5206), .Z(n5205) );
  XOR U5029 ( .A(p_input[1459]), .B(p_input[1443]), .Z(n5206) );
  XNOR U5030 ( .A(n4804), .B(n5201), .Z(n5203) );
  XOR U5031 ( .A(n5207), .B(n5208), .Z(n4804) );
  AND U5032 ( .A(n163), .B(n5209), .Z(n5208) );
  XOR U5033 ( .A(p_input[1427]), .B(p_input[1411]), .Z(n5209) );
  XOR U5034 ( .A(n5210), .B(n5211), .Z(n5201) );
  AND U5035 ( .A(n5212), .B(n5213), .Z(n5211) );
  XOR U5036 ( .A(n4819), .B(n5210), .Z(n5213) );
  XNOR U5037 ( .A(p_input[1442]), .B(n5214), .Z(n4819) );
  AND U5038 ( .A(n166), .B(n5215), .Z(n5214) );
  XOR U5039 ( .A(p_input[1458]), .B(p_input[1442]), .Z(n5215) );
  XNOR U5040 ( .A(n5210), .B(n4816), .Z(n5212) );
  XOR U5041 ( .A(n5216), .B(n5217), .Z(n4816) );
  AND U5042 ( .A(n163), .B(n5218), .Z(n5217) );
  XOR U5043 ( .A(p_input[1426]), .B(p_input[1410]), .Z(n5218) );
  XOR U5044 ( .A(n5219), .B(n5220), .Z(n5210) );
  AND U5045 ( .A(n5221), .B(n5222), .Z(n5220) );
  XNOR U5046 ( .A(n5223), .B(n4832), .Z(n5222) );
  XNOR U5047 ( .A(p_input[1441]), .B(n5224), .Z(n4832) );
  AND U5048 ( .A(n166), .B(n5225), .Z(n5224) );
  XNOR U5049 ( .A(p_input[1457]), .B(n5226), .Z(n5225) );
  IV U5050 ( .A(p_input[1441]), .Z(n5226) );
  XNOR U5051 ( .A(n4829), .B(n5219), .Z(n5221) );
  XNOR U5052 ( .A(p_input[1409]), .B(n5227), .Z(n4829) );
  AND U5053 ( .A(n163), .B(n5228), .Z(n5227) );
  XOR U5054 ( .A(p_input[1425]), .B(p_input[1409]), .Z(n5228) );
  IV U5055 ( .A(n5223), .Z(n5219) );
  AND U5056 ( .A(n5094), .B(n5097), .Z(n5223) );
  XOR U5057 ( .A(p_input[1440]), .B(n5229), .Z(n5097) );
  AND U5058 ( .A(n166), .B(n5230), .Z(n5229) );
  XOR U5059 ( .A(p_input[1456]), .B(p_input[1440]), .Z(n5230) );
  XOR U5060 ( .A(n5231), .B(n5232), .Z(n166) );
  AND U5061 ( .A(n5233), .B(n5234), .Z(n5232) );
  XNOR U5062 ( .A(p_input[1471]), .B(n5231), .Z(n5234) );
  XOR U5063 ( .A(n5231), .B(p_input[1455]), .Z(n5233) );
  XOR U5064 ( .A(n5235), .B(n5236), .Z(n5231) );
  AND U5065 ( .A(n5237), .B(n5238), .Z(n5236) );
  XNOR U5066 ( .A(p_input[1470]), .B(n5235), .Z(n5238) );
  XOR U5067 ( .A(n5235), .B(p_input[1454]), .Z(n5237) );
  XOR U5068 ( .A(n5239), .B(n5240), .Z(n5235) );
  AND U5069 ( .A(n5241), .B(n5242), .Z(n5240) );
  XNOR U5070 ( .A(p_input[1469]), .B(n5239), .Z(n5242) );
  XOR U5071 ( .A(n5239), .B(p_input[1453]), .Z(n5241) );
  XOR U5072 ( .A(n5243), .B(n5244), .Z(n5239) );
  AND U5073 ( .A(n5245), .B(n5246), .Z(n5244) );
  XNOR U5074 ( .A(p_input[1468]), .B(n5243), .Z(n5246) );
  XOR U5075 ( .A(n5243), .B(p_input[1452]), .Z(n5245) );
  XOR U5076 ( .A(n5247), .B(n5248), .Z(n5243) );
  AND U5077 ( .A(n5249), .B(n5250), .Z(n5248) );
  XNOR U5078 ( .A(p_input[1467]), .B(n5247), .Z(n5250) );
  XOR U5079 ( .A(n5247), .B(p_input[1451]), .Z(n5249) );
  XOR U5080 ( .A(n5251), .B(n5252), .Z(n5247) );
  AND U5081 ( .A(n5253), .B(n5254), .Z(n5252) );
  XNOR U5082 ( .A(p_input[1466]), .B(n5251), .Z(n5254) );
  XOR U5083 ( .A(n5251), .B(p_input[1450]), .Z(n5253) );
  XOR U5084 ( .A(n5255), .B(n5256), .Z(n5251) );
  AND U5085 ( .A(n5257), .B(n5258), .Z(n5256) );
  XNOR U5086 ( .A(p_input[1465]), .B(n5255), .Z(n5258) );
  XOR U5087 ( .A(n5255), .B(p_input[1449]), .Z(n5257) );
  XOR U5088 ( .A(n5259), .B(n5260), .Z(n5255) );
  AND U5089 ( .A(n5261), .B(n5262), .Z(n5260) );
  XNOR U5090 ( .A(p_input[1464]), .B(n5259), .Z(n5262) );
  XOR U5091 ( .A(n5259), .B(p_input[1448]), .Z(n5261) );
  XOR U5092 ( .A(n5263), .B(n5264), .Z(n5259) );
  AND U5093 ( .A(n5265), .B(n5266), .Z(n5264) );
  XNOR U5094 ( .A(p_input[1463]), .B(n5263), .Z(n5266) );
  XOR U5095 ( .A(n5263), .B(p_input[1447]), .Z(n5265) );
  XOR U5096 ( .A(n5267), .B(n5268), .Z(n5263) );
  AND U5097 ( .A(n5269), .B(n5270), .Z(n5268) );
  XNOR U5098 ( .A(p_input[1462]), .B(n5267), .Z(n5270) );
  XOR U5099 ( .A(n5267), .B(p_input[1446]), .Z(n5269) );
  XOR U5100 ( .A(n5271), .B(n5272), .Z(n5267) );
  AND U5101 ( .A(n5273), .B(n5274), .Z(n5272) );
  XNOR U5102 ( .A(p_input[1461]), .B(n5271), .Z(n5274) );
  XOR U5103 ( .A(n5271), .B(p_input[1445]), .Z(n5273) );
  XOR U5104 ( .A(n5275), .B(n5276), .Z(n5271) );
  AND U5105 ( .A(n5277), .B(n5278), .Z(n5276) );
  XNOR U5106 ( .A(p_input[1460]), .B(n5275), .Z(n5278) );
  XOR U5107 ( .A(n5275), .B(p_input[1444]), .Z(n5277) );
  XOR U5108 ( .A(n5279), .B(n5280), .Z(n5275) );
  AND U5109 ( .A(n5281), .B(n5282), .Z(n5280) );
  XNOR U5110 ( .A(p_input[1459]), .B(n5279), .Z(n5282) );
  XOR U5111 ( .A(n5279), .B(p_input[1443]), .Z(n5281) );
  XOR U5112 ( .A(n5283), .B(n5284), .Z(n5279) );
  AND U5113 ( .A(n5285), .B(n5286), .Z(n5284) );
  XNOR U5114 ( .A(p_input[1458]), .B(n5283), .Z(n5286) );
  XOR U5115 ( .A(n5283), .B(p_input[1442]), .Z(n5285) );
  XNOR U5116 ( .A(n5287), .B(n5288), .Z(n5283) );
  AND U5117 ( .A(n5289), .B(n5290), .Z(n5288) );
  XOR U5118 ( .A(p_input[1457]), .B(n5287), .Z(n5290) );
  XNOR U5119 ( .A(p_input[1441]), .B(n5287), .Z(n5289) );
  AND U5120 ( .A(p_input[1456]), .B(n5291), .Z(n5287) );
  IV U5121 ( .A(p_input[1440]), .Z(n5291) );
  XNOR U5122 ( .A(p_input[1408]), .B(n5292), .Z(n5094) );
  AND U5123 ( .A(n163), .B(n5293), .Z(n5292) );
  XOR U5124 ( .A(p_input[1424]), .B(p_input[1408]), .Z(n5293) );
  XOR U5125 ( .A(n5294), .B(n5295), .Z(n163) );
  AND U5126 ( .A(n5296), .B(n5297), .Z(n5295) );
  XNOR U5127 ( .A(p_input[1439]), .B(n5294), .Z(n5297) );
  XOR U5128 ( .A(n5294), .B(p_input[1423]), .Z(n5296) );
  XOR U5129 ( .A(n5298), .B(n5299), .Z(n5294) );
  AND U5130 ( .A(n5300), .B(n5301), .Z(n5299) );
  XNOR U5131 ( .A(p_input[1438]), .B(n5298), .Z(n5301) );
  XNOR U5132 ( .A(n5298), .B(n5108), .Z(n5300) );
  IV U5133 ( .A(p_input[1422]), .Z(n5108) );
  XOR U5134 ( .A(n5302), .B(n5303), .Z(n5298) );
  AND U5135 ( .A(n5304), .B(n5305), .Z(n5303) );
  XNOR U5136 ( .A(p_input[1437]), .B(n5302), .Z(n5305) );
  XNOR U5137 ( .A(n5302), .B(n5117), .Z(n5304) );
  IV U5138 ( .A(p_input[1421]), .Z(n5117) );
  XOR U5139 ( .A(n5306), .B(n5307), .Z(n5302) );
  AND U5140 ( .A(n5308), .B(n5309), .Z(n5307) );
  XNOR U5141 ( .A(p_input[1436]), .B(n5306), .Z(n5309) );
  XNOR U5142 ( .A(n5306), .B(n5126), .Z(n5308) );
  IV U5143 ( .A(p_input[1420]), .Z(n5126) );
  XOR U5144 ( .A(n5310), .B(n5311), .Z(n5306) );
  AND U5145 ( .A(n5312), .B(n5313), .Z(n5311) );
  XNOR U5146 ( .A(p_input[1435]), .B(n5310), .Z(n5313) );
  XNOR U5147 ( .A(n5310), .B(n5135), .Z(n5312) );
  IV U5148 ( .A(p_input[1419]), .Z(n5135) );
  XOR U5149 ( .A(n5314), .B(n5315), .Z(n5310) );
  AND U5150 ( .A(n5316), .B(n5317), .Z(n5315) );
  XNOR U5151 ( .A(p_input[1434]), .B(n5314), .Z(n5317) );
  XNOR U5152 ( .A(n5314), .B(n5144), .Z(n5316) );
  IV U5153 ( .A(p_input[1418]), .Z(n5144) );
  XOR U5154 ( .A(n5318), .B(n5319), .Z(n5314) );
  AND U5155 ( .A(n5320), .B(n5321), .Z(n5319) );
  XNOR U5156 ( .A(p_input[1433]), .B(n5318), .Z(n5321) );
  XNOR U5157 ( .A(n5318), .B(n5153), .Z(n5320) );
  IV U5158 ( .A(p_input[1417]), .Z(n5153) );
  XOR U5159 ( .A(n5322), .B(n5323), .Z(n5318) );
  AND U5160 ( .A(n5324), .B(n5325), .Z(n5323) );
  XNOR U5161 ( .A(p_input[1432]), .B(n5322), .Z(n5325) );
  XNOR U5162 ( .A(n5322), .B(n5162), .Z(n5324) );
  IV U5163 ( .A(p_input[1416]), .Z(n5162) );
  XOR U5164 ( .A(n5326), .B(n5327), .Z(n5322) );
  AND U5165 ( .A(n5328), .B(n5329), .Z(n5327) );
  XNOR U5166 ( .A(p_input[1431]), .B(n5326), .Z(n5329) );
  XNOR U5167 ( .A(n5326), .B(n5171), .Z(n5328) );
  IV U5168 ( .A(p_input[1415]), .Z(n5171) );
  XOR U5169 ( .A(n5330), .B(n5331), .Z(n5326) );
  AND U5170 ( .A(n5332), .B(n5333), .Z(n5331) );
  XNOR U5171 ( .A(p_input[1430]), .B(n5330), .Z(n5333) );
  XNOR U5172 ( .A(n5330), .B(n5180), .Z(n5332) );
  IV U5173 ( .A(p_input[1414]), .Z(n5180) );
  XOR U5174 ( .A(n5334), .B(n5335), .Z(n5330) );
  AND U5175 ( .A(n5336), .B(n5337), .Z(n5335) );
  XNOR U5176 ( .A(p_input[1429]), .B(n5334), .Z(n5337) );
  XNOR U5177 ( .A(n5334), .B(n5189), .Z(n5336) );
  IV U5178 ( .A(p_input[1413]), .Z(n5189) );
  XOR U5179 ( .A(n5338), .B(n5339), .Z(n5334) );
  AND U5180 ( .A(n5340), .B(n5341), .Z(n5339) );
  XNOR U5181 ( .A(p_input[1428]), .B(n5338), .Z(n5341) );
  XNOR U5182 ( .A(n5338), .B(n5198), .Z(n5340) );
  IV U5183 ( .A(p_input[1412]), .Z(n5198) );
  XOR U5184 ( .A(n5342), .B(n5343), .Z(n5338) );
  AND U5185 ( .A(n5344), .B(n5345), .Z(n5343) );
  XNOR U5186 ( .A(p_input[1427]), .B(n5342), .Z(n5345) );
  XNOR U5187 ( .A(n5342), .B(n5207), .Z(n5344) );
  IV U5188 ( .A(p_input[1411]), .Z(n5207) );
  XOR U5189 ( .A(n5346), .B(n5347), .Z(n5342) );
  AND U5190 ( .A(n5348), .B(n5349), .Z(n5347) );
  XNOR U5191 ( .A(p_input[1426]), .B(n5346), .Z(n5349) );
  XNOR U5192 ( .A(n5346), .B(n5216), .Z(n5348) );
  IV U5193 ( .A(p_input[1410]), .Z(n5216) );
  XNOR U5194 ( .A(n5350), .B(n5351), .Z(n5346) );
  AND U5195 ( .A(n5352), .B(n5353), .Z(n5351) );
  XOR U5196 ( .A(p_input[1425]), .B(n5350), .Z(n5353) );
  XNOR U5197 ( .A(p_input[1409]), .B(n5350), .Z(n5352) );
  AND U5198 ( .A(p_input[1424]), .B(n5354), .Z(n5350) );
  IV U5199 ( .A(p_input[1408]), .Z(n5354) );
  XOR U5200 ( .A(n5355), .B(n5356), .Z(n4470) );
  AND U5201 ( .A(n420), .B(n5357), .Z(n5356) );
  XNOR U5202 ( .A(n5358), .B(n5355), .Z(n5357) );
  XOR U5203 ( .A(n5359), .B(n5360), .Z(n420) );
  AND U5204 ( .A(n5361), .B(n5362), .Z(n5360) );
  XNOR U5205 ( .A(n4482), .B(n5359), .Z(n5362) );
  AND U5206 ( .A(n5363), .B(n5364), .Z(n4482) );
  XOR U5207 ( .A(n5359), .B(n4481), .Z(n5361) );
  AND U5208 ( .A(n5365), .B(n5366), .Z(n4481) );
  XOR U5209 ( .A(n5367), .B(n5368), .Z(n5359) );
  AND U5210 ( .A(n5369), .B(n5370), .Z(n5368) );
  XOR U5211 ( .A(n5367), .B(n4494), .Z(n5370) );
  XOR U5212 ( .A(n5371), .B(n5372), .Z(n4494) );
  AND U5213 ( .A(n258), .B(n5373), .Z(n5372) );
  XOR U5214 ( .A(n5374), .B(n5371), .Z(n5373) );
  XNOR U5215 ( .A(n4491), .B(n5367), .Z(n5369) );
  XOR U5216 ( .A(n5375), .B(n5376), .Z(n4491) );
  AND U5217 ( .A(n255), .B(n5377), .Z(n5376) );
  XOR U5218 ( .A(n5378), .B(n5375), .Z(n5377) );
  XOR U5219 ( .A(n5379), .B(n5380), .Z(n5367) );
  AND U5220 ( .A(n5381), .B(n5382), .Z(n5380) );
  XOR U5221 ( .A(n5379), .B(n4506), .Z(n5382) );
  XOR U5222 ( .A(n5383), .B(n5384), .Z(n4506) );
  AND U5223 ( .A(n258), .B(n5385), .Z(n5384) );
  XOR U5224 ( .A(n5386), .B(n5383), .Z(n5385) );
  XNOR U5225 ( .A(n4503), .B(n5379), .Z(n5381) );
  XOR U5226 ( .A(n5387), .B(n5388), .Z(n4503) );
  AND U5227 ( .A(n255), .B(n5389), .Z(n5388) );
  XOR U5228 ( .A(n5390), .B(n5387), .Z(n5389) );
  XOR U5229 ( .A(n5391), .B(n5392), .Z(n5379) );
  AND U5230 ( .A(n5393), .B(n5394), .Z(n5392) );
  XOR U5231 ( .A(n5391), .B(n4518), .Z(n5394) );
  XOR U5232 ( .A(n5395), .B(n5396), .Z(n4518) );
  AND U5233 ( .A(n258), .B(n5397), .Z(n5396) );
  XOR U5234 ( .A(n5398), .B(n5395), .Z(n5397) );
  XNOR U5235 ( .A(n4515), .B(n5391), .Z(n5393) );
  XOR U5236 ( .A(n5399), .B(n5400), .Z(n4515) );
  AND U5237 ( .A(n255), .B(n5401), .Z(n5400) );
  XOR U5238 ( .A(n5402), .B(n5399), .Z(n5401) );
  XOR U5239 ( .A(n5403), .B(n5404), .Z(n5391) );
  AND U5240 ( .A(n5405), .B(n5406), .Z(n5404) );
  XOR U5241 ( .A(n5403), .B(n4530), .Z(n5406) );
  XOR U5242 ( .A(n5407), .B(n5408), .Z(n4530) );
  AND U5243 ( .A(n258), .B(n5409), .Z(n5408) );
  XOR U5244 ( .A(n5410), .B(n5407), .Z(n5409) );
  XNOR U5245 ( .A(n4527), .B(n5403), .Z(n5405) );
  XOR U5246 ( .A(n5411), .B(n5412), .Z(n4527) );
  AND U5247 ( .A(n255), .B(n5413), .Z(n5412) );
  XOR U5248 ( .A(n5414), .B(n5411), .Z(n5413) );
  XOR U5249 ( .A(n5415), .B(n5416), .Z(n5403) );
  AND U5250 ( .A(n5417), .B(n5418), .Z(n5416) );
  XOR U5251 ( .A(n5415), .B(n4542), .Z(n5418) );
  XOR U5252 ( .A(n5419), .B(n5420), .Z(n4542) );
  AND U5253 ( .A(n258), .B(n5421), .Z(n5420) );
  XOR U5254 ( .A(n5422), .B(n5419), .Z(n5421) );
  XNOR U5255 ( .A(n4539), .B(n5415), .Z(n5417) );
  XOR U5256 ( .A(n5423), .B(n5424), .Z(n4539) );
  AND U5257 ( .A(n255), .B(n5425), .Z(n5424) );
  XOR U5258 ( .A(n5426), .B(n5423), .Z(n5425) );
  XOR U5259 ( .A(n5427), .B(n5428), .Z(n5415) );
  AND U5260 ( .A(n5429), .B(n5430), .Z(n5428) );
  XOR U5261 ( .A(n5427), .B(n4554), .Z(n5430) );
  XOR U5262 ( .A(n5431), .B(n5432), .Z(n4554) );
  AND U5263 ( .A(n258), .B(n5433), .Z(n5432) );
  XOR U5264 ( .A(n5434), .B(n5431), .Z(n5433) );
  XNOR U5265 ( .A(n4551), .B(n5427), .Z(n5429) );
  XOR U5266 ( .A(n5435), .B(n5436), .Z(n4551) );
  AND U5267 ( .A(n255), .B(n5437), .Z(n5436) );
  XOR U5268 ( .A(n5438), .B(n5435), .Z(n5437) );
  XOR U5269 ( .A(n5439), .B(n5440), .Z(n5427) );
  AND U5270 ( .A(n5441), .B(n5442), .Z(n5440) );
  XOR U5271 ( .A(n5439), .B(n4566), .Z(n5442) );
  XOR U5272 ( .A(n5443), .B(n5444), .Z(n4566) );
  AND U5273 ( .A(n258), .B(n5445), .Z(n5444) );
  XOR U5274 ( .A(n5446), .B(n5443), .Z(n5445) );
  XNOR U5275 ( .A(n4563), .B(n5439), .Z(n5441) );
  XOR U5276 ( .A(n5447), .B(n5448), .Z(n4563) );
  AND U5277 ( .A(n255), .B(n5449), .Z(n5448) );
  XOR U5278 ( .A(n5450), .B(n5447), .Z(n5449) );
  XOR U5279 ( .A(n5451), .B(n5452), .Z(n5439) );
  AND U5280 ( .A(n5453), .B(n5454), .Z(n5452) );
  XOR U5281 ( .A(n5451), .B(n4578), .Z(n5454) );
  XOR U5282 ( .A(n5455), .B(n5456), .Z(n4578) );
  AND U5283 ( .A(n258), .B(n5457), .Z(n5456) );
  XOR U5284 ( .A(n5458), .B(n5455), .Z(n5457) );
  XNOR U5285 ( .A(n4575), .B(n5451), .Z(n5453) );
  XOR U5286 ( .A(n5459), .B(n5460), .Z(n4575) );
  AND U5287 ( .A(n255), .B(n5461), .Z(n5460) );
  XOR U5288 ( .A(n5462), .B(n5459), .Z(n5461) );
  XOR U5289 ( .A(n5463), .B(n5464), .Z(n5451) );
  AND U5290 ( .A(n5465), .B(n5466), .Z(n5464) );
  XOR U5291 ( .A(n5463), .B(n4590), .Z(n5466) );
  XOR U5292 ( .A(n5467), .B(n5468), .Z(n4590) );
  AND U5293 ( .A(n258), .B(n5469), .Z(n5468) );
  XOR U5294 ( .A(n5470), .B(n5467), .Z(n5469) );
  XNOR U5295 ( .A(n4587), .B(n5463), .Z(n5465) );
  XOR U5296 ( .A(n5471), .B(n5472), .Z(n4587) );
  AND U5297 ( .A(n255), .B(n5473), .Z(n5472) );
  XOR U5298 ( .A(n5474), .B(n5471), .Z(n5473) );
  XOR U5299 ( .A(n5475), .B(n5476), .Z(n5463) );
  AND U5300 ( .A(n5477), .B(n5478), .Z(n5476) );
  XOR U5301 ( .A(n5475), .B(n4602), .Z(n5478) );
  XOR U5302 ( .A(n5479), .B(n5480), .Z(n4602) );
  AND U5303 ( .A(n258), .B(n5481), .Z(n5480) );
  XOR U5304 ( .A(n5482), .B(n5479), .Z(n5481) );
  XNOR U5305 ( .A(n4599), .B(n5475), .Z(n5477) );
  XOR U5306 ( .A(n5483), .B(n5484), .Z(n4599) );
  AND U5307 ( .A(n255), .B(n5485), .Z(n5484) );
  XOR U5308 ( .A(n5486), .B(n5483), .Z(n5485) );
  XOR U5309 ( .A(n5487), .B(n5488), .Z(n5475) );
  AND U5310 ( .A(n5489), .B(n5490), .Z(n5488) );
  XOR U5311 ( .A(n5487), .B(n4614), .Z(n5490) );
  XOR U5312 ( .A(n5491), .B(n5492), .Z(n4614) );
  AND U5313 ( .A(n258), .B(n5493), .Z(n5492) );
  XOR U5314 ( .A(n5494), .B(n5491), .Z(n5493) );
  XNOR U5315 ( .A(n4611), .B(n5487), .Z(n5489) );
  XOR U5316 ( .A(n5495), .B(n5496), .Z(n4611) );
  AND U5317 ( .A(n255), .B(n5497), .Z(n5496) );
  XOR U5318 ( .A(n5498), .B(n5495), .Z(n5497) );
  XOR U5319 ( .A(n5499), .B(n5500), .Z(n5487) );
  AND U5320 ( .A(n5501), .B(n5502), .Z(n5500) );
  XOR U5321 ( .A(n5499), .B(n4626), .Z(n5502) );
  XOR U5322 ( .A(n5503), .B(n5504), .Z(n4626) );
  AND U5323 ( .A(n258), .B(n5505), .Z(n5504) );
  XOR U5324 ( .A(n5506), .B(n5503), .Z(n5505) );
  XNOR U5325 ( .A(n4623), .B(n5499), .Z(n5501) );
  XOR U5326 ( .A(n5507), .B(n5508), .Z(n4623) );
  AND U5327 ( .A(n255), .B(n5509), .Z(n5508) );
  XOR U5328 ( .A(n5510), .B(n5507), .Z(n5509) );
  XOR U5329 ( .A(n5511), .B(n5512), .Z(n5499) );
  AND U5330 ( .A(n5513), .B(n5514), .Z(n5512) );
  XOR U5331 ( .A(n4638), .B(n5511), .Z(n5514) );
  XOR U5332 ( .A(n5515), .B(n5516), .Z(n4638) );
  AND U5333 ( .A(n258), .B(n5517), .Z(n5516) );
  XOR U5334 ( .A(n5515), .B(n5518), .Z(n5517) );
  XNOR U5335 ( .A(n5511), .B(n4635), .Z(n5513) );
  XOR U5336 ( .A(n5519), .B(n5520), .Z(n4635) );
  AND U5337 ( .A(n255), .B(n5521), .Z(n5520) );
  XOR U5338 ( .A(n5519), .B(n5522), .Z(n5521) );
  XOR U5339 ( .A(n5523), .B(n5524), .Z(n5511) );
  AND U5340 ( .A(n5525), .B(n5526), .Z(n5524) );
  XNOR U5341 ( .A(n5527), .B(n4651), .Z(n5526) );
  XOR U5342 ( .A(n5528), .B(n5529), .Z(n4651) );
  AND U5343 ( .A(n258), .B(n5530), .Z(n5529) );
  XOR U5344 ( .A(n5531), .B(n5528), .Z(n5530) );
  XNOR U5345 ( .A(n4648), .B(n5523), .Z(n5525) );
  XOR U5346 ( .A(n5532), .B(n5533), .Z(n4648) );
  AND U5347 ( .A(n255), .B(n5534), .Z(n5533) );
  XOR U5348 ( .A(n5535), .B(n5532), .Z(n5534) );
  IV U5349 ( .A(n5527), .Z(n5523) );
  AND U5350 ( .A(n5355), .B(n5358), .Z(n5527) );
  XNOR U5351 ( .A(n5536), .B(n5537), .Z(n5358) );
  AND U5352 ( .A(n258), .B(n5538), .Z(n5537) );
  XNOR U5353 ( .A(n5539), .B(n5536), .Z(n5538) );
  XOR U5354 ( .A(n5540), .B(n5541), .Z(n258) );
  AND U5355 ( .A(n5542), .B(n5543), .Z(n5541) );
  XNOR U5356 ( .A(n5363), .B(n5540), .Z(n5543) );
  AND U5357 ( .A(p_input[1407]), .B(p_input[1391]), .Z(n5363) );
  XOR U5358 ( .A(n5540), .B(n5364), .Z(n5542) );
  AND U5359 ( .A(p_input[1375]), .B(p_input[1359]), .Z(n5364) );
  XOR U5360 ( .A(n5544), .B(n5545), .Z(n5540) );
  AND U5361 ( .A(n5546), .B(n5547), .Z(n5545) );
  XOR U5362 ( .A(n5544), .B(n5374), .Z(n5547) );
  XNOR U5363 ( .A(p_input[1390]), .B(n5548), .Z(n5374) );
  AND U5364 ( .A(n174), .B(n5549), .Z(n5548) );
  XOR U5365 ( .A(p_input[1406]), .B(p_input[1390]), .Z(n5549) );
  XNOR U5366 ( .A(n5371), .B(n5544), .Z(n5546) );
  XOR U5367 ( .A(n5550), .B(n5551), .Z(n5371) );
  AND U5368 ( .A(n172), .B(n5552), .Z(n5551) );
  XOR U5369 ( .A(p_input[1374]), .B(p_input[1358]), .Z(n5552) );
  XOR U5370 ( .A(n5553), .B(n5554), .Z(n5544) );
  AND U5371 ( .A(n5555), .B(n5556), .Z(n5554) );
  XOR U5372 ( .A(n5553), .B(n5386), .Z(n5556) );
  XNOR U5373 ( .A(p_input[1389]), .B(n5557), .Z(n5386) );
  AND U5374 ( .A(n174), .B(n5558), .Z(n5557) );
  XOR U5375 ( .A(p_input[1405]), .B(p_input[1389]), .Z(n5558) );
  XNOR U5376 ( .A(n5383), .B(n5553), .Z(n5555) );
  XOR U5377 ( .A(n5559), .B(n5560), .Z(n5383) );
  AND U5378 ( .A(n172), .B(n5561), .Z(n5560) );
  XOR U5379 ( .A(p_input[1373]), .B(p_input[1357]), .Z(n5561) );
  XOR U5380 ( .A(n5562), .B(n5563), .Z(n5553) );
  AND U5381 ( .A(n5564), .B(n5565), .Z(n5563) );
  XOR U5382 ( .A(n5562), .B(n5398), .Z(n5565) );
  XNOR U5383 ( .A(p_input[1388]), .B(n5566), .Z(n5398) );
  AND U5384 ( .A(n174), .B(n5567), .Z(n5566) );
  XOR U5385 ( .A(p_input[1404]), .B(p_input[1388]), .Z(n5567) );
  XNOR U5386 ( .A(n5395), .B(n5562), .Z(n5564) );
  XOR U5387 ( .A(n5568), .B(n5569), .Z(n5395) );
  AND U5388 ( .A(n172), .B(n5570), .Z(n5569) );
  XOR U5389 ( .A(p_input[1372]), .B(p_input[1356]), .Z(n5570) );
  XOR U5390 ( .A(n5571), .B(n5572), .Z(n5562) );
  AND U5391 ( .A(n5573), .B(n5574), .Z(n5572) );
  XOR U5392 ( .A(n5571), .B(n5410), .Z(n5574) );
  XNOR U5393 ( .A(p_input[1387]), .B(n5575), .Z(n5410) );
  AND U5394 ( .A(n174), .B(n5576), .Z(n5575) );
  XOR U5395 ( .A(p_input[1403]), .B(p_input[1387]), .Z(n5576) );
  XNOR U5396 ( .A(n5407), .B(n5571), .Z(n5573) );
  XOR U5397 ( .A(n5577), .B(n5578), .Z(n5407) );
  AND U5398 ( .A(n172), .B(n5579), .Z(n5578) );
  XOR U5399 ( .A(p_input[1371]), .B(p_input[1355]), .Z(n5579) );
  XOR U5400 ( .A(n5580), .B(n5581), .Z(n5571) );
  AND U5401 ( .A(n5582), .B(n5583), .Z(n5581) );
  XOR U5402 ( .A(n5580), .B(n5422), .Z(n5583) );
  XNOR U5403 ( .A(p_input[1386]), .B(n5584), .Z(n5422) );
  AND U5404 ( .A(n174), .B(n5585), .Z(n5584) );
  XOR U5405 ( .A(p_input[1402]), .B(p_input[1386]), .Z(n5585) );
  XNOR U5406 ( .A(n5419), .B(n5580), .Z(n5582) );
  XOR U5407 ( .A(n5586), .B(n5587), .Z(n5419) );
  AND U5408 ( .A(n172), .B(n5588), .Z(n5587) );
  XOR U5409 ( .A(p_input[1370]), .B(p_input[1354]), .Z(n5588) );
  XOR U5410 ( .A(n5589), .B(n5590), .Z(n5580) );
  AND U5411 ( .A(n5591), .B(n5592), .Z(n5590) );
  XOR U5412 ( .A(n5589), .B(n5434), .Z(n5592) );
  XNOR U5413 ( .A(p_input[1385]), .B(n5593), .Z(n5434) );
  AND U5414 ( .A(n174), .B(n5594), .Z(n5593) );
  XOR U5415 ( .A(p_input[1401]), .B(p_input[1385]), .Z(n5594) );
  XNOR U5416 ( .A(n5431), .B(n5589), .Z(n5591) );
  XOR U5417 ( .A(n5595), .B(n5596), .Z(n5431) );
  AND U5418 ( .A(n172), .B(n5597), .Z(n5596) );
  XOR U5419 ( .A(p_input[1369]), .B(p_input[1353]), .Z(n5597) );
  XOR U5420 ( .A(n5598), .B(n5599), .Z(n5589) );
  AND U5421 ( .A(n5600), .B(n5601), .Z(n5599) );
  XOR U5422 ( .A(n5598), .B(n5446), .Z(n5601) );
  XNOR U5423 ( .A(p_input[1384]), .B(n5602), .Z(n5446) );
  AND U5424 ( .A(n174), .B(n5603), .Z(n5602) );
  XOR U5425 ( .A(p_input[1400]), .B(p_input[1384]), .Z(n5603) );
  XNOR U5426 ( .A(n5443), .B(n5598), .Z(n5600) );
  XOR U5427 ( .A(n5604), .B(n5605), .Z(n5443) );
  AND U5428 ( .A(n172), .B(n5606), .Z(n5605) );
  XOR U5429 ( .A(p_input[1368]), .B(p_input[1352]), .Z(n5606) );
  XOR U5430 ( .A(n5607), .B(n5608), .Z(n5598) );
  AND U5431 ( .A(n5609), .B(n5610), .Z(n5608) );
  XOR U5432 ( .A(n5607), .B(n5458), .Z(n5610) );
  XNOR U5433 ( .A(p_input[1383]), .B(n5611), .Z(n5458) );
  AND U5434 ( .A(n174), .B(n5612), .Z(n5611) );
  XOR U5435 ( .A(p_input[1399]), .B(p_input[1383]), .Z(n5612) );
  XNOR U5436 ( .A(n5455), .B(n5607), .Z(n5609) );
  XOR U5437 ( .A(n5613), .B(n5614), .Z(n5455) );
  AND U5438 ( .A(n172), .B(n5615), .Z(n5614) );
  XOR U5439 ( .A(p_input[1367]), .B(p_input[1351]), .Z(n5615) );
  XOR U5440 ( .A(n5616), .B(n5617), .Z(n5607) );
  AND U5441 ( .A(n5618), .B(n5619), .Z(n5617) );
  XOR U5442 ( .A(n5616), .B(n5470), .Z(n5619) );
  XNOR U5443 ( .A(p_input[1382]), .B(n5620), .Z(n5470) );
  AND U5444 ( .A(n174), .B(n5621), .Z(n5620) );
  XOR U5445 ( .A(p_input[1398]), .B(p_input[1382]), .Z(n5621) );
  XNOR U5446 ( .A(n5467), .B(n5616), .Z(n5618) );
  XOR U5447 ( .A(n5622), .B(n5623), .Z(n5467) );
  AND U5448 ( .A(n172), .B(n5624), .Z(n5623) );
  XOR U5449 ( .A(p_input[1366]), .B(p_input[1350]), .Z(n5624) );
  XOR U5450 ( .A(n5625), .B(n5626), .Z(n5616) );
  AND U5451 ( .A(n5627), .B(n5628), .Z(n5626) );
  XOR U5452 ( .A(n5625), .B(n5482), .Z(n5628) );
  XNOR U5453 ( .A(p_input[1381]), .B(n5629), .Z(n5482) );
  AND U5454 ( .A(n174), .B(n5630), .Z(n5629) );
  XOR U5455 ( .A(p_input[1397]), .B(p_input[1381]), .Z(n5630) );
  XNOR U5456 ( .A(n5479), .B(n5625), .Z(n5627) );
  XOR U5457 ( .A(n5631), .B(n5632), .Z(n5479) );
  AND U5458 ( .A(n172), .B(n5633), .Z(n5632) );
  XOR U5459 ( .A(p_input[1365]), .B(p_input[1349]), .Z(n5633) );
  XOR U5460 ( .A(n5634), .B(n5635), .Z(n5625) );
  AND U5461 ( .A(n5636), .B(n5637), .Z(n5635) );
  XOR U5462 ( .A(n5634), .B(n5494), .Z(n5637) );
  XNOR U5463 ( .A(p_input[1380]), .B(n5638), .Z(n5494) );
  AND U5464 ( .A(n174), .B(n5639), .Z(n5638) );
  XOR U5465 ( .A(p_input[1396]), .B(p_input[1380]), .Z(n5639) );
  XNOR U5466 ( .A(n5491), .B(n5634), .Z(n5636) );
  XOR U5467 ( .A(n5640), .B(n5641), .Z(n5491) );
  AND U5468 ( .A(n172), .B(n5642), .Z(n5641) );
  XOR U5469 ( .A(p_input[1364]), .B(p_input[1348]), .Z(n5642) );
  XOR U5470 ( .A(n5643), .B(n5644), .Z(n5634) );
  AND U5471 ( .A(n5645), .B(n5646), .Z(n5644) );
  XOR U5472 ( .A(n5643), .B(n5506), .Z(n5646) );
  XNOR U5473 ( .A(p_input[1379]), .B(n5647), .Z(n5506) );
  AND U5474 ( .A(n174), .B(n5648), .Z(n5647) );
  XOR U5475 ( .A(p_input[1395]), .B(p_input[1379]), .Z(n5648) );
  XNOR U5476 ( .A(n5503), .B(n5643), .Z(n5645) );
  XOR U5477 ( .A(n5649), .B(n5650), .Z(n5503) );
  AND U5478 ( .A(n172), .B(n5651), .Z(n5650) );
  XOR U5479 ( .A(p_input[1363]), .B(p_input[1347]), .Z(n5651) );
  XOR U5480 ( .A(n5652), .B(n5653), .Z(n5643) );
  AND U5481 ( .A(n5654), .B(n5655), .Z(n5653) );
  XOR U5482 ( .A(n5518), .B(n5652), .Z(n5655) );
  XNOR U5483 ( .A(p_input[1378]), .B(n5656), .Z(n5518) );
  AND U5484 ( .A(n174), .B(n5657), .Z(n5656) );
  XOR U5485 ( .A(p_input[1394]), .B(p_input[1378]), .Z(n5657) );
  XNOR U5486 ( .A(n5652), .B(n5515), .Z(n5654) );
  XOR U5487 ( .A(n5658), .B(n5659), .Z(n5515) );
  AND U5488 ( .A(n172), .B(n5660), .Z(n5659) );
  XOR U5489 ( .A(p_input[1362]), .B(p_input[1346]), .Z(n5660) );
  XOR U5490 ( .A(n5661), .B(n5662), .Z(n5652) );
  AND U5491 ( .A(n5663), .B(n5664), .Z(n5662) );
  XNOR U5492 ( .A(n5665), .B(n5531), .Z(n5664) );
  XNOR U5493 ( .A(p_input[1377]), .B(n5666), .Z(n5531) );
  AND U5494 ( .A(n174), .B(n5667), .Z(n5666) );
  XNOR U5495 ( .A(p_input[1393]), .B(n5668), .Z(n5667) );
  IV U5496 ( .A(p_input[1377]), .Z(n5668) );
  XNOR U5497 ( .A(n5528), .B(n5661), .Z(n5663) );
  XNOR U5498 ( .A(p_input[1345]), .B(n5669), .Z(n5528) );
  AND U5499 ( .A(n172), .B(n5670), .Z(n5669) );
  XOR U5500 ( .A(p_input[1361]), .B(p_input[1345]), .Z(n5670) );
  IV U5501 ( .A(n5665), .Z(n5661) );
  AND U5502 ( .A(n5536), .B(n5539), .Z(n5665) );
  XOR U5503 ( .A(p_input[1376]), .B(n5671), .Z(n5539) );
  AND U5504 ( .A(n174), .B(n5672), .Z(n5671) );
  XOR U5505 ( .A(p_input[1392]), .B(p_input[1376]), .Z(n5672) );
  XOR U5506 ( .A(n5673), .B(n5674), .Z(n174) );
  AND U5507 ( .A(n5675), .B(n5676), .Z(n5674) );
  XNOR U5508 ( .A(p_input[1407]), .B(n5673), .Z(n5676) );
  XOR U5509 ( .A(n5673), .B(p_input[1391]), .Z(n5675) );
  XOR U5510 ( .A(n5677), .B(n5678), .Z(n5673) );
  AND U5511 ( .A(n5679), .B(n5680), .Z(n5678) );
  XNOR U5512 ( .A(p_input[1406]), .B(n5677), .Z(n5680) );
  XOR U5513 ( .A(n5677), .B(p_input[1390]), .Z(n5679) );
  XOR U5514 ( .A(n5681), .B(n5682), .Z(n5677) );
  AND U5515 ( .A(n5683), .B(n5684), .Z(n5682) );
  XNOR U5516 ( .A(p_input[1405]), .B(n5681), .Z(n5684) );
  XOR U5517 ( .A(n5681), .B(p_input[1389]), .Z(n5683) );
  XOR U5518 ( .A(n5685), .B(n5686), .Z(n5681) );
  AND U5519 ( .A(n5687), .B(n5688), .Z(n5686) );
  XNOR U5520 ( .A(p_input[1404]), .B(n5685), .Z(n5688) );
  XOR U5521 ( .A(n5685), .B(p_input[1388]), .Z(n5687) );
  XOR U5522 ( .A(n5689), .B(n5690), .Z(n5685) );
  AND U5523 ( .A(n5691), .B(n5692), .Z(n5690) );
  XNOR U5524 ( .A(p_input[1403]), .B(n5689), .Z(n5692) );
  XOR U5525 ( .A(n5689), .B(p_input[1387]), .Z(n5691) );
  XOR U5526 ( .A(n5693), .B(n5694), .Z(n5689) );
  AND U5527 ( .A(n5695), .B(n5696), .Z(n5694) );
  XNOR U5528 ( .A(p_input[1402]), .B(n5693), .Z(n5696) );
  XOR U5529 ( .A(n5693), .B(p_input[1386]), .Z(n5695) );
  XOR U5530 ( .A(n5697), .B(n5698), .Z(n5693) );
  AND U5531 ( .A(n5699), .B(n5700), .Z(n5698) );
  XNOR U5532 ( .A(p_input[1401]), .B(n5697), .Z(n5700) );
  XOR U5533 ( .A(n5697), .B(p_input[1385]), .Z(n5699) );
  XOR U5534 ( .A(n5701), .B(n5702), .Z(n5697) );
  AND U5535 ( .A(n5703), .B(n5704), .Z(n5702) );
  XNOR U5536 ( .A(p_input[1400]), .B(n5701), .Z(n5704) );
  XOR U5537 ( .A(n5701), .B(p_input[1384]), .Z(n5703) );
  XOR U5538 ( .A(n5705), .B(n5706), .Z(n5701) );
  AND U5539 ( .A(n5707), .B(n5708), .Z(n5706) );
  XNOR U5540 ( .A(p_input[1399]), .B(n5705), .Z(n5708) );
  XOR U5541 ( .A(n5705), .B(p_input[1383]), .Z(n5707) );
  XOR U5542 ( .A(n5709), .B(n5710), .Z(n5705) );
  AND U5543 ( .A(n5711), .B(n5712), .Z(n5710) );
  XNOR U5544 ( .A(p_input[1398]), .B(n5709), .Z(n5712) );
  XOR U5545 ( .A(n5709), .B(p_input[1382]), .Z(n5711) );
  XOR U5546 ( .A(n5713), .B(n5714), .Z(n5709) );
  AND U5547 ( .A(n5715), .B(n5716), .Z(n5714) );
  XNOR U5548 ( .A(p_input[1397]), .B(n5713), .Z(n5716) );
  XOR U5549 ( .A(n5713), .B(p_input[1381]), .Z(n5715) );
  XOR U5550 ( .A(n5717), .B(n5718), .Z(n5713) );
  AND U5551 ( .A(n5719), .B(n5720), .Z(n5718) );
  XNOR U5552 ( .A(p_input[1396]), .B(n5717), .Z(n5720) );
  XOR U5553 ( .A(n5717), .B(p_input[1380]), .Z(n5719) );
  XOR U5554 ( .A(n5721), .B(n5722), .Z(n5717) );
  AND U5555 ( .A(n5723), .B(n5724), .Z(n5722) );
  XNOR U5556 ( .A(p_input[1395]), .B(n5721), .Z(n5724) );
  XOR U5557 ( .A(n5721), .B(p_input[1379]), .Z(n5723) );
  XOR U5558 ( .A(n5725), .B(n5726), .Z(n5721) );
  AND U5559 ( .A(n5727), .B(n5728), .Z(n5726) );
  XNOR U5560 ( .A(p_input[1394]), .B(n5725), .Z(n5728) );
  XOR U5561 ( .A(n5725), .B(p_input[1378]), .Z(n5727) );
  XNOR U5562 ( .A(n5729), .B(n5730), .Z(n5725) );
  AND U5563 ( .A(n5731), .B(n5732), .Z(n5730) );
  XOR U5564 ( .A(p_input[1393]), .B(n5729), .Z(n5732) );
  XNOR U5565 ( .A(p_input[1377]), .B(n5729), .Z(n5731) );
  AND U5566 ( .A(p_input[1392]), .B(n5733), .Z(n5729) );
  IV U5567 ( .A(p_input[1376]), .Z(n5733) );
  XNOR U5568 ( .A(p_input[1344]), .B(n5734), .Z(n5536) );
  AND U5569 ( .A(n172), .B(n5735), .Z(n5734) );
  XOR U5570 ( .A(p_input[1360]), .B(p_input[1344]), .Z(n5735) );
  XOR U5571 ( .A(n5736), .B(n5737), .Z(n172) );
  AND U5572 ( .A(n5738), .B(n5739), .Z(n5737) );
  XNOR U5573 ( .A(p_input[1375]), .B(n5736), .Z(n5739) );
  XOR U5574 ( .A(n5736), .B(p_input[1359]), .Z(n5738) );
  XOR U5575 ( .A(n5740), .B(n5741), .Z(n5736) );
  AND U5576 ( .A(n5742), .B(n5743), .Z(n5741) );
  XNOR U5577 ( .A(p_input[1374]), .B(n5740), .Z(n5743) );
  XNOR U5578 ( .A(n5740), .B(n5550), .Z(n5742) );
  IV U5579 ( .A(p_input[1358]), .Z(n5550) );
  XOR U5580 ( .A(n5744), .B(n5745), .Z(n5740) );
  AND U5581 ( .A(n5746), .B(n5747), .Z(n5745) );
  XNOR U5582 ( .A(p_input[1373]), .B(n5744), .Z(n5747) );
  XNOR U5583 ( .A(n5744), .B(n5559), .Z(n5746) );
  IV U5584 ( .A(p_input[1357]), .Z(n5559) );
  XOR U5585 ( .A(n5748), .B(n5749), .Z(n5744) );
  AND U5586 ( .A(n5750), .B(n5751), .Z(n5749) );
  XNOR U5587 ( .A(p_input[1372]), .B(n5748), .Z(n5751) );
  XNOR U5588 ( .A(n5748), .B(n5568), .Z(n5750) );
  IV U5589 ( .A(p_input[1356]), .Z(n5568) );
  XOR U5590 ( .A(n5752), .B(n5753), .Z(n5748) );
  AND U5591 ( .A(n5754), .B(n5755), .Z(n5753) );
  XNOR U5592 ( .A(p_input[1371]), .B(n5752), .Z(n5755) );
  XNOR U5593 ( .A(n5752), .B(n5577), .Z(n5754) );
  IV U5594 ( .A(p_input[1355]), .Z(n5577) );
  XOR U5595 ( .A(n5756), .B(n5757), .Z(n5752) );
  AND U5596 ( .A(n5758), .B(n5759), .Z(n5757) );
  XNOR U5597 ( .A(p_input[1370]), .B(n5756), .Z(n5759) );
  XNOR U5598 ( .A(n5756), .B(n5586), .Z(n5758) );
  IV U5599 ( .A(p_input[1354]), .Z(n5586) );
  XOR U5600 ( .A(n5760), .B(n5761), .Z(n5756) );
  AND U5601 ( .A(n5762), .B(n5763), .Z(n5761) );
  XNOR U5602 ( .A(p_input[1369]), .B(n5760), .Z(n5763) );
  XNOR U5603 ( .A(n5760), .B(n5595), .Z(n5762) );
  IV U5604 ( .A(p_input[1353]), .Z(n5595) );
  XOR U5605 ( .A(n5764), .B(n5765), .Z(n5760) );
  AND U5606 ( .A(n5766), .B(n5767), .Z(n5765) );
  XNOR U5607 ( .A(p_input[1368]), .B(n5764), .Z(n5767) );
  XNOR U5608 ( .A(n5764), .B(n5604), .Z(n5766) );
  IV U5609 ( .A(p_input[1352]), .Z(n5604) );
  XOR U5610 ( .A(n5768), .B(n5769), .Z(n5764) );
  AND U5611 ( .A(n5770), .B(n5771), .Z(n5769) );
  XNOR U5612 ( .A(p_input[1367]), .B(n5768), .Z(n5771) );
  XNOR U5613 ( .A(n5768), .B(n5613), .Z(n5770) );
  IV U5614 ( .A(p_input[1351]), .Z(n5613) );
  XOR U5615 ( .A(n5772), .B(n5773), .Z(n5768) );
  AND U5616 ( .A(n5774), .B(n5775), .Z(n5773) );
  XNOR U5617 ( .A(p_input[1366]), .B(n5772), .Z(n5775) );
  XNOR U5618 ( .A(n5772), .B(n5622), .Z(n5774) );
  IV U5619 ( .A(p_input[1350]), .Z(n5622) );
  XOR U5620 ( .A(n5776), .B(n5777), .Z(n5772) );
  AND U5621 ( .A(n5778), .B(n5779), .Z(n5777) );
  XNOR U5622 ( .A(p_input[1365]), .B(n5776), .Z(n5779) );
  XNOR U5623 ( .A(n5776), .B(n5631), .Z(n5778) );
  IV U5624 ( .A(p_input[1349]), .Z(n5631) );
  XOR U5625 ( .A(n5780), .B(n5781), .Z(n5776) );
  AND U5626 ( .A(n5782), .B(n5783), .Z(n5781) );
  XNOR U5627 ( .A(p_input[1364]), .B(n5780), .Z(n5783) );
  XNOR U5628 ( .A(n5780), .B(n5640), .Z(n5782) );
  IV U5629 ( .A(p_input[1348]), .Z(n5640) );
  XOR U5630 ( .A(n5784), .B(n5785), .Z(n5780) );
  AND U5631 ( .A(n5786), .B(n5787), .Z(n5785) );
  XNOR U5632 ( .A(p_input[1363]), .B(n5784), .Z(n5787) );
  XNOR U5633 ( .A(n5784), .B(n5649), .Z(n5786) );
  IV U5634 ( .A(p_input[1347]), .Z(n5649) );
  XOR U5635 ( .A(n5788), .B(n5789), .Z(n5784) );
  AND U5636 ( .A(n5790), .B(n5791), .Z(n5789) );
  XNOR U5637 ( .A(p_input[1362]), .B(n5788), .Z(n5791) );
  XNOR U5638 ( .A(n5788), .B(n5658), .Z(n5790) );
  IV U5639 ( .A(p_input[1346]), .Z(n5658) );
  XNOR U5640 ( .A(n5792), .B(n5793), .Z(n5788) );
  AND U5641 ( .A(n5794), .B(n5795), .Z(n5793) );
  XOR U5642 ( .A(p_input[1361]), .B(n5792), .Z(n5795) );
  XNOR U5643 ( .A(p_input[1345]), .B(n5792), .Z(n5794) );
  AND U5644 ( .A(p_input[1360]), .B(n5796), .Z(n5792) );
  IV U5645 ( .A(p_input[1344]), .Z(n5796) );
  XOR U5646 ( .A(n5797), .B(n5798), .Z(n5355) );
  AND U5647 ( .A(n255), .B(n5799), .Z(n5798) );
  XNOR U5648 ( .A(n5800), .B(n5797), .Z(n5799) );
  XOR U5649 ( .A(n5801), .B(n5802), .Z(n255) );
  AND U5650 ( .A(n5803), .B(n5804), .Z(n5802) );
  XNOR U5651 ( .A(n5366), .B(n5801), .Z(n5804) );
  AND U5652 ( .A(p_input[1343]), .B(p_input[1327]), .Z(n5366) );
  XOR U5653 ( .A(n5801), .B(n5365), .Z(n5803) );
  AND U5654 ( .A(p_input[1295]), .B(p_input[1311]), .Z(n5365) );
  XOR U5655 ( .A(n5805), .B(n5806), .Z(n5801) );
  AND U5656 ( .A(n5807), .B(n5808), .Z(n5806) );
  XOR U5657 ( .A(n5805), .B(n5378), .Z(n5808) );
  XNOR U5658 ( .A(p_input[1326]), .B(n5809), .Z(n5378) );
  AND U5659 ( .A(n178), .B(n5810), .Z(n5809) );
  XOR U5660 ( .A(p_input[1342]), .B(p_input[1326]), .Z(n5810) );
  XNOR U5661 ( .A(n5375), .B(n5805), .Z(n5807) );
  XOR U5662 ( .A(n5811), .B(n5812), .Z(n5375) );
  AND U5663 ( .A(n175), .B(n5813), .Z(n5812) );
  XOR U5664 ( .A(p_input[1310]), .B(p_input[1294]), .Z(n5813) );
  XOR U5665 ( .A(n5814), .B(n5815), .Z(n5805) );
  AND U5666 ( .A(n5816), .B(n5817), .Z(n5815) );
  XOR U5667 ( .A(n5814), .B(n5390), .Z(n5817) );
  XNOR U5668 ( .A(p_input[1325]), .B(n5818), .Z(n5390) );
  AND U5669 ( .A(n178), .B(n5819), .Z(n5818) );
  XOR U5670 ( .A(p_input[1341]), .B(p_input[1325]), .Z(n5819) );
  XNOR U5671 ( .A(n5387), .B(n5814), .Z(n5816) );
  XOR U5672 ( .A(n5820), .B(n5821), .Z(n5387) );
  AND U5673 ( .A(n175), .B(n5822), .Z(n5821) );
  XOR U5674 ( .A(p_input[1309]), .B(p_input[1293]), .Z(n5822) );
  XOR U5675 ( .A(n5823), .B(n5824), .Z(n5814) );
  AND U5676 ( .A(n5825), .B(n5826), .Z(n5824) );
  XOR U5677 ( .A(n5823), .B(n5402), .Z(n5826) );
  XNOR U5678 ( .A(p_input[1324]), .B(n5827), .Z(n5402) );
  AND U5679 ( .A(n178), .B(n5828), .Z(n5827) );
  XOR U5680 ( .A(p_input[1340]), .B(p_input[1324]), .Z(n5828) );
  XNOR U5681 ( .A(n5399), .B(n5823), .Z(n5825) );
  XOR U5682 ( .A(n5829), .B(n5830), .Z(n5399) );
  AND U5683 ( .A(n175), .B(n5831), .Z(n5830) );
  XOR U5684 ( .A(p_input[1308]), .B(p_input[1292]), .Z(n5831) );
  XOR U5685 ( .A(n5832), .B(n5833), .Z(n5823) );
  AND U5686 ( .A(n5834), .B(n5835), .Z(n5833) );
  XOR U5687 ( .A(n5832), .B(n5414), .Z(n5835) );
  XNOR U5688 ( .A(p_input[1323]), .B(n5836), .Z(n5414) );
  AND U5689 ( .A(n178), .B(n5837), .Z(n5836) );
  XOR U5690 ( .A(p_input[1339]), .B(p_input[1323]), .Z(n5837) );
  XNOR U5691 ( .A(n5411), .B(n5832), .Z(n5834) );
  XOR U5692 ( .A(n5838), .B(n5839), .Z(n5411) );
  AND U5693 ( .A(n175), .B(n5840), .Z(n5839) );
  XOR U5694 ( .A(p_input[1307]), .B(p_input[1291]), .Z(n5840) );
  XOR U5695 ( .A(n5841), .B(n5842), .Z(n5832) );
  AND U5696 ( .A(n5843), .B(n5844), .Z(n5842) );
  XOR U5697 ( .A(n5841), .B(n5426), .Z(n5844) );
  XNOR U5698 ( .A(p_input[1322]), .B(n5845), .Z(n5426) );
  AND U5699 ( .A(n178), .B(n5846), .Z(n5845) );
  XOR U5700 ( .A(p_input[1338]), .B(p_input[1322]), .Z(n5846) );
  XNOR U5701 ( .A(n5423), .B(n5841), .Z(n5843) );
  XOR U5702 ( .A(n5847), .B(n5848), .Z(n5423) );
  AND U5703 ( .A(n175), .B(n5849), .Z(n5848) );
  XOR U5704 ( .A(p_input[1306]), .B(p_input[1290]), .Z(n5849) );
  XOR U5705 ( .A(n5850), .B(n5851), .Z(n5841) );
  AND U5706 ( .A(n5852), .B(n5853), .Z(n5851) );
  XOR U5707 ( .A(n5850), .B(n5438), .Z(n5853) );
  XNOR U5708 ( .A(p_input[1321]), .B(n5854), .Z(n5438) );
  AND U5709 ( .A(n178), .B(n5855), .Z(n5854) );
  XOR U5710 ( .A(p_input[1337]), .B(p_input[1321]), .Z(n5855) );
  XNOR U5711 ( .A(n5435), .B(n5850), .Z(n5852) );
  XOR U5712 ( .A(n5856), .B(n5857), .Z(n5435) );
  AND U5713 ( .A(n175), .B(n5858), .Z(n5857) );
  XOR U5714 ( .A(p_input[1305]), .B(p_input[1289]), .Z(n5858) );
  XOR U5715 ( .A(n5859), .B(n5860), .Z(n5850) );
  AND U5716 ( .A(n5861), .B(n5862), .Z(n5860) );
  XOR U5717 ( .A(n5859), .B(n5450), .Z(n5862) );
  XNOR U5718 ( .A(p_input[1320]), .B(n5863), .Z(n5450) );
  AND U5719 ( .A(n178), .B(n5864), .Z(n5863) );
  XOR U5720 ( .A(p_input[1336]), .B(p_input[1320]), .Z(n5864) );
  XNOR U5721 ( .A(n5447), .B(n5859), .Z(n5861) );
  XOR U5722 ( .A(n5865), .B(n5866), .Z(n5447) );
  AND U5723 ( .A(n175), .B(n5867), .Z(n5866) );
  XOR U5724 ( .A(p_input[1304]), .B(p_input[1288]), .Z(n5867) );
  XOR U5725 ( .A(n5868), .B(n5869), .Z(n5859) );
  AND U5726 ( .A(n5870), .B(n5871), .Z(n5869) );
  XOR U5727 ( .A(n5868), .B(n5462), .Z(n5871) );
  XNOR U5728 ( .A(p_input[1319]), .B(n5872), .Z(n5462) );
  AND U5729 ( .A(n178), .B(n5873), .Z(n5872) );
  XOR U5730 ( .A(p_input[1335]), .B(p_input[1319]), .Z(n5873) );
  XNOR U5731 ( .A(n5459), .B(n5868), .Z(n5870) );
  XOR U5732 ( .A(n5874), .B(n5875), .Z(n5459) );
  AND U5733 ( .A(n175), .B(n5876), .Z(n5875) );
  XOR U5734 ( .A(p_input[1303]), .B(p_input[1287]), .Z(n5876) );
  XOR U5735 ( .A(n5877), .B(n5878), .Z(n5868) );
  AND U5736 ( .A(n5879), .B(n5880), .Z(n5878) );
  XOR U5737 ( .A(n5877), .B(n5474), .Z(n5880) );
  XNOR U5738 ( .A(p_input[1318]), .B(n5881), .Z(n5474) );
  AND U5739 ( .A(n178), .B(n5882), .Z(n5881) );
  XOR U5740 ( .A(p_input[1334]), .B(p_input[1318]), .Z(n5882) );
  XNOR U5741 ( .A(n5471), .B(n5877), .Z(n5879) );
  XOR U5742 ( .A(n5883), .B(n5884), .Z(n5471) );
  AND U5743 ( .A(n175), .B(n5885), .Z(n5884) );
  XOR U5744 ( .A(p_input[1302]), .B(p_input[1286]), .Z(n5885) );
  XOR U5745 ( .A(n5886), .B(n5887), .Z(n5877) );
  AND U5746 ( .A(n5888), .B(n5889), .Z(n5887) );
  XOR U5747 ( .A(n5886), .B(n5486), .Z(n5889) );
  XNOR U5748 ( .A(p_input[1317]), .B(n5890), .Z(n5486) );
  AND U5749 ( .A(n178), .B(n5891), .Z(n5890) );
  XOR U5750 ( .A(p_input[1333]), .B(p_input[1317]), .Z(n5891) );
  XNOR U5751 ( .A(n5483), .B(n5886), .Z(n5888) );
  XOR U5752 ( .A(n5892), .B(n5893), .Z(n5483) );
  AND U5753 ( .A(n175), .B(n5894), .Z(n5893) );
  XOR U5754 ( .A(p_input[1301]), .B(p_input[1285]), .Z(n5894) );
  XOR U5755 ( .A(n5895), .B(n5896), .Z(n5886) );
  AND U5756 ( .A(n5897), .B(n5898), .Z(n5896) );
  XOR U5757 ( .A(n5895), .B(n5498), .Z(n5898) );
  XNOR U5758 ( .A(p_input[1316]), .B(n5899), .Z(n5498) );
  AND U5759 ( .A(n178), .B(n5900), .Z(n5899) );
  XOR U5760 ( .A(p_input[1332]), .B(p_input[1316]), .Z(n5900) );
  XNOR U5761 ( .A(n5495), .B(n5895), .Z(n5897) );
  XOR U5762 ( .A(n5901), .B(n5902), .Z(n5495) );
  AND U5763 ( .A(n175), .B(n5903), .Z(n5902) );
  XOR U5764 ( .A(p_input[1300]), .B(p_input[1284]), .Z(n5903) );
  XOR U5765 ( .A(n5904), .B(n5905), .Z(n5895) );
  AND U5766 ( .A(n5906), .B(n5907), .Z(n5905) );
  XOR U5767 ( .A(n5904), .B(n5510), .Z(n5907) );
  XNOR U5768 ( .A(p_input[1315]), .B(n5908), .Z(n5510) );
  AND U5769 ( .A(n178), .B(n5909), .Z(n5908) );
  XOR U5770 ( .A(p_input[1331]), .B(p_input[1315]), .Z(n5909) );
  XNOR U5771 ( .A(n5507), .B(n5904), .Z(n5906) );
  XOR U5772 ( .A(n5910), .B(n5911), .Z(n5507) );
  AND U5773 ( .A(n175), .B(n5912), .Z(n5911) );
  XOR U5774 ( .A(p_input[1299]), .B(p_input[1283]), .Z(n5912) );
  XOR U5775 ( .A(n5913), .B(n5914), .Z(n5904) );
  AND U5776 ( .A(n5915), .B(n5916), .Z(n5914) );
  XOR U5777 ( .A(n5522), .B(n5913), .Z(n5916) );
  XNOR U5778 ( .A(p_input[1314]), .B(n5917), .Z(n5522) );
  AND U5779 ( .A(n178), .B(n5918), .Z(n5917) );
  XOR U5780 ( .A(p_input[1330]), .B(p_input[1314]), .Z(n5918) );
  XNOR U5781 ( .A(n5913), .B(n5519), .Z(n5915) );
  XOR U5782 ( .A(n5919), .B(n5920), .Z(n5519) );
  AND U5783 ( .A(n175), .B(n5921), .Z(n5920) );
  XOR U5784 ( .A(p_input[1298]), .B(p_input[1282]), .Z(n5921) );
  XOR U5785 ( .A(n5922), .B(n5923), .Z(n5913) );
  AND U5786 ( .A(n5924), .B(n5925), .Z(n5923) );
  XNOR U5787 ( .A(n5926), .B(n5535), .Z(n5925) );
  XNOR U5788 ( .A(p_input[1313]), .B(n5927), .Z(n5535) );
  AND U5789 ( .A(n178), .B(n5928), .Z(n5927) );
  XNOR U5790 ( .A(p_input[1329]), .B(n5929), .Z(n5928) );
  IV U5791 ( .A(p_input[1313]), .Z(n5929) );
  XNOR U5792 ( .A(n5532), .B(n5922), .Z(n5924) );
  XNOR U5793 ( .A(p_input[1281]), .B(n5930), .Z(n5532) );
  AND U5794 ( .A(n175), .B(n5931), .Z(n5930) );
  XOR U5795 ( .A(p_input[1297]), .B(p_input[1281]), .Z(n5931) );
  IV U5796 ( .A(n5926), .Z(n5922) );
  AND U5797 ( .A(n5797), .B(n5800), .Z(n5926) );
  XOR U5798 ( .A(p_input[1312]), .B(n5932), .Z(n5800) );
  AND U5799 ( .A(n178), .B(n5933), .Z(n5932) );
  XOR U5800 ( .A(p_input[1328]), .B(p_input[1312]), .Z(n5933) );
  XOR U5801 ( .A(n5934), .B(n5935), .Z(n178) );
  AND U5802 ( .A(n5936), .B(n5937), .Z(n5935) );
  XNOR U5803 ( .A(p_input[1343]), .B(n5934), .Z(n5937) );
  XOR U5804 ( .A(n5934), .B(p_input[1327]), .Z(n5936) );
  XOR U5805 ( .A(n5938), .B(n5939), .Z(n5934) );
  AND U5806 ( .A(n5940), .B(n5941), .Z(n5939) );
  XNOR U5807 ( .A(p_input[1342]), .B(n5938), .Z(n5941) );
  XOR U5808 ( .A(n5938), .B(p_input[1326]), .Z(n5940) );
  XOR U5809 ( .A(n5942), .B(n5943), .Z(n5938) );
  AND U5810 ( .A(n5944), .B(n5945), .Z(n5943) );
  XNOR U5811 ( .A(p_input[1341]), .B(n5942), .Z(n5945) );
  XOR U5812 ( .A(n5942), .B(p_input[1325]), .Z(n5944) );
  XOR U5813 ( .A(n5946), .B(n5947), .Z(n5942) );
  AND U5814 ( .A(n5948), .B(n5949), .Z(n5947) );
  XNOR U5815 ( .A(p_input[1340]), .B(n5946), .Z(n5949) );
  XOR U5816 ( .A(n5946), .B(p_input[1324]), .Z(n5948) );
  XOR U5817 ( .A(n5950), .B(n5951), .Z(n5946) );
  AND U5818 ( .A(n5952), .B(n5953), .Z(n5951) );
  XNOR U5819 ( .A(p_input[1339]), .B(n5950), .Z(n5953) );
  XOR U5820 ( .A(n5950), .B(p_input[1323]), .Z(n5952) );
  XOR U5821 ( .A(n5954), .B(n5955), .Z(n5950) );
  AND U5822 ( .A(n5956), .B(n5957), .Z(n5955) );
  XNOR U5823 ( .A(p_input[1338]), .B(n5954), .Z(n5957) );
  XOR U5824 ( .A(n5954), .B(p_input[1322]), .Z(n5956) );
  XOR U5825 ( .A(n5958), .B(n5959), .Z(n5954) );
  AND U5826 ( .A(n5960), .B(n5961), .Z(n5959) );
  XNOR U5827 ( .A(p_input[1337]), .B(n5958), .Z(n5961) );
  XOR U5828 ( .A(n5958), .B(p_input[1321]), .Z(n5960) );
  XOR U5829 ( .A(n5962), .B(n5963), .Z(n5958) );
  AND U5830 ( .A(n5964), .B(n5965), .Z(n5963) );
  XNOR U5831 ( .A(p_input[1336]), .B(n5962), .Z(n5965) );
  XOR U5832 ( .A(n5962), .B(p_input[1320]), .Z(n5964) );
  XOR U5833 ( .A(n5966), .B(n5967), .Z(n5962) );
  AND U5834 ( .A(n5968), .B(n5969), .Z(n5967) );
  XNOR U5835 ( .A(p_input[1335]), .B(n5966), .Z(n5969) );
  XOR U5836 ( .A(n5966), .B(p_input[1319]), .Z(n5968) );
  XOR U5837 ( .A(n5970), .B(n5971), .Z(n5966) );
  AND U5838 ( .A(n5972), .B(n5973), .Z(n5971) );
  XNOR U5839 ( .A(p_input[1334]), .B(n5970), .Z(n5973) );
  XOR U5840 ( .A(n5970), .B(p_input[1318]), .Z(n5972) );
  XOR U5841 ( .A(n5974), .B(n5975), .Z(n5970) );
  AND U5842 ( .A(n5976), .B(n5977), .Z(n5975) );
  XNOR U5843 ( .A(p_input[1333]), .B(n5974), .Z(n5977) );
  XOR U5844 ( .A(n5974), .B(p_input[1317]), .Z(n5976) );
  XOR U5845 ( .A(n5978), .B(n5979), .Z(n5974) );
  AND U5846 ( .A(n5980), .B(n5981), .Z(n5979) );
  XNOR U5847 ( .A(p_input[1332]), .B(n5978), .Z(n5981) );
  XOR U5848 ( .A(n5978), .B(p_input[1316]), .Z(n5980) );
  XOR U5849 ( .A(n5982), .B(n5983), .Z(n5978) );
  AND U5850 ( .A(n5984), .B(n5985), .Z(n5983) );
  XNOR U5851 ( .A(p_input[1331]), .B(n5982), .Z(n5985) );
  XOR U5852 ( .A(n5982), .B(p_input[1315]), .Z(n5984) );
  XOR U5853 ( .A(n5986), .B(n5987), .Z(n5982) );
  AND U5854 ( .A(n5988), .B(n5989), .Z(n5987) );
  XNOR U5855 ( .A(p_input[1330]), .B(n5986), .Z(n5989) );
  XOR U5856 ( .A(n5986), .B(p_input[1314]), .Z(n5988) );
  XNOR U5857 ( .A(n5990), .B(n5991), .Z(n5986) );
  AND U5858 ( .A(n5992), .B(n5993), .Z(n5991) );
  XOR U5859 ( .A(p_input[1329]), .B(n5990), .Z(n5993) );
  XNOR U5860 ( .A(p_input[1313]), .B(n5990), .Z(n5992) );
  AND U5861 ( .A(p_input[1328]), .B(n5994), .Z(n5990) );
  IV U5862 ( .A(p_input[1312]), .Z(n5994) );
  XNOR U5863 ( .A(p_input[1280]), .B(n5995), .Z(n5797) );
  AND U5864 ( .A(n175), .B(n5996), .Z(n5995) );
  XOR U5865 ( .A(p_input[1296]), .B(p_input[1280]), .Z(n5996) );
  XOR U5866 ( .A(n5997), .B(n5998), .Z(n175) );
  AND U5867 ( .A(n5999), .B(n6000), .Z(n5998) );
  XNOR U5868 ( .A(p_input[1311]), .B(n5997), .Z(n6000) );
  XOR U5869 ( .A(n5997), .B(p_input[1295]), .Z(n5999) );
  XOR U5870 ( .A(n6001), .B(n6002), .Z(n5997) );
  AND U5871 ( .A(n6003), .B(n6004), .Z(n6002) );
  XNOR U5872 ( .A(p_input[1310]), .B(n6001), .Z(n6004) );
  XNOR U5873 ( .A(n6001), .B(n5811), .Z(n6003) );
  IV U5874 ( .A(p_input[1294]), .Z(n5811) );
  XOR U5875 ( .A(n6005), .B(n6006), .Z(n6001) );
  AND U5876 ( .A(n6007), .B(n6008), .Z(n6006) );
  XNOR U5877 ( .A(p_input[1309]), .B(n6005), .Z(n6008) );
  XNOR U5878 ( .A(n6005), .B(n5820), .Z(n6007) );
  IV U5879 ( .A(p_input[1293]), .Z(n5820) );
  XOR U5880 ( .A(n6009), .B(n6010), .Z(n6005) );
  AND U5881 ( .A(n6011), .B(n6012), .Z(n6010) );
  XNOR U5882 ( .A(p_input[1308]), .B(n6009), .Z(n6012) );
  XNOR U5883 ( .A(n6009), .B(n5829), .Z(n6011) );
  IV U5884 ( .A(p_input[1292]), .Z(n5829) );
  XOR U5885 ( .A(n6013), .B(n6014), .Z(n6009) );
  AND U5886 ( .A(n6015), .B(n6016), .Z(n6014) );
  XNOR U5887 ( .A(p_input[1307]), .B(n6013), .Z(n6016) );
  XNOR U5888 ( .A(n6013), .B(n5838), .Z(n6015) );
  IV U5889 ( .A(p_input[1291]), .Z(n5838) );
  XOR U5890 ( .A(n6017), .B(n6018), .Z(n6013) );
  AND U5891 ( .A(n6019), .B(n6020), .Z(n6018) );
  XNOR U5892 ( .A(p_input[1306]), .B(n6017), .Z(n6020) );
  XNOR U5893 ( .A(n6017), .B(n5847), .Z(n6019) );
  IV U5894 ( .A(p_input[1290]), .Z(n5847) );
  XOR U5895 ( .A(n6021), .B(n6022), .Z(n6017) );
  AND U5896 ( .A(n6023), .B(n6024), .Z(n6022) );
  XNOR U5897 ( .A(p_input[1305]), .B(n6021), .Z(n6024) );
  XNOR U5898 ( .A(n6021), .B(n5856), .Z(n6023) );
  IV U5899 ( .A(p_input[1289]), .Z(n5856) );
  XOR U5900 ( .A(n6025), .B(n6026), .Z(n6021) );
  AND U5901 ( .A(n6027), .B(n6028), .Z(n6026) );
  XNOR U5902 ( .A(p_input[1304]), .B(n6025), .Z(n6028) );
  XNOR U5903 ( .A(n6025), .B(n5865), .Z(n6027) );
  IV U5904 ( .A(p_input[1288]), .Z(n5865) );
  XOR U5905 ( .A(n6029), .B(n6030), .Z(n6025) );
  AND U5906 ( .A(n6031), .B(n6032), .Z(n6030) );
  XNOR U5907 ( .A(p_input[1303]), .B(n6029), .Z(n6032) );
  XNOR U5908 ( .A(n6029), .B(n5874), .Z(n6031) );
  IV U5909 ( .A(p_input[1287]), .Z(n5874) );
  XOR U5910 ( .A(n6033), .B(n6034), .Z(n6029) );
  AND U5911 ( .A(n6035), .B(n6036), .Z(n6034) );
  XNOR U5912 ( .A(p_input[1302]), .B(n6033), .Z(n6036) );
  XNOR U5913 ( .A(n6033), .B(n5883), .Z(n6035) );
  IV U5914 ( .A(p_input[1286]), .Z(n5883) );
  XOR U5915 ( .A(n6037), .B(n6038), .Z(n6033) );
  AND U5916 ( .A(n6039), .B(n6040), .Z(n6038) );
  XNOR U5917 ( .A(p_input[1301]), .B(n6037), .Z(n6040) );
  XNOR U5918 ( .A(n6037), .B(n5892), .Z(n6039) );
  IV U5919 ( .A(p_input[1285]), .Z(n5892) );
  XOR U5920 ( .A(n6041), .B(n6042), .Z(n6037) );
  AND U5921 ( .A(n6043), .B(n6044), .Z(n6042) );
  XNOR U5922 ( .A(p_input[1300]), .B(n6041), .Z(n6044) );
  XNOR U5923 ( .A(n6041), .B(n5901), .Z(n6043) );
  IV U5924 ( .A(p_input[1284]), .Z(n5901) );
  XOR U5925 ( .A(n6045), .B(n6046), .Z(n6041) );
  AND U5926 ( .A(n6047), .B(n6048), .Z(n6046) );
  XNOR U5927 ( .A(p_input[1299]), .B(n6045), .Z(n6048) );
  XNOR U5928 ( .A(n6045), .B(n5910), .Z(n6047) );
  IV U5929 ( .A(p_input[1283]), .Z(n5910) );
  XOR U5930 ( .A(n6049), .B(n6050), .Z(n6045) );
  AND U5931 ( .A(n6051), .B(n6052), .Z(n6050) );
  XNOR U5932 ( .A(p_input[1298]), .B(n6049), .Z(n6052) );
  XNOR U5933 ( .A(n6049), .B(n5919), .Z(n6051) );
  IV U5934 ( .A(p_input[1282]), .Z(n5919) );
  XNOR U5935 ( .A(n6053), .B(n6054), .Z(n6049) );
  AND U5936 ( .A(n6055), .B(n6056), .Z(n6054) );
  XOR U5937 ( .A(p_input[1297]), .B(n6053), .Z(n6056) );
  XNOR U5938 ( .A(p_input[1281]), .B(n6053), .Z(n6055) );
  AND U5939 ( .A(p_input[1296]), .B(n6057), .Z(n6053) );
  IV U5940 ( .A(p_input[1280]), .Z(n6057) );
  XOR U5941 ( .A(n6058), .B(n6059), .Z(n4285) );
  AND U5942 ( .A(n499), .B(n6060), .Z(n6059) );
  XNOR U5943 ( .A(n6061), .B(n6058), .Z(n6060) );
  XOR U5944 ( .A(n6062), .B(n6063), .Z(n499) );
  AND U5945 ( .A(n6064), .B(n6065), .Z(n6063) );
  XNOR U5946 ( .A(n4300), .B(n6062), .Z(n6065) );
  AND U5947 ( .A(n6066), .B(n6067), .Z(n4300) );
  XNOR U5948 ( .A(n6062), .B(n4297), .Z(n6064) );
  IV U5949 ( .A(n6068), .Z(n4297) );
  AND U5950 ( .A(n6069), .B(n6070), .Z(n6068) );
  XOR U5951 ( .A(n6071), .B(n6072), .Z(n6062) );
  AND U5952 ( .A(n6073), .B(n6074), .Z(n6072) );
  XOR U5953 ( .A(n6071), .B(n4312), .Z(n6074) );
  XOR U5954 ( .A(n6075), .B(n6076), .Z(n4312) );
  AND U5955 ( .A(n426), .B(n6077), .Z(n6076) );
  XOR U5956 ( .A(n6078), .B(n6075), .Z(n6077) );
  XNOR U5957 ( .A(n4309), .B(n6071), .Z(n6073) );
  XOR U5958 ( .A(n6079), .B(n6080), .Z(n4309) );
  AND U5959 ( .A(n423), .B(n6081), .Z(n6080) );
  XOR U5960 ( .A(n6082), .B(n6079), .Z(n6081) );
  XOR U5961 ( .A(n6083), .B(n6084), .Z(n6071) );
  AND U5962 ( .A(n6085), .B(n6086), .Z(n6084) );
  XOR U5963 ( .A(n6083), .B(n4324), .Z(n6086) );
  XOR U5964 ( .A(n6087), .B(n6088), .Z(n4324) );
  AND U5965 ( .A(n426), .B(n6089), .Z(n6088) );
  XOR U5966 ( .A(n6090), .B(n6087), .Z(n6089) );
  XNOR U5967 ( .A(n4321), .B(n6083), .Z(n6085) );
  XOR U5968 ( .A(n6091), .B(n6092), .Z(n4321) );
  AND U5969 ( .A(n423), .B(n6093), .Z(n6092) );
  XOR U5970 ( .A(n6094), .B(n6091), .Z(n6093) );
  XOR U5971 ( .A(n6095), .B(n6096), .Z(n6083) );
  AND U5972 ( .A(n6097), .B(n6098), .Z(n6096) );
  XOR U5973 ( .A(n6095), .B(n4336), .Z(n6098) );
  XOR U5974 ( .A(n6099), .B(n6100), .Z(n4336) );
  AND U5975 ( .A(n426), .B(n6101), .Z(n6100) );
  XOR U5976 ( .A(n6102), .B(n6099), .Z(n6101) );
  XNOR U5977 ( .A(n4333), .B(n6095), .Z(n6097) );
  XOR U5978 ( .A(n6103), .B(n6104), .Z(n4333) );
  AND U5979 ( .A(n423), .B(n6105), .Z(n6104) );
  XOR U5980 ( .A(n6106), .B(n6103), .Z(n6105) );
  XOR U5981 ( .A(n6107), .B(n6108), .Z(n6095) );
  AND U5982 ( .A(n6109), .B(n6110), .Z(n6108) );
  XOR U5983 ( .A(n6107), .B(n4348), .Z(n6110) );
  XOR U5984 ( .A(n6111), .B(n6112), .Z(n4348) );
  AND U5985 ( .A(n426), .B(n6113), .Z(n6112) );
  XOR U5986 ( .A(n6114), .B(n6111), .Z(n6113) );
  XNOR U5987 ( .A(n4345), .B(n6107), .Z(n6109) );
  XOR U5988 ( .A(n6115), .B(n6116), .Z(n4345) );
  AND U5989 ( .A(n423), .B(n6117), .Z(n6116) );
  XOR U5990 ( .A(n6118), .B(n6115), .Z(n6117) );
  XOR U5991 ( .A(n6119), .B(n6120), .Z(n6107) );
  AND U5992 ( .A(n6121), .B(n6122), .Z(n6120) );
  XOR U5993 ( .A(n6119), .B(n4360), .Z(n6122) );
  XOR U5994 ( .A(n6123), .B(n6124), .Z(n4360) );
  AND U5995 ( .A(n426), .B(n6125), .Z(n6124) );
  XOR U5996 ( .A(n6126), .B(n6123), .Z(n6125) );
  XNOR U5997 ( .A(n4357), .B(n6119), .Z(n6121) );
  XOR U5998 ( .A(n6127), .B(n6128), .Z(n4357) );
  AND U5999 ( .A(n423), .B(n6129), .Z(n6128) );
  XOR U6000 ( .A(n6130), .B(n6127), .Z(n6129) );
  XOR U6001 ( .A(n6131), .B(n6132), .Z(n6119) );
  AND U6002 ( .A(n6133), .B(n6134), .Z(n6132) );
  XOR U6003 ( .A(n6131), .B(n4372), .Z(n6134) );
  XOR U6004 ( .A(n6135), .B(n6136), .Z(n4372) );
  AND U6005 ( .A(n426), .B(n6137), .Z(n6136) );
  XOR U6006 ( .A(n6138), .B(n6135), .Z(n6137) );
  XNOR U6007 ( .A(n4369), .B(n6131), .Z(n6133) );
  XOR U6008 ( .A(n6139), .B(n6140), .Z(n4369) );
  AND U6009 ( .A(n423), .B(n6141), .Z(n6140) );
  XOR U6010 ( .A(n6142), .B(n6139), .Z(n6141) );
  XOR U6011 ( .A(n6143), .B(n6144), .Z(n6131) );
  AND U6012 ( .A(n6145), .B(n6146), .Z(n6144) );
  XOR U6013 ( .A(n6143), .B(n4384), .Z(n6146) );
  XOR U6014 ( .A(n6147), .B(n6148), .Z(n4384) );
  AND U6015 ( .A(n426), .B(n6149), .Z(n6148) );
  XOR U6016 ( .A(n6150), .B(n6147), .Z(n6149) );
  XNOR U6017 ( .A(n4381), .B(n6143), .Z(n6145) );
  XOR U6018 ( .A(n6151), .B(n6152), .Z(n4381) );
  AND U6019 ( .A(n423), .B(n6153), .Z(n6152) );
  XOR U6020 ( .A(n6154), .B(n6151), .Z(n6153) );
  XOR U6021 ( .A(n6155), .B(n6156), .Z(n6143) );
  AND U6022 ( .A(n6157), .B(n6158), .Z(n6156) );
  XOR U6023 ( .A(n6155), .B(n4396), .Z(n6158) );
  XOR U6024 ( .A(n6159), .B(n6160), .Z(n4396) );
  AND U6025 ( .A(n426), .B(n6161), .Z(n6160) );
  XOR U6026 ( .A(n6162), .B(n6159), .Z(n6161) );
  XNOR U6027 ( .A(n4393), .B(n6155), .Z(n6157) );
  XOR U6028 ( .A(n6163), .B(n6164), .Z(n4393) );
  AND U6029 ( .A(n423), .B(n6165), .Z(n6164) );
  XOR U6030 ( .A(n6166), .B(n6163), .Z(n6165) );
  XOR U6031 ( .A(n6167), .B(n6168), .Z(n6155) );
  AND U6032 ( .A(n6169), .B(n6170), .Z(n6168) );
  XOR U6033 ( .A(n6167), .B(n4408), .Z(n6170) );
  XOR U6034 ( .A(n6171), .B(n6172), .Z(n4408) );
  AND U6035 ( .A(n426), .B(n6173), .Z(n6172) );
  XOR U6036 ( .A(n6174), .B(n6171), .Z(n6173) );
  XNOR U6037 ( .A(n4405), .B(n6167), .Z(n6169) );
  XOR U6038 ( .A(n6175), .B(n6176), .Z(n4405) );
  AND U6039 ( .A(n423), .B(n6177), .Z(n6176) );
  XOR U6040 ( .A(n6178), .B(n6175), .Z(n6177) );
  XOR U6041 ( .A(n6179), .B(n6180), .Z(n6167) );
  AND U6042 ( .A(n6181), .B(n6182), .Z(n6180) );
  XOR U6043 ( .A(n6179), .B(n4420), .Z(n6182) );
  XOR U6044 ( .A(n6183), .B(n6184), .Z(n4420) );
  AND U6045 ( .A(n426), .B(n6185), .Z(n6184) );
  XOR U6046 ( .A(n6186), .B(n6183), .Z(n6185) );
  XNOR U6047 ( .A(n4417), .B(n6179), .Z(n6181) );
  XOR U6048 ( .A(n6187), .B(n6188), .Z(n4417) );
  AND U6049 ( .A(n423), .B(n6189), .Z(n6188) );
  XOR U6050 ( .A(n6190), .B(n6187), .Z(n6189) );
  XOR U6051 ( .A(n6191), .B(n6192), .Z(n6179) );
  AND U6052 ( .A(n6193), .B(n6194), .Z(n6192) );
  XOR U6053 ( .A(n6191), .B(n4432), .Z(n6194) );
  XOR U6054 ( .A(n6195), .B(n6196), .Z(n4432) );
  AND U6055 ( .A(n426), .B(n6197), .Z(n6196) );
  XOR U6056 ( .A(n6198), .B(n6195), .Z(n6197) );
  XNOR U6057 ( .A(n4429), .B(n6191), .Z(n6193) );
  XOR U6058 ( .A(n6199), .B(n6200), .Z(n4429) );
  AND U6059 ( .A(n423), .B(n6201), .Z(n6200) );
  XOR U6060 ( .A(n6202), .B(n6199), .Z(n6201) );
  XOR U6061 ( .A(n6203), .B(n6204), .Z(n6191) );
  AND U6062 ( .A(n6205), .B(n6206), .Z(n6204) );
  XOR U6063 ( .A(n6203), .B(n4444), .Z(n6206) );
  XOR U6064 ( .A(n6207), .B(n6208), .Z(n4444) );
  AND U6065 ( .A(n426), .B(n6209), .Z(n6208) );
  XOR U6066 ( .A(n6210), .B(n6207), .Z(n6209) );
  XNOR U6067 ( .A(n4441), .B(n6203), .Z(n6205) );
  XOR U6068 ( .A(n6211), .B(n6212), .Z(n4441) );
  AND U6069 ( .A(n423), .B(n6213), .Z(n6212) );
  XOR U6070 ( .A(n6214), .B(n6211), .Z(n6213) );
  XOR U6071 ( .A(n6215), .B(n6216), .Z(n6203) );
  AND U6072 ( .A(n6217), .B(n6218), .Z(n6216) );
  XOR U6073 ( .A(n4456), .B(n6215), .Z(n6218) );
  XOR U6074 ( .A(n6219), .B(n6220), .Z(n4456) );
  AND U6075 ( .A(n426), .B(n6221), .Z(n6220) );
  XOR U6076 ( .A(n6219), .B(n6222), .Z(n6221) );
  XNOR U6077 ( .A(n6215), .B(n4453), .Z(n6217) );
  XOR U6078 ( .A(n6223), .B(n6224), .Z(n4453) );
  AND U6079 ( .A(n423), .B(n6225), .Z(n6224) );
  XOR U6080 ( .A(n6223), .B(n6226), .Z(n6225) );
  XOR U6081 ( .A(n6227), .B(n6228), .Z(n6215) );
  AND U6082 ( .A(n6229), .B(n6230), .Z(n6228) );
  XNOR U6083 ( .A(n6231), .B(n4469), .Z(n6230) );
  XOR U6084 ( .A(n6232), .B(n6233), .Z(n4469) );
  AND U6085 ( .A(n426), .B(n6234), .Z(n6233) );
  XOR U6086 ( .A(n6235), .B(n6232), .Z(n6234) );
  XNOR U6087 ( .A(n4466), .B(n6227), .Z(n6229) );
  XOR U6088 ( .A(n6236), .B(n6237), .Z(n4466) );
  AND U6089 ( .A(n423), .B(n6238), .Z(n6237) );
  XOR U6090 ( .A(n6239), .B(n6236), .Z(n6238) );
  IV U6091 ( .A(n6231), .Z(n6227) );
  AND U6092 ( .A(n6058), .B(n6061), .Z(n6231) );
  XNOR U6093 ( .A(n6240), .B(n6241), .Z(n6061) );
  AND U6094 ( .A(n426), .B(n6242), .Z(n6241) );
  XNOR U6095 ( .A(n6243), .B(n6240), .Z(n6242) );
  XOR U6096 ( .A(n6244), .B(n6245), .Z(n426) );
  AND U6097 ( .A(n6246), .B(n6247), .Z(n6245) );
  XNOR U6098 ( .A(n6066), .B(n6244), .Z(n6247) );
  AND U6099 ( .A(n6248), .B(n6249), .Z(n6066) );
  XOR U6100 ( .A(n6244), .B(n6067), .Z(n6246) );
  AND U6101 ( .A(n6250), .B(n6251), .Z(n6067) );
  XOR U6102 ( .A(n6252), .B(n6253), .Z(n6244) );
  AND U6103 ( .A(n6254), .B(n6255), .Z(n6253) );
  XOR U6104 ( .A(n6252), .B(n6078), .Z(n6255) );
  XOR U6105 ( .A(n6256), .B(n6257), .Z(n6078) );
  AND U6106 ( .A(n266), .B(n6258), .Z(n6257) );
  XOR U6107 ( .A(n6259), .B(n6256), .Z(n6258) );
  XNOR U6108 ( .A(n6075), .B(n6252), .Z(n6254) );
  XOR U6109 ( .A(n6260), .B(n6261), .Z(n6075) );
  AND U6110 ( .A(n264), .B(n6262), .Z(n6261) );
  XOR U6111 ( .A(n6263), .B(n6260), .Z(n6262) );
  XOR U6112 ( .A(n6264), .B(n6265), .Z(n6252) );
  AND U6113 ( .A(n6266), .B(n6267), .Z(n6265) );
  XOR U6114 ( .A(n6264), .B(n6090), .Z(n6267) );
  XOR U6115 ( .A(n6268), .B(n6269), .Z(n6090) );
  AND U6116 ( .A(n266), .B(n6270), .Z(n6269) );
  XOR U6117 ( .A(n6271), .B(n6268), .Z(n6270) );
  XNOR U6118 ( .A(n6087), .B(n6264), .Z(n6266) );
  XOR U6119 ( .A(n6272), .B(n6273), .Z(n6087) );
  AND U6120 ( .A(n264), .B(n6274), .Z(n6273) );
  XOR U6121 ( .A(n6275), .B(n6272), .Z(n6274) );
  XOR U6122 ( .A(n6276), .B(n6277), .Z(n6264) );
  AND U6123 ( .A(n6278), .B(n6279), .Z(n6277) );
  XOR U6124 ( .A(n6276), .B(n6102), .Z(n6279) );
  XOR U6125 ( .A(n6280), .B(n6281), .Z(n6102) );
  AND U6126 ( .A(n266), .B(n6282), .Z(n6281) );
  XOR U6127 ( .A(n6283), .B(n6280), .Z(n6282) );
  XNOR U6128 ( .A(n6099), .B(n6276), .Z(n6278) );
  XOR U6129 ( .A(n6284), .B(n6285), .Z(n6099) );
  AND U6130 ( .A(n264), .B(n6286), .Z(n6285) );
  XOR U6131 ( .A(n6287), .B(n6284), .Z(n6286) );
  XOR U6132 ( .A(n6288), .B(n6289), .Z(n6276) );
  AND U6133 ( .A(n6290), .B(n6291), .Z(n6289) );
  XOR U6134 ( .A(n6288), .B(n6114), .Z(n6291) );
  XOR U6135 ( .A(n6292), .B(n6293), .Z(n6114) );
  AND U6136 ( .A(n266), .B(n6294), .Z(n6293) );
  XOR U6137 ( .A(n6295), .B(n6292), .Z(n6294) );
  XNOR U6138 ( .A(n6111), .B(n6288), .Z(n6290) );
  XOR U6139 ( .A(n6296), .B(n6297), .Z(n6111) );
  AND U6140 ( .A(n264), .B(n6298), .Z(n6297) );
  XOR U6141 ( .A(n6299), .B(n6296), .Z(n6298) );
  XOR U6142 ( .A(n6300), .B(n6301), .Z(n6288) );
  AND U6143 ( .A(n6302), .B(n6303), .Z(n6301) );
  XOR U6144 ( .A(n6300), .B(n6126), .Z(n6303) );
  XOR U6145 ( .A(n6304), .B(n6305), .Z(n6126) );
  AND U6146 ( .A(n266), .B(n6306), .Z(n6305) );
  XOR U6147 ( .A(n6307), .B(n6304), .Z(n6306) );
  XNOR U6148 ( .A(n6123), .B(n6300), .Z(n6302) );
  XOR U6149 ( .A(n6308), .B(n6309), .Z(n6123) );
  AND U6150 ( .A(n264), .B(n6310), .Z(n6309) );
  XOR U6151 ( .A(n6311), .B(n6308), .Z(n6310) );
  XOR U6152 ( .A(n6312), .B(n6313), .Z(n6300) );
  AND U6153 ( .A(n6314), .B(n6315), .Z(n6313) );
  XOR U6154 ( .A(n6312), .B(n6138), .Z(n6315) );
  XOR U6155 ( .A(n6316), .B(n6317), .Z(n6138) );
  AND U6156 ( .A(n266), .B(n6318), .Z(n6317) );
  XOR U6157 ( .A(n6319), .B(n6316), .Z(n6318) );
  XNOR U6158 ( .A(n6135), .B(n6312), .Z(n6314) );
  XOR U6159 ( .A(n6320), .B(n6321), .Z(n6135) );
  AND U6160 ( .A(n264), .B(n6322), .Z(n6321) );
  XOR U6161 ( .A(n6323), .B(n6320), .Z(n6322) );
  XOR U6162 ( .A(n6324), .B(n6325), .Z(n6312) );
  AND U6163 ( .A(n6326), .B(n6327), .Z(n6325) );
  XOR U6164 ( .A(n6324), .B(n6150), .Z(n6327) );
  XOR U6165 ( .A(n6328), .B(n6329), .Z(n6150) );
  AND U6166 ( .A(n266), .B(n6330), .Z(n6329) );
  XOR U6167 ( .A(n6331), .B(n6328), .Z(n6330) );
  XNOR U6168 ( .A(n6147), .B(n6324), .Z(n6326) );
  XOR U6169 ( .A(n6332), .B(n6333), .Z(n6147) );
  AND U6170 ( .A(n264), .B(n6334), .Z(n6333) );
  XOR U6171 ( .A(n6335), .B(n6332), .Z(n6334) );
  XOR U6172 ( .A(n6336), .B(n6337), .Z(n6324) );
  AND U6173 ( .A(n6338), .B(n6339), .Z(n6337) );
  XOR U6174 ( .A(n6336), .B(n6162), .Z(n6339) );
  XOR U6175 ( .A(n6340), .B(n6341), .Z(n6162) );
  AND U6176 ( .A(n266), .B(n6342), .Z(n6341) );
  XOR U6177 ( .A(n6343), .B(n6340), .Z(n6342) );
  XNOR U6178 ( .A(n6159), .B(n6336), .Z(n6338) );
  XOR U6179 ( .A(n6344), .B(n6345), .Z(n6159) );
  AND U6180 ( .A(n264), .B(n6346), .Z(n6345) );
  XOR U6181 ( .A(n6347), .B(n6344), .Z(n6346) );
  XOR U6182 ( .A(n6348), .B(n6349), .Z(n6336) );
  AND U6183 ( .A(n6350), .B(n6351), .Z(n6349) );
  XOR U6184 ( .A(n6348), .B(n6174), .Z(n6351) );
  XOR U6185 ( .A(n6352), .B(n6353), .Z(n6174) );
  AND U6186 ( .A(n266), .B(n6354), .Z(n6353) );
  XOR U6187 ( .A(n6355), .B(n6352), .Z(n6354) );
  XNOR U6188 ( .A(n6171), .B(n6348), .Z(n6350) );
  XOR U6189 ( .A(n6356), .B(n6357), .Z(n6171) );
  AND U6190 ( .A(n264), .B(n6358), .Z(n6357) );
  XOR U6191 ( .A(n6359), .B(n6356), .Z(n6358) );
  XOR U6192 ( .A(n6360), .B(n6361), .Z(n6348) );
  AND U6193 ( .A(n6362), .B(n6363), .Z(n6361) );
  XOR U6194 ( .A(n6360), .B(n6186), .Z(n6363) );
  XOR U6195 ( .A(n6364), .B(n6365), .Z(n6186) );
  AND U6196 ( .A(n266), .B(n6366), .Z(n6365) );
  XOR U6197 ( .A(n6367), .B(n6364), .Z(n6366) );
  XNOR U6198 ( .A(n6183), .B(n6360), .Z(n6362) );
  XOR U6199 ( .A(n6368), .B(n6369), .Z(n6183) );
  AND U6200 ( .A(n264), .B(n6370), .Z(n6369) );
  XOR U6201 ( .A(n6371), .B(n6368), .Z(n6370) );
  XOR U6202 ( .A(n6372), .B(n6373), .Z(n6360) );
  AND U6203 ( .A(n6374), .B(n6375), .Z(n6373) );
  XOR U6204 ( .A(n6372), .B(n6198), .Z(n6375) );
  XOR U6205 ( .A(n6376), .B(n6377), .Z(n6198) );
  AND U6206 ( .A(n266), .B(n6378), .Z(n6377) );
  XOR U6207 ( .A(n6379), .B(n6376), .Z(n6378) );
  XNOR U6208 ( .A(n6195), .B(n6372), .Z(n6374) );
  XOR U6209 ( .A(n6380), .B(n6381), .Z(n6195) );
  AND U6210 ( .A(n264), .B(n6382), .Z(n6381) );
  XOR U6211 ( .A(n6383), .B(n6380), .Z(n6382) );
  XOR U6212 ( .A(n6384), .B(n6385), .Z(n6372) );
  AND U6213 ( .A(n6386), .B(n6387), .Z(n6385) );
  XOR U6214 ( .A(n6384), .B(n6210), .Z(n6387) );
  XOR U6215 ( .A(n6388), .B(n6389), .Z(n6210) );
  AND U6216 ( .A(n266), .B(n6390), .Z(n6389) );
  XOR U6217 ( .A(n6391), .B(n6388), .Z(n6390) );
  XNOR U6218 ( .A(n6207), .B(n6384), .Z(n6386) );
  XOR U6219 ( .A(n6392), .B(n6393), .Z(n6207) );
  AND U6220 ( .A(n264), .B(n6394), .Z(n6393) );
  XOR U6221 ( .A(n6395), .B(n6392), .Z(n6394) );
  XOR U6222 ( .A(n6396), .B(n6397), .Z(n6384) );
  AND U6223 ( .A(n6398), .B(n6399), .Z(n6397) );
  XOR U6224 ( .A(n6222), .B(n6396), .Z(n6399) );
  XOR U6225 ( .A(n6400), .B(n6401), .Z(n6222) );
  AND U6226 ( .A(n266), .B(n6402), .Z(n6401) );
  XOR U6227 ( .A(n6400), .B(n6403), .Z(n6402) );
  XNOR U6228 ( .A(n6396), .B(n6219), .Z(n6398) );
  XOR U6229 ( .A(n6404), .B(n6405), .Z(n6219) );
  AND U6230 ( .A(n264), .B(n6406), .Z(n6405) );
  XOR U6231 ( .A(n6404), .B(n6407), .Z(n6406) );
  XOR U6232 ( .A(n6408), .B(n6409), .Z(n6396) );
  AND U6233 ( .A(n6410), .B(n6411), .Z(n6409) );
  XNOR U6234 ( .A(n6412), .B(n6235), .Z(n6411) );
  XOR U6235 ( .A(n6413), .B(n6414), .Z(n6235) );
  AND U6236 ( .A(n266), .B(n6415), .Z(n6414) );
  XOR U6237 ( .A(n6416), .B(n6413), .Z(n6415) );
  XNOR U6238 ( .A(n6232), .B(n6408), .Z(n6410) );
  XOR U6239 ( .A(n6417), .B(n6418), .Z(n6232) );
  AND U6240 ( .A(n264), .B(n6419), .Z(n6418) );
  XOR U6241 ( .A(n6420), .B(n6417), .Z(n6419) );
  IV U6242 ( .A(n6412), .Z(n6408) );
  AND U6243 ( .A(n6240), .B(n6243), .Z(n6412) );
  XNOR U6244 ( .A(n6421), .B(n6422), .Z(n6243) );
  AND U6245 ( .A(n266), .B(n6423), .Z(n6422) );
  XNOR U6246 ( .A(n6424), .B(n6421), .Z(n6423) );
  XOR U6247 ( .A(n6425), .B(n6426), .Z(n266) );
  AND U6248 ( .A(n6427), .B(n6428), .Z(n6426) );
  XNOR U6249 ( .A(n6248), .B(n6425), .Z(n6428) );
  AND U6250 ( .A(p_input[1279]), .B(p_input[1263]), .Z(n6248) );
  XOR U6251 ( .A(n6425), .B(n6249), .Z(n6427) );
  AND U6252 ( .A(p_input[1247]), .B(p_input[1231]), .Z(n6249) );
  XOR U6253 ( .A(n6429), .B(n6430), .Z(n6425) );
  AND U6254 ( .A(n6431), .B(n6432), .Z(n6430) );
  XOR U6255 ( .A(n6429), .B(n6259), .Z(n6432) );
  XNOR U6256 ( .A(p_input[1262]), .B(n6433), .Z(n6259) );
  AND U6257 ( .A(n190), .B(n6434), .Z(n6433) );
  XOR U6258 ( .A(p_input[1278]), .B(p_input[1262]), .Z(n6434) );
  XNOR U6259 ( .A(n6256), .B(n6429), .Z(n6431) );
  XOR U6260 ( .A(n6435), .B(n6436), .Z(n6256) );
  AND U6261 ( .A(n188), .B(n6437), .Z(n6436) );
  XOR U6262 ( .A(p_input[1246]), .B(p_input[1230]), .Z(n6437) );
  XOR U6263 ( .A(n6438), .B(n6439), .Z(n6429) );
  AND U6264 ( .A(n6440), .B(n6441), .Z(n6439) );
  XOR U6265 ( .A(n6438), .B(n6271), .Z(n6441) );
  XNOR U6266 ( .A(p_input[1261]), .B(n6442), .Z(n6271) );
  AND U6267 ( .A(n190), .B(n6443), .Z(n6442) );
  XOR U6268 ( .A(p_input[1277]), .B(p_input[1261]), .Z(n6443) );
  XNOR U6269 ( .A(n6268), .B(n6438), .Z(n6440) );
  XOR U6270 ( .A(n6444), .B(n6445), .Z(n6268) );
  AND U6271 ( .A(n188), .B(n6446), .Z(n6445) );
  XOR U6272 ( .A(p_input[1245]), .B(p_input[1229]), .Z(n6446) );
  XOR U6273 ( .A(n6447), .B(n6448), .Z(n6438) );
  AND U6274 ( .A(n6449), .B(n6450), .Z(n6448) );
  XOR U6275 ( .A(n6447), .B(n6283), .Z(n6450) );
  XNOR U6276 ( .A(p_input[1260]), .B(n6451), .Z(n6283) );
  AND U6277 ( .A(n190), .B(n6452), .Z(n6451) );
  XOR U6278 ( .A(p_input[1276]), .B(p_input[1260]), .Z(n6452) );
  XNOR U6279 ( .A(n6280), .B(n6447), .Z(n6449) );
  XOR U6280 ( .A(n6453), .B(n6454), .Z(n6280) );
  AND U6281 ( .A(n188), .B(n6455), .Z(n6454) );
  XOR U6282 ( .A(p_input[1244]), .B(p_input[1228]), .Z(n6455) );
  XOR U6283 ( .A(n6456), .B(n6457), .Z(n6447) );
  AND U6284 ( .A(n6458), .B(n6459), .Z(n6457) );
  XOR U6285 ( .A(n6456), .B(n6295), .Z(n6459) );
  XNOR U6286 ( .A(p_input[1259]), .B(n6460), .Z(n6295) );
  AND U6287 ( .A(n190), .B(n6461), .Z(n6460) );
  XOR U6288 ( .A(p_input[1275]), .B(p_input[1259]), .Z(n6461) );
  XNOR U6289 ( .A(n6292), .B(n6456), .Z(n6458) );
  XOR U6290 ( .A(n6462), .B(n6463), .Z(n6292) );
  AND U6291 ( .A(n188), .B(n6464), .Z(n6463) );
  XOR U6292 ( .A(p_input[1243]), .B(p_input[1227]), .Z(n6464) );
  XOR U6293 ( .A(n6465), .B(n6466), .Z(n6456) );
  AND U6294 ( .A(n6467), .B(n6468), .Z(n6466) );
  XOR U6295 ( .A(n6465), .B(n6307), .Z(n6468) );
  XNOR U6296 ( .A(p_input[1258]), .B(n6469), .Z(n6307) );
  AND U6297 ( .A(n190), .B(n6470), .Z(n6469) );
  XOR U6298 ( .A(p_input[1274]), .B(p_input[1258]), .Z(n6470) );
  XNOR U6299 ( .A(n6304), .B(n6465), .Z(n6467) );
  XOR U6300 ( .A(n6471), .B(n6472), .Z(n6304) );
  AND U6301 ( .A(n188), .B(n6473), .Z(n6472) );
  XOR U6302 ( .A(p_input[1242]), .B(p_input[1226]), .Z(n6473) );
  XOR U6303 ( .A(n6474), .B(n6475), .Z(n6465) );
  AND U6304 ( .A(n6476), .B(n6477), .Z(n6475) );
  XOR U6305 ( .A(n6474), .B(n6319), .Z(n6477) );
  XNOR U6306 ( .A(p_input[1257]), .B(n6478), .Z(n6319) );
  AND U6307 ( .A(n190), .B(n6479), .Z(n6478) );
  XOR U6308 ( .A(p_input[1273]), .B(p_input[1257]), .Z(n6479) );
  XNOR U6309 ( .A(n6316), .B(n6474), .Z(n6476) );
  XOR U6310 ( .A(n6480), .B(n6481), .Z(n6316) );
  AND U6311 ( .A(n188), .B(n6482), .Z(n6481) );
  XOR U6312 ( .A(p_input[1241]), .B(p_input[1225]), .Z(n6482) );
  XOR U6313 ( .A(n6483), .B(n6484), .Z(n6474) );
  AND U6314 ( .A(n6485), .B(n6486), .Z(n6484) );
  XOR U6315 ( .A(n6483), .B(n6331), .Z(n6486) );
  XNOR U6316 ( .A(p_input[1256]), .B(n6487), .Z(n6331) );
  AND U6317 ( .A(n190), .B(n6488), .Z(n6487) );
  XOR U6318 ( .A(p_input[1272]), .B(p_input[1256]), .Z(n6488) );
  XNOR U6319 ( .A(n6328), .B(n6483), .Z(n6485) );
  XOR U6320 ( .A(n6489), .B(n6490), .Z(n6328) );
  AND U6321 ( .A(n188), .B(n6491), .Z(n6490) );
  XOR U6322 ( .A(p_input[1240]), .B(p_input[1224]), .Z(n6491) );
  XOR U6323 ( .A(n6492), .B(n6493), .Z(n6483) );
  AND U6324 ( .A(n6494), .B(n6495), .Z(n6493) );
  XOR U6325 ( .A(n6492), .B(n6343), .Z(n6495) );
  XNOR U6326 ( .A(p_input[1255]), .B(n6496), .Z(n6343) );
  AND U6327 ( .A(n190), .B(n6497), .Z(n6496) );
  XOR U6328 ( .A(p_input[1271]), .B(p_input[1255]), .Z(n6497) );
  XNOR U6329 ( .A(n6340), .B(n6492), .Z(n6494) );
  XOR U6330 ( .A(n6498), .B(n6499), .Z(n6340) );
  AND U6331 ( .A(n188), .B(n6500), .Z(n6499) );
  XOR U6332 ( .A(p_input[1239]), .B(p_input[1223]), .Z(n6500) );
  XOR U6333 ( .A(n6501), .B(n6502), .Z(n6492) );
  AND U6334 ( .A(n6503), .B(n6504), .Z(n6502) );
  XOR U6335 ( .A(n6501), .B(n6355), .Z(n6504) );
  XNOR U6336 ( .A(p_input[1254]), .B(n6505), .Z(n6355) );
  AND U6337 ( .A(n190), .B(n6506), .Z(n6505) );
  XOR U6338 ( .A(p_input[1270]), .B(p_input[1254]), .Z(n6506) );
  XNOR U6339 ( .A(n6352), .B(n6501), .Z(n6503) );
  XOR U6340 ( .A(n6507), .B(n6508), .Z(n6352) );
  AND U6341 ( .A(n188), .B(n6509), .Z(n6508) );
  XOR U6342 ( .A(p_input[1238]), .B(p_input[1222]), .Z(n6509) );
  XOR U6343 ( .A(n6510), .B(n6511), .Z(n6501) );
  AND U6344 ( .A(n6512), .B(n6513), .Z(n6511) );
  XOR U6345 ( .A(n6510), .B(n6367), .Z(n6513) );
  XNOR U6346 ( .A(p_input[1253]), .B(n6514), .Z(n6367) );
  AND U6347 ( .A(n190), .B(n6515), .Z(n6514) );
  XOR U6348 ( .A(p_input[1269]), .B(p_input[1253]), .Z(n6515) );
  XNOR U6349 ( .A(n6364), .B(n6510), .Z(n6512) );
  XOR U6350 ( .A(n6516), .B(n6517), .Z(n6364) );
  AND U6351 ( .A(n188), .B(n6518), .Z(n6517) );
  XOR U6352 ( .A(p_input[1237]), .B(p_input[1221]), .Z(n6518) );
  XOR U6353 ( .A(n6519), .B(n6520), .Z(n6510) );
  AND U6354 ( .A(n6521), .B(n6522), .Z(n6520) );
  XOR U6355 ( .A(n6519), .B(n6379), .Z(n6522) );
  XNOR U6356 ( .A(p_input[1252]), .B(n6523), .Z(n6379) );
  AND U6357 ( .A(n190), .B(n6524), .Z(n6523) );
  XOR U6358 ( .A(p_input[1268]), .B(p_input[1252]), .Z(n6524) );
  XNOR U6359 ( .A(n6376), .B(n6519), .Z(n6521) );
  XOR U6360 ( .A(n6525), .B(n6526), .Z(n6376) );
  AND U6361 ( .A(n188), .B(n6527), .Z(n6526) );
  XOR U6362 ( .A(p_input[1236]), .B(p_input[1220]), .Z(n6527) );
  XOR U6363 ( .A(n6528), .B(n6529), .Z(n6519) );
  AND U6364 ( .A(n6530), .B(n6531), .Z(n6529) );
  XOR U6365 ( .A(n6528), .B(n6391), .Z(n6531) );
  XNOR U6366 ( .A(p_input[1251]), .B(n6532), .Z(n6391) );
  AND U6367 ( .A(n190), .B(n6533), .Z(n6532) );
  XOR U6368 ( .A(p_input[1267]), .B(p_input[1251]), .Z(n6533) );
  XNOR U6369 ( .A(n6388), .B(n6528), .Z(n6530) );
  XOR U6370 ( .A(n6534), .B(n6535), .Z(n6388) );
  AND U6371 ( .A(n188), .B(n6536), .Z(n6535) );
  XOR U6372 ( .A(p_input[1235]), .B(p_input[1219]), .Z(n6536) );
  XOR U6373 ( .A(n6537), .B(n6538), .Z(n6528) );
  AND U6374 ( .A(n6539), .B(n6540), .Z(n6538) );
  XOR U6375 ( .A(n6403), .B(n6537), .Z(n6540) );
  XNOR U6376 ( .A(p_input[1250]), .B(n6541), .Z(n6403) );
  AND U6377 ( .A(n190), .B(n6542), .Z(n6541) );
  XOR U6378 ( .A(p_input[1266]), .B(p_input[1250]), .Z(n6542) );
  XNOR U6379 ( .A(n6537), .B(n6400), .Z(n6539) );
  XOR U6380 ( .A(n6543), .B(n6544), .Z(n6400) );
  AND U6381 ( .A(n188), .B(n6545), .Z(n6544) );
  XOR U6382 ( .A(p_input[1234]), .B(p_input[1218]), .Z(n6545) );
  XOR U6383 ( .A(n6546), .B(n6547), .Z(n6537) );
  AND U6384 ( .A(n6548), .B(n6549), .Z(n6547) );
  XNOR U6385 ( .A(n6550), .B(n6416), .Z(n6549) );
  XNOR U6386 ( .A(p_input[1249]), .B(n6551), .Z(n6416) );
  AND U6387 ( .A(n190), .B(n6552), .Z(n6551) );
  XNOR U6388 ( .A(p_input[1265]), .B(n6553), .Z(n6552) );
  IV U6389 ( .A(p_input[1249]), .Z(n6553) );
  XNOR U6390 ( .A(n6413), .B(n6546), .Z(n6548) );
  XNOR U6391 ( .A(p_input[1217]), .B(n6554), .Z(n6413) );
  AND U6392 ( .A(n188), .B(n6555), .Z(n6554) );
  XOR U6393 ( .A(p_input[1233]), .B(p_input[1217]), .Z(n6555) );
  IV U6394 ( .A(n6550), .Z(n6546) );
  AND U6395 ( .A(n6421), .B(n6424), .Z(n6550) );
  XOR U6396 ( .A(p_input[1248]), .B(n6556), .Z(n6424) );
  AND U6397 ( .A(n190), .B(n6557), .Z(n6556) );
  XOR U6398 ( .A(p_input[1264]), .B(p_input[1248]), .Z(n6557) );
  XOR U6399 ( .A(n6558), .B(n6559), .Z(n190) );
  AND U6400 ( .A(n6560), .B(n6561), .Z(n6559) );
  XNOR U6401 ( .A(p_input[1279]), .B(n6558), .Z(n6561) );
  XOR U6402 ( .A(n6558), .B(p_input[1263]), .Z(n6560) );
  XOR U6403 ( .A(n6562), .B(n6563), .Z(n6558) );
  AND U6404 ( .A(n6564), .B(n6565), .Z(n6563) );
  XNOR U6405 ( .A(p_input[1278]), .B(n6562), .Z(n6565) );
  XOR U6406 ( .A(n6562), .B(p_input[1262]), .Z(n6564) );
  XOR U6407 ( .A(n6566), .B(n6567), .Z(n6562) );
  AND U6408 ( .A(n6568), .B(n6569), .Z(n6567) );
  XNOR U6409 ( .A(p_input[1277]), .B(n6566), .Z(n6569) );
  XOR U6410 ( .A(n6566), .B(p_input[1261]), .Z(n6568) );
  XOR U6411 ( .A(n6570), .B(n6571), .Z(n6566) );
  AND U6412 ( .A(n6572), .B(n6573), .Z(n6571) );
  XNOR U6413 ( .A(p_input[1276]), .B(n6570), .Z(n6573) );
  XOR U6414 ( .A(n6570), .B(p_input[1260]), .Z(n6572) );
  XOR U6415 ( .A(n6574), .B(n6575), .Z(n6570) );
  AND U6416 ( .A(n6576), .B(n6577), .Z(n6575) );
  XNOR U6417 ( .A(p_input[1275]), .B(n6574), .Z(n6577) );
  XOR U6418 ( .A(n6574), .B(p_input[1259]), .Z(n6576) );
  XOR U6419 ( .A(n6578), .B(n6579), .Z(n6574) );
  AND U6420 ( .A(n6580), .B(n6581), .Z(n6579) );
  XNOR U6421 ( .A(p_input[1274]), .B(n6578), .Z(n6581) );
  XOR U6422 ( .A(n6578), .B(p_input[1258]), .Z(n6580) );
  XOR U6423 ( .A(n6582), .B(n6583), .Z(n6578) );
  AND U6424 ( .A(n6584), .B(n6585), .Z(n6583) );
  XNOR U6425 ( .A(p_input[1273]), .B(n6582), .Z(n6585) );
  XOR U6426 ( .A(n6582), .B(p_input[1257]), .Z(n6584) );
  XOR U6427 ( .A(n6586), .B(n6587), .Z(n6582) );
  AND U6428 ( .A(n6588), .B(n6589), .Z(n6587) );
  XNOR U6429 ( .A(p_input[1272]), .B(n6586), .Z(n6589) );
  XOR U6430 ( .A(n6586), .B(p_input[1256]), .Z(n6588) );
  XOR U6431 ( .A(n6590), .B(n6591), .Z(n6586) );
  AND U6432 ( .A(n6592), .B(n6593), .Z(n6591) );
  XNOR U6433 ( .A(p_input[1271]), .B(n6590), .Z(n6593) );
  XOR U6434 ( .A(n6590), .B(p_input[1255]), .Z(n6592) );
  XOR U6435 ( .A(n6594), .B(n6595), .Z(n6590) );
  AND U6436 ( .A(n6596), .B(n6597), .Z(n6595) );
  XNOR U6437 ( .A(p_input[1270]), .B(n6594), .Z(n6597) );
  XOR U6438 ( .A(n6594), .B(p_input[1254]), .Z(n6596) );
  XOR U6439 ( .A(n6598), .B(n6599), .Z(n6594) );
  AND U6440 ( .A(n6600), .B(n6601), .Z(n6599) );
  XNOR U6441 ( .A(p_input[1269]), .B(n6598), .Z(n6601) );
  XOR U6442 ( .A(n6598), .B(p_input[1253]), .Z(n6600) );
  XOR U6443 ( .A(n6602), .B(n6603), .Z(n6598) );
  AND U6444 ( .A(n6604), .B(n6605), .Z(n6603) );
  XNOR U6445 ( .A(p_input[1268]), .B(n6602), .Z(n6605) );
  XOR U6446 ( .A(n6602), .B(p_input[1252]), .Z(n6604) );
  XOR U6447 ( .A(n6606), .B(n6607), .Z(n6602) );
  AND U6448 ( .A(n6608), .B(n6609), .Z(n6607) );
  XNOR U6449 ( .A(p_input[1267]), .B(n6606), .Z(n6609) );
  XOR U6450 ( .A(n6606), .B(p_input[1251]), .Z(n6608) );
  XOR U6451 ( .A(n6610), .B(n6611), .Z(n6606) );
  AND U6452 ( .A(n6612), .B(n6613), .Z(n6611) );
  XNOR U6453 ( .A(p_input[1266]), .B(n6610), .Z(n6613) );
  XOR U6454 ( .A(n6610), .B(p_input[1250]), .Z(n6612) );
  XNOR U6455 ( .A(n6614), .B(n6615), .Z(n6610) );
  AND U6456 ( .A(n6616), .B(n6617), .Z(n6615) );
  XOR U6457 ( .A(p_input[1265]), .B(n6614), .Z(n6617) );
  XNOR U6458 ( .A(p_input[1249]), .B(n6614), .Z(n6616) );
  AND U6459 ( .A(p_input[1264]), .B(n6618), .Z(n6614) );
  IV U6460 ( .A(p_input[1248]), .Z(n6618) );
  XNOR U6461 ( .A(p_input[1216]), .B(n6619), .Z(n6421) );
  AND U6462 ( .A(n188), .B(n6620), .Z(n6619) );
  XOR U6463 ( .A(p_input[1232]), .B(p_input[1216]), .Z(n6620) );
  XOR U6464 ( .A(n6621), .B(n6622), .Z(n188) );
  AND U6465 ( .A(n6623), .B(n6624), .Z(n6622) );
  XNOR U6466 ( .A(p_input[1247]), .B(n6621), .Z(n6624) );
  XOR U6467 ( .A(n6621), .B(p_input[1231]), .Z(n6623) );
  XOR U6468 ( .A(n6625), .B(n6626), .Z(n6621) );
  AND U6469 ( .A(n6627), .B(n6628), .Z(n6626) );
  XNOR U6470 ( .A(p_input[1246]), .B(n6625), .Z(n6628) );
  XNOR U6471 ( .A(n6625), .B(n6435), .Z(n6627) );
  IV U6472 ( .A(p_input[1230]), .Z(n6435) );
  XOR U6473 ( .A(n6629), .B(n6630), .Z(n6625) );
  AND U6474 ( .A(n6631), .B(n6632), .Z(n6630) );
  XNOR U6475 ( .A(p_input[1245]), .B(n6629), .Z(n6632) );
  XNOR U6476 ( .A(n6629), .B(n6444), .Z(n6631) );
  IV U6477 ( .A(p_input[1229]), .Z(n6444) );
  XOR U6478 ( .A(n6633), .B(n6634), .Z(n6629) );
  AND U6479 ( .A(n6635), .B(n6636), .Z(n6634) );
  XNOR U6480 ( .A(p_input[1244]), .B(n6633), .Z(n6636) );
  XNOR U6481 ( .A(n6633), .B(n6453), .Z(n6635) );
  IV U6482 ( .A(p_input[1228]), .Z(n6453) );
  XOR U6483 ( .A(n6637), .B(n6638), .Z(n6633) );
  AND U6484 ( .A(n6639), .B(n6640), .Z(n6638) );
  XNOR U6485 ( .A(p_input[1243]), .B(n6637), .Z(n6640) );
  XNOR U6486 ( .A(n6637), .B(n6462), .Z(n6639) );
  IV U6487 ( .A(p_input[1227]), .Z(n6462) );
  XOR U6488 ( .A(n6641), .B(n6642), .Z(n6637) );
  AND U6489 ( .A(n6643), .B(n6644), .Z(n6642) );
  XNOR U6490 ( .A(p_input[1242]), .B(n6641), .Z(n6644) );
  XNOR U6491 ( .A(n6641), .B(n6471), .Z(n6643) );
  IV U6492 ( .A(p_input[1226]), .Z(n6471) );
  XOR U6493 ( .A(n6645), .B(n6646), .Z(n6641) );
  AND U6494 ( .A(n6647), .B(n6648), .Z(n6646) );
  XNOR U6495 ( .A(p_input[1241]), .B(n6645), .Z(n6648) );
  XNOR U6496 ( .A(n6645), .B(n6480), .Z(n6647) );
  IV U6497 ( .A(p_input[1225]), .Z(n6480) );
  XOR U6498 ( .A(n6649), .B(n6650), .Z(n6645) );
  AND U6499 ( .A(n6651), .B(n6652), .Z(n6650) );
  XNOR U6500 ( .A(p_input[1240]), .B(n6649), .Z(n6652) );
  XNOR U6501 ( .A(n6649), .B(n6489), .Z(n6651) );
  IV U6502 ( .A(p_input[1224]), .Z(n6489) );
  XOR U6503 ( .A(n6653), .B(n6654), .Z(n6649) );
  AND U6504 ( .A(n6655), .B(n6656), .Z(n6654) );
  XNOR U6505 ( .A(p_input[1239]), .B(n6653), .Z(n6656) );
  XNOR U6506 ( .A(n6653), .B(n6498), .Z(n6655) );
  IV U6507 ( .A(p_input[1223]), .Z(n6498) );
  XOR U6508 ( .A(n6657), .B(n6658), .Z(n6653) );
  AND U6509 ( .A(n6659), .B(n6660), .Z(n6658) );
  XNOR U6510 ( .A(p_input[1238]), .B(n6657), .Z(n6660) );
  XNOR U6511 ( .A(n6657), .B(n6507), .Z(n6659) );
  IV U6512 ( .A(p_input[1222]), .Z(n6507) );
  XOR U6513 ( .A(n6661), .B(n6662), .Z(n6657) );
  AND U6514 ( .A(n6663), .B(n6664), .Z(n6662) );
  XNOR U6515 ( .A(p_input[1237]), .B(n6661), .Z(n6664) );
  XNOR U6516 ( .A(n6661), .B(n6516), .Z(n6663) );
  IV U6517 ( .A(p_input[1221]), .Z(n6516) );
  XOR U6518 ( .A(n6665), .B(n6666), .Z(n6661) );
  AND U6519 ( .A(n6667), .B(n6668), .Z(n6666) );
  XNOR U6520 ( .A(p_input[1236]), .B(n6665), .Z(n6668) );
  XNOR U6521 ( .A(n6665), .B(n6525), .Z(n6667) );
  IV U6522 ( .A(p_input[1220]), .Z(n6525) );
  XOR U6523 ( .A(n6669), .B(n6670), .Z(n6665) );
  AND U6524 ( .A(n6671), .B(n6672), .Z(n6670) );
  XNOR U6525 ( .A(p_input[1235]), .B(n6669), .Z(n6672) );
  XNOR U6526 ( .A(n6669), .B(n6534), .Z(n6671) );
  IV U6527 ( .A(p_input[1219]), .Z(n6534) );
  XOR U6528 ( .A(n6673), .B(n6674), .Z(n6669) );
  AND U6529 ( .A(n6675), .B(n6676), .Z(n6674) );
  XNOR U6530 ( .A(p_input[1234]), .B(n6673), .Z(n6676) );
  XNOR U6531 ( .A(n6673), .B(n6543), .Z(n6675) );
  IV U6532 ( .A(p_input[1218]), .Z(n6543) );
  XNOR U6533 ( .A(n6677), .B(n6678), .Z(n6673) );
  AND U6534 ( .A(n6679), .B(n6680), .Z(n6678) );
  XOR U6535 ( .A(p_input[1233]), .B(n6677), .Z(n6680) );
  XNOR U6536 ( .A(p_input[1217]), .B(n6677), .Z(n6679) );
  AND U6537 ( .A(p_input[1232]), .B(n6681), .Z(n6677) );
  IV U6538 ( .A(p_input[1216]), .Z(n6681) );
  XOR U6539 ( .A(n6682), .B(n6683), .Z(n6240) );
  AND U6540 ( .A(n264), .B(n6684), .Z(n6683) );
  XNOR U6541 ( .A(n6685), .B(n6682), .Z(n6684) );
  XOR U6542 ( .A(n6686), .B(n6687), .Z(n264) );
  AND U6543 ( .A(n6688), .B(n6689), .Z(n6687) );
  XNOR U6544 ( .A(n6250), .B(n6686), .Z(n6689) );
  AND U6545 ( .A(p_input[1215]), .B(p_input[1199]), .Z(n6250) );
  XOR U6546 ( .A(n6686), .B(n6251), .Z(n6688) );
  AND U6547 ( .A(p_input[1183]), .B(p_input[1167]), .Z(n6251) );
  XOR U6548 ( .A(n6690), .B(n6691), .Z(n6686) );
  AND U6549 ( .A(n6692), .B(n6693), .Z(n6691) );
  XOR U6550 ( .A(n6690), .B(n6263), .Z(n6693) );
  XNOR U6551 ( .A(p_input[1198]), .B(n6694), .Z(n6263) );
  AND U6552 ( .A(n194), .B(n6695), .Z(n6694) );
  XOR U6553 ( .A(p_input[1214]), .B(p_input[1198]), .Z(n6695) );
  XNOR U6554 ( .A(n6260), .B(n6690), .Z(n6692) );
  XOR U6555 ( .A(n6696), .B(n6697), .Z(n6260) );
  AND U6556 ( .A(n191), .B(n6698), .Z(n6697) );
  XOR U6557 ( .A(p_input[1182]), .B(p_input[1166]), .Z(n6698) );
  XOR U6558 ( .A(n6699), .B(n6700), .Z(n6690) );
  AND U6559 ( .A(n6701), .B(n6702), .Z(n6700) );
  XOR U6560 ( .A(n6699), .B(n6275), .Z(n6702) );
  XNOR U6561 ( .A(p_input[1197]), .B(n6703), .Z(n6275) );
  AND U6562 ( .A(n194), .B(n6704), .Z(n6703) );
  XOR U6563 ( .A(p_input[1213]), .B(p_input[1197]), .Z(n6704) );
  XNOR U6564 ( .A(n6272), .B(n6699), .Z(n6701) );
  XOR U6565 ( .A(n6705), .B(n6706), .Z(n6272) );
  AND U6566 ( .A(n191), .B(n6707), .Z(n6706) );
  XOR U6567 ( .A(p_input[1181]), .B(p_input[1165]), .Z(n6707) );
  XOR U6568 ( .A(n6708), .B(n6709), .Z(n6699) );
  AND U6569 ( .A(n6710), .B(n6711), .Z(n6709) );
  XOR U6570 ( .A(n6708), .B(n6287), .Z(n6711) );
  XNOR U6571 ( .A(p_input[1196]), .B(n6712), .Z(n6287) );
  AND U6572 ( .A(n194), .B(n6713), .Z(n6712) );
  XOR U6573 ( .A(p_input[1212]), .B(p_input[1196]), .Z(n6713) );
  XNOR U6574 ( .A(n6284), .B(n6708), .Z(n6710) );
  XOR U6575 ( .A(n6714), .B(n6715), .Z(n6284) );
  AND U6576 ( .A(n191), .B(n6716), .Z(n6715) );
  XOR U6577 ( .A(p_input[1180]), .B(p_input[1164]), .Z(n6716) );
  XOR U6578 ( .A(n6717), .B(n6718), .Z(n6708) );
  AND U6579 ( .A(n6719), .B(n6720), .Z(n6718) );
  XOR U6580 ( .A(n6717), .B(n6299), .Z(n6720) );
  XNOR U6581 ( .A(p_input[1195]), .B(n6721), .Z(n6299) );
  AND U6582 ( .A(n194), .B(n6722), .Z(n6721) );
  XOR U6583 ( .A(p_input[1211]), .B(p_input[1195]), .Z(n6722) );
  XNOR U6584 ( .A(n6296), .B(n6717), .Z(n6719) );
  XOR U6585 ( .A(n6723), .B(n6724), .Z(n6296) );
  AND U6586 ( .A(n191), .B(n6725), .Z(n6724) );
  XOR U6587 ( .A(p_input[1179]), .B(p_input[1163]), .Z(n6725) );
  XOR U6588 ( .A(n6726), .B(n6727), .Z(n6717) );
  AND U6589 ( .A(n6728), .B(n6729), .Z(n6727) );
  XOR U6590 ( .A(n6726), .B(n6311), .Z(n6729) );
  XNOR U6591 ( .A(p_input[1194]), .B(n6730), .Z(n6311) );
  AND U6592 ( .A(n194), .B(n6731), .Z(n6730) );
  XOR U6593 ( .A(p_input[1210]), .B(p_input[1194]), .Z(n6731) );
  XNOR U6594 ( .A(n6308), .B(n6726), .Z(n6728) );
  XOR U6595 ( .A(n6732), .B(n6733), .Z(n6308) );
  AND U6596 ( .A(n191), .B(n6734), .Z(n6733) );
  XOR U6597 ( .A(p_input[1178]), .B(p_input[1162]), .Z(n6734) );
  XOR U6598 ( .A(n6735), .B(n6736), .Z(n6726) );
  AND U6599 ( .A(n6737), .B(n6738), .Z(n6736) );
  XOR U6600 ( .A(n6735), .B(n6323), .Z(n6738) );
  XNOR U6601 ( .A(p_input[1193]), .B(n6739), .Z(n6323) );
  AND U6602 ( .A(n194), .B(n6740), .Z(n6739) );
  XOR U6603 ( .A(p_input[1209]), .B(p_input[1193]), .Z(n6740) );
  XNOR U6604 ( .A(n6320), .B(n6735), .Z(n6737) );
  XOR U6605 ( .A(n6741), .B(n6742), .Z(n6320) );
  AND U6606 ( .A(n191), .B(n6743), .Z(n6742) );
  XOR U6607 ( .A(p_input[1177]), .B(p_input[1161]), .Z(n6743) );
  XOR U6608 ( .A(n6744), .B(n6745), .Z(n6735) );
  AND U6609 ( .A(n6746), .B(n6747), .Z(n6745) );
  XOR U6610 ( .A(n6744), .B(n6335), .Z(n6747) );
  XNOR U6611 ( .A(p_input[1192]), .B(n6748), .Z(n6335) );
  AND U6612 ( .A(n194), .B(n6749), .Z(n6748) );
  XOR U6613 ( .A(p_input[1208]), .B(p_input[1192]), .Z(n6749) );
  XNOR U6614 ( .A(n6332), .B(n6744), .Z(n6746) );
  XOR U6615 ( .A(n6750), .B(n6751), .Z(n6332) );
  AND U6616 ( .A(n191), .B(n6752), .Z(n6751) );
  XOR U6617 ( .A(p_input[1176]), .B(p_input[1160]), .Z(n6752) );
  XOR U6618 ( .A(n6753), .B(n6754), .Z(n6744) );
  AND U6619 ( .A(n6755), .B(n6756), .Z(n6754) );
  XOR U6620 ( .A(n6753), .B(n6347), .Z(n6756) );
  XNOR U6621 ( .A(p_input[1191]), .B(n6757), .Z(n6347) );
  AND U6622 ( .A(n194), .B(n6758), .Z(n6757) );
  XOR U6623 ( .A(p_input[1207]), .B(p_input[1191]), .Z(n6758) );
  XNOR U6624 ( .A(n6344), .B(n6753), .Z(n6755) );
  XOR U6625 ( .A(n6759), .B(n6760), .Z(n6344) );
  AND U6626 ( .A(n191), .B(n6761), .Z(n6760) );
  XOR U6627 ( .A(p_input[1175]), .B(p_input[1159]), .Z(n6761) );
  XOR U6628 ( .A(n6762), .B(n6763), .Z(n6753) );
  AND U6629 ( .A(n6764), .B(n6765), .Z(n6763) );
  XOR U6630 ( .A(n6762), .B(n6359), .Z(n6765) );
  XNOR U6631 ( .A(p_input[1190]), .B(n6766), .Z(n6359) );
  AND U6632 ( .A(n194), .B(n6767), .Z(n6766) );
  XOR U6633 ( .A(p_input[1206]), .B(p_input[1190]), .Z(n6767) );
  XNOR U6634 ( .A(n6356), .B(n6762), .Z(n6764) );
  XOR U6635 ( .A(n6768), .B(n6769), .Z(n6356) );
  AND U6636 ( .A(n191), .B(n6770), .Z(n6769) );
  XOR U6637 ( .A(p_input[1174]), .B(p_input[1158]), .Z(n6770) );
  XOR U6638 ( .A(n6771), .B(n6772), .Z(n6762) );
  AND U6639 ( .A(n6773), .B(n6774), .Z(n6772) );
  XOR U6640 ( .A(n6771), .B(n6371), .Z(n6774) );
  XNOR U6641 ( .A(p_input[1189]), .B(n6775), .Z(n6371) );
  AND U6642 ( .A(n194), .B(n6776), .Z(n6775) );
  XOR U6643 ( .A(p_input[1205]), .B(p_input[1189]), .Z(n6776) );
  XNOR U6644 ( .A(n6368), .B(n6771), .Z(n6773) );
  XOR U6645 ( .A(n6777), .B(n6778), .Z(n6368) );
  AND U6646 ( .A(n191), .B(n6779), .Z(n6778) );
  XOR U6647 ( .A(p_input[1173]), .B(p_input[1157]), .Z(n6779) );
  XOR U6648 ( .A(n6780), .B(n6781), .Z(n6771) );
  AND U6649 ( .A(n6782), .B(n6783), .Z(n6781) );
  XOR U6650 ( .A(n6780), .B(n6383), .Z(n6783) );
  XNOR U6651 ( .A(p_input[1188]), .B(n6784), .Z(n6383) );
  AND U6652 ( .A(n194), .B(n6785), .Z(n6784) );
  XOR U6653 ( .A(p_input[1204]), .B(p_input[1188]), .Z(n6785) );
  XNOR U6654 ( .A(n6380), .B(n6780), .Z(n6782) );
  XOR U6655 ( .A(n6786), .B(n6787), .Z(n6380) );
  AND U6656 ( .A(n191), .B(n6788), .Z(n6787) );
  XOR U6657 ( .A(p_input[1172]), .B(p_input[1156]), .Z(n6788) );
  XOR U6658 ( .A(n6789), .B(n6790), .Z(n6780) );
  AND U6659 ( .A(n6791), .B(n6792), .Z(n6790) );
  XOR U6660 ( .A(n6789), .B(n6395), .Z(n6792) );
  XNOR U6661 ( .A(p_input[1187]), .B(n6793), .Z(n6395) );
  AND U6662 ( .A(n194), .B(n6794), .Z(n6793) );
  XOR U6663 ( .A(p_input[1203]), .B(p_input[1187]), .Z(n6794) );
  XNOR U6664 ( .A(n6392), .B(n6789), .Z(n6791) );
  XOR U6665 ( .A(n6795), .B(n6796), .Z(n6392) );
  AND U6666 ( .A(n191), .B(n6797), .Z(n6796) );
  XOR U6667 ( .A(p_input[1171]), .B(p_input[1155]), .Z(n6797) );
  XOR U6668 ( .A(n6798), .B(n6799), .Z(n6789) );
  AND U6669 ( .A(n6800), .B(n6801), .Z(n6799) );
  XOR U6670 ( .A(n6407), .B(n6798), .Z(n6801) );
  XNOR U6671 ( .A(p_input[1186]), .B(n6802), .Z(n6407) );
  AND U6672 ( .A(n194), .B(n6803), .Z(n6802) );
  XOR U6673 ( .A(p_input[1202]), .B(p_input[1186]), .Z(n6803) );
  XNOR U6674 ( .A(n6798), .B(n6404), .Z(n6800) );
  XOR U6675 ( .A(n6804), .B(n6805), .Z(n6404) );
  AND U6676 ( .A(n191), .B(n6806), .Z(n6805) );
  XOR U6677 ( .A(p_input[1170]), .B(p_input[1154]), .Z(n6806) );
  XOR U6678 ( .A(n6807), .B(n6808), .Z(n6798) );
  AND U6679 ( .A(n6809), .B(n6810), .Z(n6808) );
  XNOR U6680 ( .A(n6811), .B(n6420), .Z(n6810) );
  XNOR U6681 ( .A(p_input[1185]), .B(n6812), .Z(n6420) );
  AND U6682 ( .A(n194), .B(n6813), .Z(n6812) );
  XNOR U6683 ( .A(p_input[1201]), .B(n6814), .Z(n6813) );
  IV U6684 ( .A(p_input[1185]), .Z(n6814) );
  XNOR U6685 ( .A(n6417), .B(n6807), .Z(n6809) );
  XNOR U6686 ( .A(p_input[1153]), .B(n6815), .Z(n6417) );
  AND U6687 ( .A(n191), .B(n6816), .Z(n6815) );
  XOR U6688 ( .A(p_input[1169]), .B(p_input[1153]), .Z(n6816) );
  IV U6689 ( .A(n6811), .Z(n6807) );
  AND U6690 ( .A(n6682), .B(n6685), .Z(n6811) );
  XOR U6691 ( .A(p_input[1184]), .B(n6817), .Z(n6685) );
  AND U6692 ( .A(n194), .B(n6818), .Z(n6817) );
  XOR U6693 ( .A(p_input[1200]), .B(p_input[1184]), .Z(n6818) );
  XOR U6694 ( .A(n6819), .B(n6820), .Z(n194) );
  AND U6695 ( .A(n6821), .B(n6822), .Z(n6820) );
  XNOR U6696 ( .A(p_input[1215]), .B(n6819), .Z(n6822) );
  XOR U6697 ( .A(n6819), .B(p_input[1199]), .Z(n6821) );
  XOR U6698 ( .A(n6823), .B(n6824), .Z(n6819) );
  AND U6699 ( .A(n6825), .B(n6826), .Z(n6824) );
  XNOR U6700 ( .A(p_input[1214]), .B(n6823), .Z(n6826) );
  XOR U6701 ( .A(n6823), .B(p_input[1198]), .Z(n6825) );
  XOR U6702 ( .A(n6827), .B(n6828), .Z(n6823) );
  AND U6703 ( .A(n6829), .B(n6830), .Z(n6828) );
  XNOR U6704 ( .A(p_input[1213]), .B(n6827), .Z(n6830) );
  XOR U6705 ( .A(n6827), .B(p_input[1197]), .Z(n6829) );
  XOR U6706 ( .A(n6831), .B(n6832), .Z(n6827) );
  AND U6707 ( .A(n6833), .B(n6834), .Z(n6832) );
  XNOR U6708 ( .A(p_input[1212]), .B(n6831), .Z(n6834) );
  XOR U6709 ( .A(n6831), .B(p_input[1196]), .Z(n6833) );
  XOR U6710 ( .A(n6835), .B(n6836), .Z(n6831) );
  AND U6711 ( .A(n6837), .B(n6838), .Z(n6836) );
  XNOR U6712 ( .A(p_input[1211]), .B(n6835), .Z(n6838) );
  XOR U6713 ( .A(n6835), .B(p_input[1195]), .Z(n6837) );
  XOR U6714 ( .A(n6839), .B(n6840), .Z(n6835) );
  AND U6715 ( .A(n6841), .B(n6842), .Z(n6840) );
  XNOR U6716 ( .A(p_input[1210]), .B(n6839), .Z(n6842) );
  XOR U6717 ( .A(n6839), .B(p_input[1194]), .Z(n6841) );
  XOR U6718 ( .A(n6843), .B(n6844), .Z(n6839) );
  AND U6719 ( .A(n6845), .B(n6846), .Z(n6844) );
  XNOR U6720 ( .A(p_input[1209]), .B(n6843), .Z(n6846) );
  XOR U6721 ( .A(n6843), .B(p_input[1193]), .Z(n6845) );
  XOR U6722 ( .A(n6847), .B(n6848), .Z(n6843) );
  AND U6723 ( .A(n6849), .B(n6850), .Z(n6848) );
  XNOR U6724 ( .A(p_input[1208]), .B(n6847), .Z(n6850) );
  XOR U6725 ( .A(n6847), .B(p_input[1192]), .Z(n6849) );
  XOR U6726 ( .A(n6851), .B(n6852), .Z(n6847) );
  AND U6727 ( .A(n6853), .B(n6854), .Z(n6852) );
  XNOR U6728 ( .A(p_input[1207]), .B(n6851), .Z(n6854) );
  XOR U6729 ( .A(n6851), .B(p_input[1191]), .Z(n6853) );
  XOR U6730 ( .A(n6855), .B(n6856), .Z(n6851) );
  AND U6731 ( .A(n6857), .B(n6858), .Z(n6856) );
  XNOR U6732 ( .A(p_input[1206]), .B(n6855), .Z(n6858) );
  XOR U6733 ( .A(n6855), .B(p_input[1190]), .Z(n6857) );
  XOR U6734 ( .A(n6859), .B(n6860), .Z(n6855) );
  AND U6735 ( .A(n6861), .B(n6862), .Z(n6860) );
  XNOR U6736 ( .A(p_input[1205]), .B(n6859), .Z(n6862) );
  XOR U6737 ( .A(n6859), .B(p_input[1189]), .Z(n6861) );
  XOR U6738 ( .A(n6863), .B(n6864), .Z(n6859) );
  AND U6739 ( .A(n6865), .B(n6866), .Z(n6864) );
  XNOR U6740 ( .A(p_input[1204]), .B(n6863), .Z(n6866) );
  XOR U6741 ( .A(n6863), .B(p_input[1188]), .Z(n6865) );
  XOR U6742 ( .A(n6867), .B(n6868), .Z(n6863) );
  AND U6743 ( .A(n6869), .B(n6870), .Z(n6868) );
  XNOR U6744 ( .A(p_input[1203]), .B(n6867), .Z(n6870) );
  XOR U6745 ( .A(n6867), .B(p_input[1187]), .Z(n6869) );
  XOR U6746 ( .A(n6871), .B(n6872), .Z(n6867) );
  AND U6747 ( .A(n6873), .B(n6874), .Z(n6872) );
  XNOR U6748 ( .A(p_input[1202]), .B(n6871), .Z(n6874) );
  XOR U6749 ( .A(n6871), .B(p_input[1186]), .Z(n6873) );
  XNOR U6750 ( .A(n6875), .B(n6876), .Z(n6871) );
  AND U6751 ( .A(n6877), .B(n6878), .Z(n6876) );
  XOR U6752 ( .A(p_input[1201]), .B(n6875), .Z(n6878) );
  XNOR U6753 ( .A(p_input[1185]), .B(n6875), .Z(n6877) );
  AND U6754 ( .A(p_input[1200]), .B(n6879), .Z(n6875) );
  IV U6755 ( .A(p_input[1184]), .Z(n6879) );
  XNOR U6756 ( .A(p_input[1152]), .B(n6880), .Z(n6682) );
  AND U6757 ( .A(n191), .B(n6881), .Z(n6880) );
  XOR U6758 ( .A(p_input[1168]), .B(p_input[1152]), .Z(n6881) );
  XOR U6759 ( .A(n6882), .B(n6883), .Z(n191) );
  AND U6760 ( .A(n6884), .B(n6885), .Z(n6883) );
  XNOR U6761 ( .A(p_input[1183]), .B(n6882), .Z(n6885) );
  XOR U6762 ( .A(n6882), .B(p_input[1167]), .Z(n6884) );
  XOR U6763 ( .A(n6886), .B(n6887), .Z(n6882) );
  AND U6764 ( .A(n6888), .B(n6889), .Z(n6887) );
  XNOR U6765 ( .A(p_input[1182]), .B(n6886), .Z(n6889) );
  XNOR U6766 ( .A(n6886), .B(n6696), .Z(n6888) );
  IV U6767 ( .A(p_input[1166]), .Z(n6696) );
  XOR U6768 ( .A(n6890), .B(n6891), .Z(n6886) );
  AND U6769 ( .A(n6892), .B(n6893), .Z(n6891) );
  XNOR U6770 ( .A(p_input[1181]), .B(n6890), .Z(n6893) );
  XNOR U6771 ( .A(n6890), .B(n6705), .Z(n6892) );
  IV U6772 ( .A(p_input[1165]), .Z(n6705) );
  XOR U6773 ( .A(n6894), .B(n6895), .Z(n6890) );
  AND U6774 ( .A(n6896), .B(n6897), .Z(n6895) );
  XNOR U6775 ( .A(p_input[1180]), .B(n6894), .Z(n6897) );
  XNOR U6776 ( .A(n6894), .B(n6714), .Z(n6896) );
  IV U6777 ( .A(p_input[1164]), .Z(n6714) );
  XOR U6778 ( .A(n6898), .B(n6899), .Z(n6894) );
  AND U6779 ( .A(n6900), .B(n6901), .Z(n6899) );
  XNOR U6780 ( .A(p_input[1179]), .B(n6898), .Z(n6901) );
  XNOR U6781 ( .A(n6898), .B(n6723), .Z(n6900) );
  IV U6782 ( .A(p_input[1163]), .Z(n6723) );
  XOR U6783 ( .A(n6902), .B(n6903), .Z(n6898) );
  AND U6784 ( .A(n6904), .B(n6905), .Z(n6903) );
  XNOR U6785 ( .A(p_input[1178]), .B(n6902), .Z(n6905) );
  XNOR U6786 ( .A(n6902), .B(n6732), .Z(n6904) );
  IV U6787 ( .A(p_input[1162]), .Z(n6732) );
  XOR U6788 ( .A(n6906), .B(n6907), .Z(n6902) );
  AND U6789 ( .A(n6908), .B(n6909), .Z(n6907) );
  XNOR U6790 ( .A(p_input[1177]), .B(n6906), .Z(n6909) );
  XNOR U6791 ( .A(n6906), .B(n6741), .Z(n6908) );
  IV U6792 ( .A(p_input[1161]), .Z(n6741) );
  XOR U6793 ( .A(n6910), .B(n6911), .Z(n6906) );
  AND U6794 ( .A(n6912), .B(n6913), .Z(n6911) );
  XNOR U6795 ( .A(p_input[1176]), .B(n6910), .Z(n6913) );
  XNOR U6796 ( .A(n6910), .B(n6750), .Z(n6912) );
  IV U6797 ( .A(p_input[1160]), .Z(n6750) );
  XOR U6798 ( .A(n6914), .B(n6915), .Z(n6910) );
  AND U6799 ( .A(n6916), .B(n6917), .Z(n6915) );
  XNOR U6800 ( .A(p_input[1175]), .B(n6914), .Z(n6917) );
  XNOR U6801 ( .A(n6914), .B(n6759), .Z(n6916) );
  IV U6802 ( .A(p_input[1159]), .Z(n6759) );
  XOR U6803 ( .A(n6918), .B(n6919), .Z(n6914) );
  AND U6804 ( .A(n6920), .B(n6921), .Z(n6919) );
  XNOR U6805 ( .A(p_input[1174]), .B(n6918), .Z(n6921) );
  XNOR U6806 ( .A(n6918), .B(n6768), .Z(n6920) );
  IV U6807 ( .A(p_input[1158]), .Z(n6768) );
  XOR U6808 ( .A(n6922), .B(n6923), .Z(n6918) );
  AND U6809 ( .A(n6924), .B(n6925), .Z(n6923) );
  XNOR U6810 ( .A(p_input[1173]), .B(n6922), .Z(n6925) );
  XNOR U6811 ( .A(n6922), .B(n6777), .Z(n6924) );
  IV U6812 ( .A(p_input[1157]), .Z(n6777) );
  XOR U6813 ( .A(n6926), .B(n6927), .Z(n6922) );
  AND U6814 ( .A(n6928), .B(n6929), .Z(n6927) );
  XNOR U6815 ( .A(p_input[1172]), .B(n6926), .Z(n6929) );
  XNOR U6816 ( .A(n6926), .B(n6786), .Z(n6928) );
  IV U6817 ( .A(p_input[1156]), .Z(n6786) );
  XOR U6818 ( .A(n6930), .B(n6931), .Z(n6926) );
  AND U6819 ( .A(n6932), .B(n6933), .Z(n6931) );
  XNOR U6820 ( .A(p_input[1171]), .B(n6930), .Z(n6933) );
  XNOR U6821 ( .A(n6930), .B(n6795), .Z(n6932) );
  IV U6822 ( .A(p_input[1155]), .Z(n6795) );
  XOR U6823 ( .A(n6934), .B(n6935), .Z(n6930) );
  AND U6824 ( .A(n6936), .B(n6937), .Z(n6935) );
  XNOR U6825 ( .A(p_input[1170]), .B(n6934), .Z(n6937) );
  XNOR U6826 ( .A(n6934), .B(n6804), .Z(n6936) );
  IV U6827 ( .A(p_input[1154]), .Z(n6804) );
  XNOR U6828 ( .A(n6938), .B(n6939), .Z(n6934) );
  AND U6829 ( .A(n6940), .B(n6941), .Z(n6939) );
  XOR U6830 ( .A(p_input[1169]), .B(n6938), .Z(n6941) );
  XNOR U6831 ( .A(p_input[1153]), .B(n6938), .Z(n6940) );
  AND U6832 ( .A(p_input[1168]), .B(n6942), .Z(n6938) );
  IV U6833 ( .A(p_input[1152]), .Z(n6942) );
  XOR U6834 ( .A(n6943), .B(n6944), .Z(n6058) );
  AND U6835 ( .A(n423), .B(n6945), .Z(n6944) );
  XNOR U6836 ( .A(n6946), .B(n6943), .Z(n6945) );
  XOR U6837 ( .A(n6947), .B(n6948), .Z(n423) );
  AND U6838 ( .A(n6949), .B(n6950), .Z(n6948) );
  XNOR U6839 ( .A(n6070), .B(n6947), .Z(n6950) );
  AND U6840 ( .A(n6951), .B(n6952), .Z(n6070) );
  XOR U6841 ( .A(n6947), .B(n6069), .Z(n6949) );
  AND U6842 ( .A(n6953), .B(n6954), .Z(n6069) );
  XOR U6843 ( .A(n6955), .B(n6956), .Z(n6947) );
  AND U6844 ( .A(n6957), .B(n6958), .Z(n6956) );
  XOR U6845 ( .A(n6955), .B(n6082), .Z(n6958) );
  XOR U6846 ( .A(n6959), .B(n6960), .Z(n6082) );
  AND U6847 ( .A(n270), .B(n6961), .Z(n6960) );
  XOR U6848 ( .A(n6962), .B(n6959), .Z(n6961) );
  XNOR U6849 ( .A(n6079), .B(n6955), .Z(n6957) );
  XOR U6850 ( .A(n6963), .B(n6964), .Z(n6079) );
  AND U6851 ( .A(n267), .B(n6965), .Z(n6964) );
  XOR U6852 ( .A(n6966), .B(n6963), .Z(n6965) );
  XOR U6853 ( .A(n6967), .B(n6968), .Z(n6955) );
  AND U6854 ( .A(n6969), .B(n6970), .Z(n6968) );
  XOR U6855 ( .A(n6967), .B(n6094), .Z(n6970) );
  XOR U6856 ( .A(n6971), .B(n6972), .Z(n6094) );
  AND U6857 ( .A(n270), .B(n6973), .Z(n6972) );
  XOR U6858 ( .A(n6974), .B(n6971), .Z(n6973) );
  XNOR U6859 ( .A(n6091), .B(n6967), .Z(n6969) );
  XOR U6860 ( .A(n6975), .B(n6976), .Z(n6091) );
  AND U6861 ( .A(n267), .B(n6977), .Z(n6976) );
  XOR U6862 ( .A(n6978), .B(n6975), .Z(n6977) );
  XOR U6863 ( .A(n6979), .B(n6980), .Z(n6967) );
  AND U6864 ( .A(n6981), .B(n6982), .Z(n6980) );
  XOR U6865 ( .A(n6979), .B(n6106), .Z(n6982) );
  XOR U6866 ( .A(n6983), .B(n6984), .Z(n6106) );
  AND U6867 ( .A(n270), .B(n6985), .Z(n6984) );
  XOR U6868 ( .A(n6986), .B(n6983), .Z(n6985) );
  XNOR U6869 ( .A(n6103), .B(n6979), .Z(n6981) );
  XOR U6870 ( .A(n6987), .B(n6988), .Z(n6103) );
  AND U6871 ( .A(n267), .B(n6989), .Z(n6988) );
  XOR U6872 ( .A(n6990), .B(n6987), .Z(n6989) );
  XOR U6873 ( .A(n6991), .B(n6992), .Z(n6979) );
  AND U6874 ( .A(n6993), .B(n6994), .Z(n6992) );
  XOR U6875 ( .A(n6991), .B(n6118), .Z(n6994) );
  XOR U6876 ( .A(n6995), .B(n6996), .Z(n6118) );
  AND U6877 ( .A(n270), .B(n6997), .Z(n6996) );
  XOR U6878 ( .A(n6998), .B(n6995), .Z(n6997) );
  XNOR U6879 ( .A(n6115), .B(n6991), .Z(n6993) );
  XOR U6880 ( .A(n6999), .B(n7000), .Z(n6115) );
  AND U6881 ( .A(n267), .B(n7001), .Z(n7000) );
  XOR U6882 ( .A(n7002), .B(n6999), .Z(n7001) );
  XOR U6883 ( .A(n7003), .B(n7004), .Z(n6991) );
  AND U6884 ( .A(n7005), .B(n7006), .Z(n7004) );
  XOR U6885 ( .A(n7003), .B(n6130), .Z(n7006) );
  XOR U6886 ( .A(n7007), .B(n7008), .Z(n6130) );
  AND U6887 ( .A(n270), .B(n7009), .Z(n7008) );
  XOR U6888 ( .A(n7010), .B(n7007), .Z(n7009) );
  XNOR U6889 ( .A(n6127), .B(n7003), .Z(n7005) );
  XOR U6890 ( .A(n7011), .B(n7012), .Z(n6127) );
  AND U6891 ( .A(n267), .B(n7013), .Z(n7012) );
  XOR U6892 ( .A(n7014), .B(n7011), .Z(n7013) );
  XOR U6893 ( .A(n7015), .B(n7016), .Z(n7003) );
  AND U6894 ( .A(n7017), .B(n7018), .Z(n7016) );
  XOR U6895 ( .A(n7015), .B(n6142), .Z(n7018) );
  XOR U6896 ( .A(n7019), .B(n7020), .Z(n6142) );
  AND U6897 ( .A(n270), .B(n7021), .Z(n7020) );
  XOR U6898 ( .A(n7022), .B(n7019), .Z(n7021) );
  XNOR U6899 ( .A(n6139), .B(n7015), .Z(n7017) );
  XOR U6900 ( .A(n7023), .B(n7024), .Z(n6139) );
  AND U6901 ( .A(n267), .B(n7025), .Z(n7024) );
  XOR U6902 ( .A(n7026), .B(n7023), .Z(n7025) );
  XOR U6903 ( .A(n7027), .B(n7028), .Z(n7015) );
  AND U6904 ( .A(n7029), .B(n7030), .Z(n7028) );
  XOR U6905 ( .A(n7027), .B(n6154), .Z(n7030) );
  XOR U6906 ( .A(n7031), .B(n7032), .Z(n6154) );
  AND U6907 ( .A(n270), .B(n7033), .Z(n7032) );
  XOR U6908 ( .A(n7034), .B(n7031), .Z(n7033) );
  XNOR U6909 ( .A(n6151), .B(n7027), .Z(n7029) );
  XOR U6910 ( .A(n7035), .B(n7036), .Z(n6151) );
  AND U6911 ( .A(n267), .B(n7037), .Z(n7036) );
  XOR U6912 ( .A(n7038), .B(n7035), .Z(n7037) );
  XOR U6913 ( .A(n7039), .B(n7040), .Z(n7027) );
  AND U6914 ( .A(n7041), .B(n7042), .Z(n7040) );
  XOR U6915 ( .A(n7039), .B(n6166), .Z(n7042) );
  XOR U6916 ( .A(n7043), .B(n7044), .Z(n6166) );
  AND U6917 ( .A(n270), .B(n7045), .Z(n7044) );
  XOR U6918 ( .A(n7046), .B(n7043), .Z(n7045) );
  XNOR U6919 ( .A(n6163), .B(n7039), .Z(n7041) );
  XOR U6920 ( .A(n7047), .B(n7048), .Z(n6163) );
  AND U6921 ( .A(n267), .B(n7049), .Z(n7048) );
  XOR U6922 ( .A(n7050), .B(n7047), .Z(n7049) );
  XOR U6923 ( .A(n7051), .B(n7052), .Z(n7039) );
  AND U6924 ( .A(n7053), .B(n7054), .Z(n7052) );
  XOR U6925 ( .A(n7051), .B(n6178), .Z(n7054) );
  XOR U6926 ( .A(n7055), .B(n7056), .Z(n6178) );
  AND U6927 ( .A(n270), .B(n7057), .Z(n7056) );
  XOR U6928 ( .A(n7058), .B(n7055), .Z(n7057) );
  XNOR U6929 ( .A(n6175), .B(n7051), .Z(n7053) );
  XOR U6930 ( .A(n7059), .B(n7060), .Z(n6175) );
  AND U6931 ( .A(n267), .B(n7061), .Z(n7060) );
  XOR U6932 ( .A(n7062), .B(n7059), .Z(n7061) );
  XOR U6933 ( .A(n7063), .B(n7064), .Z(n7051) );
  AND U6934 ( .A(n7065), .B(n7066), .Z(n7064) );
  XOR U6935 ( .A(n7063), .B(n6190), .Z(n7066) );
  XOR U6936 ( .A(n7067), .B(n7068), .Z(n6190) );
  AND U6937 ( .A(n270), .B(n7069), .Z(n7068) );
  XOR U6938 ( .A(n7070), .B(n7067), .Z(n7069) );
  XNOR U6939 ( .A(n6187), .B(n7063), .Z(n7065) );
  XOR U6940 ( .A(n7071), .B(n7072), .Z(n6187) );
  AND U6941 ( .A(n267), .B(n7073), .Z(n7072) );
  XOR U6942 ( .A(n7074), .B(n7071), .Z(n7073) );
  XOR U6943 ( .A(n7075), .B(n7076), .Z(n7063) );
  AND U6944 ( .A(n7077), .B(n7078), .Z(n7076) );
  XOR U6945 ( .A(n7075), .B(n6202), .Z(n7078) );
  XOR U6946 ( .A(n7079), .B(n7080), .Z(n6202) );
  AND U6947 ( .A(n270), .B(n7081), .Z(n7080) );
  XOR U6948 ( .A(n7082), .B(n7079), .Z(n7081) );
  XNOR U6949 ( .A(n6199), .B(n7075), .Z(n7077) );
  XOR U6950 ( .A(n7083), .B(n7084), .Z(n6199) );
  AND U6951 ( .A(n267), .B(n7085), .Z(n7084) );
  XOR U6952 ( .A(n7086), .B(n7083), .Z(n7085) );
  XOR U6953 ( .A(n7087), .B(n7088), .Z(n7075) );
  AND U6954 ( .A(n7089), .B(n7090), .Z(n7088) );
  XOR U6955 ( .A(n7087), .B(n6214), .Z(n7090) );
  XOR U6956 ( .A(n7091), .B(n7092), .Z(n6214) );
  AND U6957 ( .A(n270), .B(n7093), .Z(n7092) );
  XOR U6958 ( .A(n7094), .B(n7091), .Z(n7093) );
  XNOR U6959 ( .A(n6211), .B(n7087), .Z(n7089) );
  XOR U6960 ( .A(n7095), .B(n7096), .Z(n6211) );
  AND U6961 ( .A(n267), .B(n7097), .Z(n7096) );
  XOR U6962 ( .A(n7098), .B(n7095), .Z(n7097) );
  XOR U6963 ( .A(n7099), .B(n7100), .Z(n7087) );
  AND U6964 ( .A(n7101), .B(n7102), .Z(n7100) );
  XOR U6965 ( .A(n6226), .B(n7099), .Z(n7102) );
  XOR U6966 ( .A(n7103), .B(n7104), .Z(n6226) );
  AND U6967 ( .A(n270), .B(n7105), .Z(n7104) );
  XOR U6968 ( .A(n7103), .B(n7106), .Z(n7105) );
  XNOR U6969 ( .A(n7099), .B(n6223), .Z(n7101) );
  XOR U6970 ( .A(n7107), .B(n7108), .Z(n6223) );
  AND U6971 ( .A(n267), .B(n7109), .Z(n7108) );
  XOR U6972 ( .A(n7107), .B(n7110), .Z(n7109) );
  XOR U6973 ( .A(n7111), .B(n7112), .Z(n7099) );
  AND U6974 ( .A(n7113), .B(n7114), .Z(n7112) );
  XNOR U6975 ( .A(n7115), .B(n6239), .Z(n7114) );
  XOR U6976 ( .A(n7116), .B(n7117), .Z(n6239) );
  AND U6977 ( .A(n270), .B(n7118), .Z(n7117) );
  XOR U6978 ( .A(n7119), .B(n7116), .Z(n7118) );
  XNOR U6979 ( .A(n6236), .B(n7111), .Z(n7113) );
  XOR U6980 ( .A(n7120), .B(n7121), .Z(n6236) );
  AND U6981 ( .A(n267), .B(n7122), .Z(n7121) );
  XOR U6982 ( .A(n7123), .B(n7120), .Z(n7122) );
  IV U6983 ( .A(n7115), .Z(n7111) );
  AND U6984 ( .A(n6943), .B(n6946), .Z(n7115) );
  XNOR U6985 ( .A(n7124), .B(n7125), .Z(n6946) );
  AND U6986 ( .A(n270), .B(n7126), .Z(n7125) );
  XNOR U6987 ( .A(n7127), .B(n7124), .Z(n7126) );
  XOR U6988 ( .A(n7128), .B(n7129), .Z(n270) );
  AND U6989 ( .A(n7130), .B(n7131), .Z(n7129) );
  XNOR U6990 ( .A(n6951), .B(n7128), .Z(n7131) );
  AND U6991 ( .A(p_input[1151]), .B(p_input[1135]), .Z(n6951) );
  XOR U6992 ( .A(n7128), .B(n6952), .Z(n7130) );
  AND U6993 ( .A(p_input[1119]), .B(p_input[1103]), .Z(n6952) );
  XOR U6994 ( .A(n7132), .B(n7133), .Z(n7128) );
  AND U6995 ( .A(n7134), .B(n7135), .Z(n7133) );
  XOR U6996 ( .A(n7132), .B(n6962), .Z(n7135) );
  XNOR U6997 ( .A(p_input[1134]), .B(n7136), .Z(n6962) );
  AND U6998 ( .A(n202), .B(n7137), .Z(n7136) );
  XOR U6999 ( .A(p_input[1150]), .B(p_input[1134]), .Z(n7137) );
  XNOR U7000 ( .A(n6959), .B(n7132), .Z(n7134) );
  XOR U7001 ( .A(n7138), .B(n7139), .Z(n6959) );
  AND U7002 ( .A(n200), .B(n7140), .Z(n7139) );
  XOR U7003 ( .A(p_input[1118]), .B(p_input[1102]), .Z(n7140) );
  XOR U7004 ( .A(n7141), .B(n7142), .Z(n7132) );
  AND U7005 ( .A(n7143), .B(n7144), .Z(n7142) );
  XOR U7006 ( .A(n7141), .B(n6974), .Z(n7144) );
  XNOR U7007 ( .A(p_input[1133]), .B(n7145), .Z(n6974) );
  AND U7008 ( .A(n202), .B(n7146), .Z(n7145) );
  XOR U7009 ( .A(p_input[1149]), .B(p_input[1133]), .Z(n7146) );
  XNOR U7010 ( .A(n6971), .B(n7141), .Z(n7143) );
  XOR U7011 ( .A(n7147), .B(n7148), .Z(n6971) );
  AND U7012 ( .A(n200), .B(n7149), .Z(n7148) );
  XOR U7013 ( .A(p_input[1117]), .B(p_input[1101]), .Z(n7149) );
  XOR U7014 ( .A(n7150), .B(n7151), .Z(n7141) );
  AND U7015 ( .A(n7152), .B(n7153), .Z(n7151) );
  XOR U7016 ( .A(n7150), .B(n6986), .Z(n7153) );
  XNOR U7017 ( .A(p_input[1132]), .B(n7154), .Z(n6986) );
  AND U7018 ( .A(n202), .B(n7155), .Z(n7154) );
  XOR U7019 ( .A(p_input[1148]), .B(p_input[1132]), .Z(n7155) );
  XNOR U7020 ( .A(n6983), .B(n7150), .Z(n7152) );
  XOR U7021 ( .A(n7156), .B(n7157), .Z(n6983) );
  AND U7022 ( .A(n200), .B(n7158), .Z(n7157) );
  XOR U7023 ( .A(p_input[1116]), .B(p_input[1100]), .Z(n7158) );
  XOR U7024 ( .A(n7159), .B(n7160), .Z(n7150) );
  AND U7025 ( .A(n7161), .B(n7162), .Z(n7160) );
  XOR U7026 ( .A(n7159), .B(n6998), .Z(n7162) );
  XNOR U7027 ( .A(p_input[1131]), .B(n7163), .Z(n6998) );
  AND U7028 ( .A(n202), .B(n7164), .Z(n7163) );
  XOR U7029 ( .A(p_input[1147]), .B(p_input[1131]), .Z(n7164) );
  XNOR U7030 ( .A(n6995), .B(n7159), .Z(n7161) );
  XOR U7031 ( .A(n7165), .B(n7166), .Z(n6995) );
  AND U7032 ( .A(n200), .B(n7167), .Z(n7166) );
  XOR U7033 ( .A(p_input[1115]), .B(p_input[1099]), .Z(n7167) );
  XOR U7034 ( .A(n7168), .B(n7169), .Z(n7159) );
  AND U7035 ( .A(n7170), .B(n7171), .Z(n7169) );
  XOR U7036 ( .A(n7168), .B(n7010), .Z(n7171) );
  XNOR U7037 ( .A(p_input[1130]), .B(n7172), .Z(n7010) );
  AND U7038 ( .A(n202), .B(n7173), .Z(n7172) );
  XOR U7039 ( .A(p_input[1146]), .B(p_input[1130]), .Z(n7173) );
  XNOR U7040 ( .A(n7007), .B(n7168), .Z(n7170) );
  XOR U7041 ( .A(n7174), .B(n7175), .Z(n7007) );
  AND U7042 ( .A(n200), .B(n7176), .Z(n7175) );
  XOR U7043 ( .A(p_input[1114]), .B(p_input[1098]), .Z(n7176) );
  XOR U7044 ( .A(n7177), .B(n7178), .Z(n7168) );
  AND U7045 ( .A(n7179), .B(n7180), .Z(n7178) );
  XOR U7046 ( .A(n7177), .B(n7022), .Z(n7180) );
  XNOR U7047 ( .A(p_input[1129]), .B(n7181), .Z(n7022) );
  AND U7048 ( .A(n202), .B(n7182), .Z(n7181) );
  XOR U7049 ( .A(p_input[1145]), .B(p_input[1129]), .Z(n7182) );
  XNOR U7050 ( .A(n7019), .B(n7177), .Z(n7179) );
  XOR U7051 ( .A(n7183), .B(n7184), .Z(n7019) );
  AND U7052 ( .A(n200), .B(n7185), .Z(n7184) );
  XOR U7053 ( .A(p_input[1113]), .B(p_input[1097]), .Z(n7185) );
  XOR U7054 ( .A(n7186), .B(n7187), .Z(n7177) );
  AND U7055 ( .A(n7188), .B(n7189), .Z(n7187) );
  XOR U7056 ( .A(n7186), .B(n7034), .Z(n7189) );
  XNOR U7057 ( .A(p_input[1128]), .B(n7190), .Z(n7034) );
  AND U7058 ( .A(n202), .B(n7191), .Z(n7190) );
  XOR U7059 ( .A(p_input[1144]), .B(p_input[1128]), .Z(n7191) );
  XNOR U7060 ( .A(n7031), .B(n7186), .Z(n7188) );
  XOR U7061 ( .A(n7192), .B(n7193), .Z(n7031) );
  AND U7062 ( .A(n200), .B(n7194), .Z(n7193) );
  XOR U7063 ( .A(p_input[1112]), .B(p_input[1096]), .Z(n7194) );
  XOR U7064 ( .A(n7195), .B(n7196), .Z(n7186) );
  AND U7065 ( .A(n7197), .B(n7198), .Z(n7196) );
  XOR U7066 ( .A(n7195), .B(n7046), .Z(n7198) );
  XNOR U7067 ( .A(p_input[1127]), .B(n7199), .Z(n7046) );
  AND U7068 ( .A(n202), .B(n7200), .Z(n7199) );
  XOR U7069 ( .A(p_input[1143]), .B(p_input[1127]), .Z(n7200) );
  XNOR U7070 ( .A(n7043), .B(n7195), .Z(n7197) );
  XOR U7071 ( .A(n7201), .B(n7202), .Z(n7043) );
  AND U7072 ( .A(n200), .B(n7203), .Z(n7202) );
  XOR U7073 ( .A(p_input[1111]), .B(p_input[1095]), .Z(n7203) );
  XOR U7074 ( .A(n7204), .B(n7205), .Z(n7195) );
  AND U7075 ( .A(n7206), .B(n7207), .Z(n7205) );
  XOR U7076 ( .A(n7204), .B(n7058), .Z(n7207) );
  XNOR U7077 ( .A(p_input[1126]), .B(n7208), .Z(n7058) );
  AND U7078 ( .A(n202), .B(n7209), .Z(n7208) );
  XOR U7079 ( .A(p_input[1142]), .B(p_input[1126]), .Z(n7209) );
  XNOR U7080 ( .A(n7055), .B(n7204), .Z(n7206) );
  XOR U7081 ( .A(n7210), .B(n7211), .Z(n7055) );
  AND U7082 ( .A(n200), .B(n7212), .Z(n7211) );
  XOR U7083 ( .A(p_input[1110]), .B(p_input[1094]), .Z(n7212) );
  XOR U7084 ( .A(n7213), .B(n7214), .Z(n7204) );
  AND U7085 ( .A(n7215), .B(n7216), .Z(n7214) );
  XOR U7086 ( .A(n7213), .B(n7070), .Z(n7216) );
  XNOR U7087 ( .A(p_input[1125]), .B(n7217), .Z(n7070) );
  AND U7088 ( .A(n202), .B(n7218), .Z(n7217) );
  XOR U7089 ( .A(p_input[1141]), .B(p_input[1125]), .Z(n7218) );
  XNOR U7090 ( .A(n7067), .B(n7213), .Z(n7215) );
  XOR U7091 ( .A(n7219), .B(n7220), .Z(n7067) );
  AND U7092 ( .A(n200), .B(n7221), .Z(n7220) );
  XOR U7093 ( .A(p_input[1109]), .B(p_input[1093]), .Z(n7221) );
  XOR U7094 ( .A(n7222), .B(n7223), .Z(n7213) );
  AND U7095 ( .A(n7224), .B(n7225), .Z(n7223) );
  XOR U7096 ( .A(n7222), .B(n7082), .Z(n7225) );
  XNOR U7097 ( .A(p_input[1124]), .B(n7226), .Z(n7082) );
  AND U7098 ( .A(n202), .B(n7227), .Z(n7226) );
  XOR U7099 ( .A(p_input[1140]), .B(p_input[1124]), .Z(n7227) );
  XNOR U7100 ( .A(n7079), .B(n7222), .Z(n7224) );
  XOR U7101 ( .A(n7228), .B(n7229), .Z(n7079) );
  AND U7102 ( .A(n200), .B(n7230), .Z(n7229) );
  XOR U7103 ( .A(p_input[1108]), .B(p_input[1092]), .Z(n7230) );
  XOR U7104 ( .A(n7231), .B(n7232), .Z(n7222) );
  AND U7105 ( .A(n7233), .B(n7234), .Z(n7232) );
  XOR U7106 ( .A(n7231), .B(n7094), .Z(n7234) );
  XNOR U7107 ( .A(p_input[1123]), .B(n7235), .Z(n7094) );
  AND U7108 ( .A(n202), .B(n7236), .Z(n7235) );
  XOR U7109 ( .A(p_input[1139]), .B(p_input[1123]), .Z(n7236) );
  XNOR U7110 ( .A(n7091), .B(n7231), .Z(n7233) );
  XOR U7111 ( .A(n7237), .B(n7238), .Z(n7091) );
  AND U7112 ( .A(n200), .B(n7239), .Z(n7238) );
  XOR U7113 ( .A(p_input[1107]), .B(p_input[1091]), .Z(n7239) );
  XOR U7114 ( .A(n7240), .B(n7241), .Z(n7231) );
  AND U7115 ( .A(n7242), .B(n7243), .Z(n7241) );
  XOR U7116 ( .A(n7106), .B(n7240), .Z(n7243) );
  XNOR U7117 ( .A(p_input[1122]), .B(n7244), .Z(n7106) );
  AND U7118 ( .A(n202), .B(n7245), .Z(n7244) );
  XOR U7119 ( .A(p_input[1138]), .B(p_input[1122]), .Z(n7245) );
  XNOR U7120 ( .A(n7240), .B(n7103), .Z(n7242) );
  XOR U7121 ( .A(n7246), .B(n7247), .Z(n7103) );
  AND U7122 ( .A(n200), .B(n7248), .Z(n7247) );
  XOR U7123 ( .A(p_input[1106]), .B(p_input[1090]), .Z(n7248) );
  XOR U7124 ( .A(n7249), .B(n7250), .Z(n7240) );
  AND U7125 ( .A(n7251), .B(n7252), .Z(n7250) );
  XNOR U7126 ( .A(n7253), .B(n7119), .Z(n7252) );
  XNOR U7127 ( .A(p_input[1121]), .B(n7254), .Z(n7119) );
  AND U7128 ( .A(n202), .B(n7255), .Z(n7254) );
  XNOR U7129 ( .A(p_input[1137]), .B(n7256), .Z(n7255) );
  IV U7130 ( .A(p_input[1121]), .Z(n7256) );
  XNOR U7131 ( .A(n7116), .B(n7249), .Z(n7251) );
  XNOR U7132 ( .A(p_input[1089]), .B(n7257), .Z(n7116) );
  AND U7133 ( .A(n200), .B(n7258), .Z(n7257) );
  XOR U7134 ( .A(p_input[1105]), .B(p_input[1089]), .Z(n7258) );
  IV U7135 ( .A(n7253), .Z(n7249) );
  AND U7136 ( .A(n7124), .B(n7127), .Z(n7253) );
  XOR U7137 ( .A(p_input[1120]), .B(n7259), .Z(n7127) );
  AND U7138 ( .A(n202), .B(n7260), .Z(n7259) );
  XOR U7139 ( .A(p_input[1136]), .B(p_input[1120]), .Z(n7260) );
  XOR U7140 ( .A(n7261), .B(n7262), .Z(n202) );
  AND U7141 ( .A(n7263), .B(n7264), .Z(n7262) );
  XNOR U7142 ( .A(p_input[1151]), .B(n7261), .Z(n7264) );
  XOR U7143 ( .A(n7261), .B(p_input[1135]), .Z(n7263) );
  XOR U7144 ( .A(n7265), .B(n7266), .Z(n7261) );
  AND U7145 ( .A(n7267), .B(n7268), .Z(n7266) );
  XNOR U7146 ( .A(p_input[1150]), .B(n7265), .Z(n7268) );
  XOR U7147 ( .A(n7265), .B(p_input[1134]), .Z(n7267) );
  XOR U7148 ( .A(n7269), .B(n7270), .Z(n7265) );
  AND U7149 ( .A(n7271), .B(n7272), .Z(n7270) );
  XNOR U7150 ( .A(p_input[1149]), .B(n7269), .Z(n7272) );
  XOR U7151 ( .A(n7269), .B(p_input[1133]), .Z(n7271) );
  XOR U7152 ( .A(n7273), .B(n7274), .Z(n7269) );
  AND U7153 ( .A(n7275), .B(n7276), .Z(n7274) );
  XNOR U7154 ( .A(p_input[1148]), .B(n7273), .Z(n7276) );
  XOR U7155 ( .A(n7273), .B(p_input[1132]), .Z(n7275) );
  XOR U7156 ( .A(n7277), .B(n7278), .Z(n7273) );
  AND U7157 ( .A(n7279), .B(n7280), .Z(n7278) );
  XNOR U7158 ( .A(p_input[1147]), .B(n7277), .Z(n7280) );
  XOR U7159 ( .A(n7277), .B(p_input[1131]), .Z(n7279) );
  XOR U7160 ( .A(n7281), .B(n7282), .Z(n7277) );
  AND U7161 ( .A(n7283), .B(n7284), .Z(n7282) );
  XNOR U7162 ( .A(p_input[1146]), .B(n7281), .Z(n7284) );
  XOR U7163 ( .A(n7281), .B(p_input[1130]), .Z(n7283) );
  XOR U7164 ( .A(n7285), .B(n7286), .Z(n7281) );
  AND U7165 ( .A(n7287), .B(n7288), .Z(n7286) );
  XNOR U7166 ( .A(p_input[1145]), .B(n7285), .Z(n7288) );
  XOR U7167 ( .A(n7285), .B(p_input[1129]), .Z(n7287) );
  XOR U7168 ( .A(n7289), .B(n7290), .Z(n7285) );
  AND U7169 ( .A(n7291), .B(n7292), .Z(n7290) );
  XNOR U7170 ( .A(p_input[1144]), .B(n7289), .Z(n7292) );
  XOR U7171 ( .A(n7289), .B(p_input[1128]), .Z(n7291) );
  XOR U7172 ( .A(n7293), .B(n7294), .Z(n7289) );
  AND U7173 ( .A(n7295), .B(n7296), .Z(n7294) );
  XNOR U7174 ( .A(p_input[1143]), .B(n7293), .Z(n7296) );
  XOR U7175 ( .A(n7293), .B(p_input[1127]), .Z(n7295) );
  XOR U7176 ( .A(n7297), .B(n7298), .Z(n7293) );
  AND U7177 ( .A(n7299), .B(n7300), .Z(n7298) );
  XNOR U7178 ( .A(p_input[1142]), .B(n7297), .Z(n7300) );
  XOR U7179 ( .A(n7297), .B(p_input[1126]), .Z(n7299) );
  XOR U7180 ( .A(n7301), .B(n7302), .Z(n7297) );
  AND U7181 ( .A(n7303), .B(n7304), .Z(n7302) );
  XNOR U7182 ( .A(p_input[1141]), .B(n7301), .Z(n7304) );
  XOR U7183 ( .A(n7301), .B(p_input[1125]), .Z(n7303) );
  XOR U7184 ( .A(n7305), .B(n7306), .Z(n7301) );
  AND U7185 ( .A(n7307), .B(n7308), .Z(n7306) );
  XNOR U7186 ( .A(p_input[1140]), .B(n7305), .Z(n7308) );
  XOR U7187 ( .A(n7305), .B(p_input[1124]), .Z(n7307) );
  XOR U7188 ( .A(n7309), .B(n7310), .Z(n7305) );
  AND U7189 ( .A(n7311), .B(n7312), .Z(n7310) );
  XNOR U7190 ( .A(p_input[1139]), .B(n7309), .Z(n7312) );
  XOR U7191 ( .A(n7309), .B(p_input[1123]), .Z(n7311) );
  XOR U7192 ( .A(n7313), .B(n7314), .Z(n7309) );
  AND U7193 ( .A(n7315), .B(n7316), .Z(n7314) );
  XNOR U7194 ( .A(p_input[1138]), .B(n7313), .Z(n7316) );
  XOR U7195 ( .A(n7313), .B(p_input[1122]), .Z(n7315) );
  XNOR U7196 ( .A(n7317), .B(n7318), .Z(n7313) );
  AND U7197 ( .A(n7319), .B(n7320), .Z(n7318) );
  XOR U7198 ( .A(p_input[1137]), .B(n7317), .Z(n7320) );
  XNOR U7199 ( .A(p_input[1121]), .B(n7317), .Z(n7319) );
  AND U7200 ( .A(p_input[1136]), .B(n7321), .Z(n7317) );
  IV U7201 ( .A(p_input[1120]), .Z(n7321) );
  XNOR U7202 ( .A(p_input[1088]), .B(n7322), .Z(n7124) );
  AND U7203 ( .A(n200), .B(n7323), .Z(n7322) );
  XOR U7204 ( .A(p_input[1104]), .B(p_input[1088]), .Z(n7323) );
  XOR U7205 ( .A(n7324), .B(n7325), .Z(n200) );
  AND U7206 ( .A(n7326), .B(n7327), .Z(n7325) );
  XNOR U7207 ( .A(p_input[1119]), .B(n7324), .Z(n7327) );
  XOR U7208 ( .A(n7324), .B(p_input[1103]), .Z(n7326) );
  XOR U7209 ( .A(n7328), .B(n7329), .Z(n7324) );
  AND U7210 ( .A(n7330), .B(n7331), .Z(n7329) );
  XNOR U7211 ( .A(p_input[1118]), .B(n7328), .Z(n7331) );
  XNOR U7212 ( .A(n7328), .B(n7138), .Z(n7330) );
  IV U7213 ( .A(p_input[1102]), .Z(n7138) );
  XOR U7214 ( .A(n7332), .B(n7333), .Z(n7328) );
  AND U7215 ( .A(n7334), .B(n7335), .Z(n7333) );
  XNOR U7216 ( .A(p_input[1117]), .B(n7332), .Z(n7335) );
  XNOR U7217 ( .A(n7332), .B(n7147), .Z(n7334) );
  IV U7218 ( .A(p_input[1101]), .Z(n7147) );
  XOR U7219 ( .A(n7336), .B(n7337), .Z(n7332) );
  AND U7220 ( .A(n7338), .B(n7339), .Z(n7337) );
  XNOR U7221 ( .A(p_input[1116]), .B(n7336), .Z(n7339) );
  XNOR U7222 ( .A(n7336), .B(n7156), .Z(n7338) );
  IV U7223 ( .A(p_input[1100]), .Z(n7156) );
  XOR U7224 ( .A(n7340), .B(n7341), .Z(n7336) );
  AND U7225 ( .A(n7342), .B(n7343), .Z(n7341) );
  XNOR U7226 ( .A(p_input[1115]), .B(n7340), .Z(n7343) );
  XNOR U7227 ( .A(n7340), .B(n7165), .Z(n7342) );
  IV U7228 ( .A(p_input[1099]), .Z(n7165) );
  XOR U7229 ( .A(n7344), .B(n7345), .Z(n7340) );
  AND U7230 ( .A(n7346), .B(n7347), .Z(n7345) );
  XNOR U7231 ( .A(p_input[1114]), .B(n7344), .Z(n7347) );
  XNOR U7232 ( .A(n7344), .B(n7174), .Z(n7346) );
  IV U7233 ( .A(p_input[1098]), .Z(n7174) );
  XOR U7234 ( .A(n7348), .B(n7349), .Z(n7344) );
  AND U7235 ( .A(n7350), .B(n7351), .Z(n7349) );
  XNOR U7236 ( .A(p_input[1113]), .B(n7348), .Z(n7351) );
  XNOR U7237 ( .A(n7348), .B(n7183), .Z(n7350) );
  IV U7238 ( .A(p_input[1097]), .Z(n7183) );
  XOR U7239 ( .A(n7352), .B(n7353), .Z(n7348) );
  AND U7240 ( .A(n7354), .B(n7355), .Z(n7353) );
  XNOR U7241 ( .A(p_input[1112]), .B(n7352), .Z(n7355) );
  XNOR U7242 ( .A(n7352), .B(n7192), .Z(n7354) );
  IV U7243 ( .A(p_input[1096]), .Z(n7192) );
  XOR U7244 ( .A(n7356), .B(n7357), .Z(n7352) );
  AND U7245 ( .A(n7358), .B(n7359), .Z(n7357) );
  XNOR U7246 ( .A(p_input[1111]), .B(n7356), .Z(n7359) );
  XNOR U7247 ( .A(n7356), .B(n7201), .Z(n7358) );
  IV U7248 ( .A(p_input[1095]), .Z(n7201) );
  XOR U7249 ( .A(n7360), .B(n7361), .Z(n7356) );
  AND U7250 ( .A(n7362), .B(n7363), .Z(n7361) );
  XNOR U7251 ( .A(p_input[1110]), .B(n7360), .Z(n7363) );
  XNOR U7252 ( .A(n7360), .B(n7210), .Z(n7362) );
  IV U7253 ( .A(p_input[1094]), .Z(n7210) );
  XOR U7254 ( .A(n7364), .B(n7365), .Z(n7360) );
  AND U7255 ( .A(n7366), .B(n7367), .Z(n7365) );
  XNOR U7256 ( .A(p_input[1109]), .B(n7364), .Z(n7367) );
  XNOR U7257 ( .A(n7364), .B(n7219), .Z(n7366) );
  IV U7258 ( .A(p_input[1093]), .Z(n7219) );
  XOR U7259 ( .A(n7368), .B(n7369), .Z(n7364) );
  AND U7260 ( .A(n7370), .B(n7371), .Z(n7369) );
  XNOR U7261 ( .A(p_input[1108]), .B(n7368), .Z(n7371) );
  XNOR U7262 ( .A(n7368), .B(n7228), .Z(n7370) );
  IV U7263 ( .A(p_input[1092]), .Z(n7228) );
  XOR U7264 ( .A(n7372), .B(n7373), .Z(n7368) );
  AND U7265 ( .A(n7374), .B(n7375), .Z(n7373) );
  XNOR U7266 ( .A(p_input[1107]), .B(n7372), .Z(n7375) );
  XNOR U7267 ( .A(n7372), .B(n7237), .Z(n7374) );
  IV U7268 ( .A(p_input[1091]), .Z(n7237) );
  XOR U7269 ( .A(n7376), .B(n7377), .Z(n7372) );
  AND U7270 ( .A(n7378), .B(n7379), .Z(n7377) );
  XNOR U7271 ( .A(p_input[1106]), .B(n7376), .Z(n7379) );
  XNOR U7272 ( .A(n7376), .B(n7246), .Z(n7378) );
  IV U7273 ( .A(p_input[1090]), .Z(n7246) );
  XNOR U7274 ( .A(n7380), .B(n7381), .Z(n7376) );
  AND U7275 ( .A(n7382), .B(n7383), .Z(n7381) );
  XOR U7276 ( .A(p_input[1105]), .B(n7380), .Z(n7383) );
  XNOR U7277 ( .A(p_input[1089]), .B(n7380), .Z(n7382) );
  AND U7278 ( .A(p_input[1104]), .B(n7384), .Z(n7380) );
  IV U7279 ( .A(p_input[1088]), .Z(n7384) );
  XOR U7280 ( .A(n7385), .B(n7386), .Z(n6943) );
  AND U7281 ( .A(n267), .B(n7387), .Z(n7386) );
  XNOR U7282 ( .A(n7388), .B(n7385), .Z(n7387) );
  XOR U7283 ( .A(n7389), .B(n7390), .Z(n267) );
  AND U7284 ( .A(n7391), .B(n7392), .Z(n7390) );
  XNOR U7285 ( .A(n6954), .B(n7389), .Z(n7392) );
  AND U7286 ( .A(p_input[1087]), .B(p_input[1071]), .Z(n6954) );
  XOR U7287 ( .A(n7389), .B(n6953), .Z(n7391) );
  AND U7288 ( .A(p_input[1039]), .B(p_input[1055]), .Z(n6953) );
  XOR U7289 ( .A(n7393), .B(n7394), .Z(n7389) );
  AND U7290 ( .A(n7395), .B(n7396), .Z(n7394) );
  XOR U7291 ( .A(n7393), .B(n6966), .Z(n7396) );
  XNOR U7292 ( .A(p_input[1070]), .B(n7397), .Z(n6966) );
  AND U7293 ( .A(n206), .B(n7398), .Z(n7397) );
  XOR U7294 ( .A(p_input[1086]), .B(p_input[1070]), .Z(n7398) );
  XNOR U7295 ( .A(n6963), .B(n7393), .Z(n7395) );
  XOR U7296 ( .A(n7399), .B(n7400), .Z(n6963) );
  AND U7297 ( .A(n203), .B(n7401), .Z(n7400) );
  XOR U7298 ( .A(p_input[1054]), .B(p_input[1038]), .Z(n7401) );
  XOR U7299 ( .A(n7402), .B(n7403), .Z(n7393) );
  AND U7300 ( .A(n7404), .B(n7405), .Z(n7403) );
  XOR U7301 ( .A(n7402), .B(n6978), .Z(n7405) );
  XNOR U7302 ( .A(p_input[1069]), .B(n7406), .Z(n6978) );
  AND U7303 ( .A(n206), .B(n7407), .Z(n7406) );
  XOR U7304 ( .A(p_input[1085]), .B(p_input[1069]), .Z(n7407) );
  XNOR U7305 ( .A(n6975), .B(n7402), .Z(n7404) );
  XOR U7306 ( .A(n7408), .B(n7409), .Z(n6975) );
  AND U7307 ( .A(n203), .B(n7410), .Z(n7409) );
  XOR U7308 ( .A(p_input[1053]), .B(p_input[1037]), .Z(n7410) );
  XOR U7309 ( .A(n7411), .B(n7412), .Z(n7402) );
  AND U7310 ( .A(n7413), .B(n7414), .Z(n7412) );
  XOR U7311 ( .A(n7411), .B(n6990), .Z(n7414) );
  XNOR U7312 ( .A(p_input[1068]), .B(n7415), .Z(n6990) );
  AND U7313 ( .A(n206), .B(n7416), .Z(n7415) );
  XOR U7314 ( .A(p_input[1084]), .B(p_input[1068]), .Z(n7416) );
  XNOR U7315 ( .A(n6987), .B(n7411), .Z(n7413) );
  XOR U7316 ( .A(n7417), .B(n7418), .Z(n6987) );
  AND U7317 ( .A(n203), .B(n7419), .Z(n7418) );
  XOR U7318 ( .A(p_input[1052]), .B(p_input[1036]), .Z(n7419) );
  XOR U7319 ( .A(n7420), .B(n7421), .Z(n7411) );
  AND U7320 ( .A(n7422), .B(n7423), .Z(n7421) );
  XOR U7321 ( .A(n7420), .B(n7002), .Z(n7423) );
  XNOR U7322 ( .A(p_input[1067]), .B(n7424), .Z(n7002) );
  AND U7323 ( .A(n206), .B(n7425), .Z(n7424) );
  XOR U7324 ( .A(p_input[1083]), .B(p_input[1067]), .Z(n7425) );
  XNOR U7325 ( .A(n6999), .B(n7420), .Z(n7422) );
  XOR U7326 ( .A(n7426), .B(n7427), .Z(n6999) );
  AND U7327 ( .A(n203), .B(n7428), .Z(n7427) );
  XOR U7328 ( .A(p_input[1051]), .B(p_input[1035]), .Z(n7428) );
  XOR U7329 ( .A(n7429), .B(n7430), .Z(n7420) );
  AND U7330 ( .A(n7431), .B(n7432), .Z(n7430) );
  XOR U7331 ( .A(n7429), .B(n7014), .Z(n7432) );
  XNOR U7332 ( .A(p_input[1066]), .B(n7433), .Z(n7014) );
  AND U7333 ( .A(n206), .B(n7434), .Z(n7433) );
  XOR U7334 ( .A(p_input[1082]), .B(p_input[1066]), .Z(n7434) );
  XNOR U7335 ( .A(n7011), .B(n7429), .Z(n7431) );
  XOR U7336 ( .A(n7435), .B(n7436), .Z(n7011) );
  AND U7337 ( .A(n203), .B(n7437), .Z(n7436) );
  XOR U7338 ( .A(p_input[1050]), .B(p_input[1034]), .Z(n7437) );
  XOR U7339 ( .A(n7438), .B(n7439), .Z(n7429) );
  AND U7340 ( .A(n7440), .B(n7441), .Z(n7439) );
  XOR U7341 ( .A(n7438), .B(n7026), .Z(n7441) );
  XNOR U7342 ( .A(p_input[1065]), .B(n7442), .Z(n7026) );
  AND U7343 ( .A(n206), .B(n7443), .Z(n7442) );
  XOR U7344 ( .A(p_input[1081]), .B(p_input[1065]), .Z(n7443) );
  XNOR U7345 ( .A(n7023), .B(n7438), .Z(n7440) );
  XOR U7346 ( .A(n7444), .B(n7445), .Z(n7023) );
  AND U7347 ( .A(n203), .B(n7446), .Z(n7445) );
  XOR U7348 ( .A(p_input[1049]), .B(p_input[1033]), .Z(n7446) );
  XOR U7349 ( .A(n7447), .B(n7448), .Z(n7438) );
  AND U7350 ( .A(n7449), .B(n7450), .Z(n7448) );
  XOR U7351 ( .A(n7447), .B(n7038), .Z(n7450) );
  XNOR U7352 ( .A(p_input[1064]), .B(n7451), .Z(n7038) );
  AND U7353 ( .A(n206), .B(n7452), .Z(n7451) );
  XOR U7354 ( .A(p_input[1080]), .B(p_input[1064]), .Z(n7452) );
  XNOR U7355 ( .A(n7035), .B(n7447), .Z(n7449) );
  XOR U7356 ( .A(n7453), .B(n7454), .Z(n7035) );
  AND U7357 ( .A(n203), .B(n7455), .Z(n7454) );
  XOR U7358 ( .A(p_input[1048]), .B(p_input[1032]), .Z(n7455) );
  XOR U7359 ( .A(n7456), .B(n7457), .Z(n7447) );
  AND U7360 ( .A(n7458), .B(n7459), .Z(n7457) );
  XOR U7361 ( .A(n7456), .B(n7050), .Z(n7459) );
  XNOR U7362 ( .A(p_input[1063]), .B(n7460), .Z(n7050) );
  AND U7363 ( .A(n206), .B(n7461), .Z(n7460) );
  XOR U7364 ( .A(p_input[1079]), .B(p_input[1063]), .Z(n7461) );
  XNOR U7365 ( .A(n7047), .B(n7456), .Z(n7458) );
  XOR U7366 ( .A(n7462), .B(n7463), .Z(n7047) );
  AND U7367 ( .A(n203), .B(n7464), .Z(n7463) );
  XOR U7368 ( .A(p_input[1047]), .B(p_input[1031]), .Z(n7464) );
  XOR U7369 ( .A(n7465), .B(n7466), .Z(n7456) );
  AND U7370 ( .A(n7467), .B(n7468), .Z(n7466) );
  XOR U7371 ( .A(n7465), .B(n7062), .Z(n7468) );
  XNOR U7372 ( .A(p_input[1062]), .B(n7469), .Z(n7062) );
  AND U7373 ( .A(n206), .B(n7470), .Z(n7469) );
  XOR U7374 ( .A(p_input[1078]), .B(p_input[1062]), .Z(n7470) );
  XNOR U7375 ( .A(n7059), .B(n7465), .Z(n7467) );
  XOR U7376 ( .A(n7471), .B(n7472), .Z(n7059) );
  AND U7377 ( .A(n203), .B(n7473), .Z(n7472) );
  XOR U7378 ( .A(p_input[1046]), .B(p_input[1030]), .Z(n7473) );
  XOR U7379 ( .A(n7474), .B(n7475), .Z(n7465) );
  AND U7380 ( .A(n7476), .B(n7477), .Z(n7475) );
  XOR U7381 ( .A(n7474), .B(n7074), .Z(n7477) );
  XNOR U7382 ( .A(p_input[1061]), .B(n7478), .Z(n7074) );
  AND U7383 ( .A(n206), .B(n7479), .Z(n7478) );
  XOR U7384 ( .A(p_input[1077]), .B(p_input[1061]), .Z(n7479) );
  XNOR U7385 ( .A(n7071), .B(n7474), .Z(n7476) );
  XOR U7386 ( .A(n7480), .B(n7481), .Z(n7071) );
  AND U7387 ( .A(n203), .B(n7482), .Z(n7481) );
  XOR U7388 ( .A(p_input[1045]), .B(p_input[1029]), .Z(n7482) );
  XOR U7389 ( .A(n7483), .B(n7484), .Z(n7474) );
  AND U7390 ( .A(n7485), .B(n7486), .Z(n7484) );
  XOR U7391 ( .A(n7483), .B(n7086), .Z(n7486) );
  XNOR U7392 ( .A(p_input[1060]), .B(n7487), .Z(n7086) );
  AND U7393 ( .A(n206), .B(n7488), .Z(n7487) );
  XOR U7394 ( .A(p_input[1076]), .B(p_input[1060]), .Z(n7488) );
  XNOR U7395 ( .A(n7083), .B(n7483), .Z(n7485) );
  XOR U7396 ( .A(n7489), .B(n7490), .Z(n7083) );
  AND U7397 ( .A(n203), .B(n7491), .Z(n7490) );
  XOR U7398 ( .A(p_input[1044]), .B(p_input[1028]), .Z(n7491) );
  XOR U7399 ( .A(n7492), .B(n7493), .Z(n7483) );
  AND U7400 ( .A(n7494), .B(n7495), .Z(n7493) );
  XOR U7401 ( .A(n7492), .B(n7098), .Z(n7495) );
  XNOR U7402 ( .A(p_input[1059]), .B(n7496), .Z(n7098) );
  AND U7403 ( .A(n206), .B(n7497), .Z(n7496) );
  XOR U7404 ( .A(p_input[1075]), .B(p_input[1059]), .Z(n7497) );
  XNOR U7405 ( .A(n7095), .B(n7492), .Z(n7494) );
  XOR U7406 ( .A(n7498), .B(n7499), .Z(n7095) );
  AND U7407 ( .A(n203), .B(n7500), .Z(n7499) );
  XOR U7408 ( .A(p_input[1043]), .B(p_input[1027]), .Z(n7500) );
  XOR U7409 ( .A(n7501), .B(n7502), .Z(n7492) );
  AND U7410 ( .A(n7503), .B(n7504), .Z(n7502) );
  XOR U7411 ( .A(n7110), .B(n7501), .Z(n7504) );
  XNOR U7412 ( .A(p_input[1058]), .B(n7505), .Z(n7110) );
  AND U7413 ( .A(n206), .B(n7506), .Z(n7505) );
  XOR U7414 ( .A(p_input[1074]), .B(p_input[1058]), .Z(n7506) );
  XNOR U7415 ( .A(n7501), .B(n7107), .Z(n7503) );
  XOR U7416 ( .A(n7507), .B(n7508), .Z(n7107) );
  AND U7417 ( .A(n203), .B(n7509), .Z(n7508) );
  XOR U7418 ( .A(p_input[1042]), .B(p_input[1026]), .Z(n7509) );
  XOR U7419 ( .A(n7510), .B(n7511), .Z(n7501) );
  AND U7420 ( .A(n7512), .B(n7513), .Z(n7511) );
  XNOR U7421 ( .A(n7514), .B(n7123), .Z(n7513) );
  XNOR U7422 ( .A(p_input[1057]), .B(n7515), .Z(n7123) );
  AND U7423 ( .A(n206), .B(n7516), .Z(n7515) );
  XNOR U7424 ( .A(p_input[1073]), .B(n7517), .Z(n7516) );
  IV U7425 ( .A(p_input[1057]), .Z(n7517) );
  XNOR U7426 ( .A(n7120), .B(n7510), .Z(n7512) );
  XNOR U7427 ( .A(p_input[1025]), .B(n7518), .Z(n7120) );
  AND U7428 ( .A(n203), .B(n7519), .Z(n7518) );
  XOR U7429 ( .A(p_input[1041]), .B(p_input[1025]), .Z(n7519) );
  IV U7430 ( .A(n7514), .Z(n7510) );
  AND U7431 ( .A(n7385), .B(n7388), .Z(n7514) );
  XOR U7432 ( .A(p_input[1056]), .B(n7520), .Z(n7388) );
  AND U7433 ( .A(n206), .B(n7521), .Z(n7520) );
  XOR U7434 ( .A(p_input[1072]), .B(p_input[1056]), .Z(n7521) );
  XOR U7435 ( .A(n7522), .B(n7523), .Z(n206) );
  AND U7436 ( .A(n7524), .B(n7525), .Z(n7523) );
  XNOR U7437 ( .A(p_input[1087]), .B(n7522), .Z(n7525) );
  XOR U7438 ( .A(n7522), .B(p_input[1071]), .Z(n7524) );
  XOR U7439 ( .A(n7526), .B(n7527), .Z(n7522) );
  AND U7440 ( .A(n7528), .B(n7529), .Z(n7527) );
  XNOR U7441 ( .A(p_input[1086]), .B(n7526), .Z(n7529) );
  XOR U7442 ( .A(n7526), .B(p_input[1070]), .Z(n7528) );
  XOR U7443 ( .A(n7530), .B(n7531), .Z(n7526) );
  AND U7444 ( .A(n7532), .B(n7533), .Z(n7531) );
  XNOR U7445 ( .A(p_input[1085]), .B(n7530), .Z(n7533) );
  XOR U7446 ( .A(n7530), .B(p_input[1069]), .Z(n7532) );
  XOR U7447 ( .A(n7534), .B(n7535), .Z(n7530) );
  AND U7448 ( .A(n7536), .B(n7537), .Z(n7535) );
  XNOR U7449 ( .A(p_input[1084]), .B(n7534), .Z(n7537) );
  XOR U7450 ( .A(n7534), .B(p_input[1068]), .Z(n7536) );
  XOR U7451 ( .A(n7538), .B(n7539), .Z(n7534) );
  AND U7452 ( .A(n7540), .B(n7541), .Z(n7539) );
  XNOR U7453 ( .A(p_input[1083]), .B(n7538), .Z(n7541) );
  XOR U7454 ( .A(n7538), .B(p_input[1067]), .Z(n7540) );
  XOR U7455 ( .A(n7542), .B(n7543), .Z(n7538) );
  AND U7456 ( .A(n7544), .B(n7545), .Z(n7543) );
  XNOR U7457 ( .A(p_input[1082]), .B(n7542), .Z(n7545) );
  XOR U7458 ( .A(n7542), .B(p_input[1066]), .Z(n7544) );
  XOR U7459 ( .A(n7546), .B(n7547), .Z(n7542) );
  AND U7460 ( .A(n7548), .B(n7549), .Z(n7547) );
  XNOR U7461 ( .A(p_input[1081]), .B(n7546), .Z(n7549) );
  XOR U7462 ( .A(n7546), .B(p_input[1065]), .Z(n7548) );
  XOR U7463 ( .A(n7550), .B(n7551), .Z(n7546) );
  AND U7464 ( .A(n7552), .B(n7553), .Z(n7551) );
  XNOR U7465 ( .A(p_input[1080]), .B(n7550), .Z(n7553) );
  XOR U7466 ( .A(n7550), .B(p_input[1064]), .Z(n7552) );
  XOR U7467 ( .A(n7554), .B(n7555), .Z(n7550) );
  AND U7468 ( .A(n7556), .B(n7557), .Z(n7555) );
  XNOR U7469 ( .A(p_input[1079]), .B(n7554), .Z(n7557) );
  XOR U7470 ( .A(n7554), .B(p_input[1063]), .Z(n7556) );
  XOR U7471 ( .A(n7558), .B(n7559), .Z(n7554) );
  AND U7472 ( .A(n7560), .B(n7561), .Z(n7559) );
  XNOR U7473 ( .A(p_input[1078]), .B(n7558), .Z(n7561) );
  XOR U7474 ( .A(n7558), .B(p_input[1062]), .Z(n7560) );
  XOR U7475 ( .A(n7562), .B(n7563), .Z(n7558) );
  AND U7476 ( .A(n7564), .B(n7565), .Z(n7563) );
  XNOR U7477 ( .A(p_input[1077]), .B(n7562), .Z(n7565) );
  XOR U7478 ( .A(n7562), .B(p_input[1061]), .Z(n7564) );
  XOR U7479 ( .A(n7566), .B(n7567), .Z(n7562) );
  AND U7480 ( .A(n7568), .B(n7569), .Z(n7567) );
  XNOR U7481 ( .A(p_input[1076]), .B(n7566), .Z(n7569) );
  XOR U7482 ( .A(n7566), .B(p_input[1060]), .Z(n7568) );
  XOR U7483 ( .A(n7570), .B(n7571), .Z(n7566) );
  AND U7484 ( .A(n7572), .B(n7573), .Z(n7571) );
  XNOR U7485 ( .A(p_input[1075]), .B(n7570), .Z(n7573) );
  XOR U7486 ( .A(n7570), .B(p_input[1059]), .Z(n7572) );
  XOR U7487 ( .A(n7574), .B(n7575), .Z(n7570) );
  AND U7488 ( .A(n7576), .B(n7577), .Z(n7575) );
  XNOR U7489 ( .A(p_input[1074]), .B(n7574), .Z(n7577) );
  XOR U7490 ( .A(n7574), .B(p_input[1058]), .Z(n7576) );
  XNOR U7491 ( .A(n7578), .B(n7579), .Z(n7574) );
  AND U7492 ( .A(n7580), .B(n7581), .Z(n7579) );
  XOR U7493 ( .A(p_input[1073]), .B(n7578), .Z(n7581) );
  XNOR U7494 ( .A(p_input[1057]), .B(n7578), .Z(n7580) );
  AND U7495 ( .A(p_input[1072]), .B(n7582), .Z(n7578) );
  IV U7496 ( .A(p_input[1056]), .Z(n7582) );
  XNOR U7497 ( .A(p_input[1024]), .B(n7583), .Z(n7385) );
  AND U7498 ( .A(n203), .B(n7584), .Z(n7583) );
  XOR U7499 ( .A(p_input[1040]), .B(p_input[1024]), .Z(n7584) );
  XOR U7500 ( .A(n7585), .B(n7586), .Z(n203) );
  AND U7501 ( .A(n7587), .B(n7588), .Z(n7586) );
  XNOR U7502 ( .A(p_input[1055]), .B(n7585), .Z(n7588) );
  XOR U7503 ( .A(n7585), .B(p_input[1039]), .Z(n7587) );
  XOR U7504 ( .A(n7589), .B(n7590), .Z(n7585) );
  AND U7505 ( .A(n7591), .B(n7592), .Z(n7590) );
  XNOR U7506 ( .A(p_input[1054]), .B(n7589), .Z(n7592) );
  XNOR U7507 ( .A(n7589), .B(n7399), .Z(n7591) );
  IV U7508 ( .A(p_input[1038]), .Z(n7399) );
  XOR U7509 ( .A(n7593), .B(n7594), .Z(n7589) );
  AND U7510 ( .A(n7595), .B(n7596), .Z(n7594) );
  XNOR U7511 ( .A(p_input[1053]), .B(n7593), .Z(n7596) );
  XNOR U7512 ( .A(n7593), .B(n7408), .Z(n7595) );
  IV U7513 ( .A(p_input[1037]), .Z(n7408) );
  XOR U7514 ( .A(n7597), .B(n7598), .Z(n7593) );
  AND U7515 ( .A(n7599), .B(n7600), .Z(n7598) );
  XNOR U7516 ( .A(p_input[1052]), .B(n7597), .Z(n7600) );
  XNOR U7517 ( .A(n7597), .B(n7417), .Z(n7599) );
  IV U7518 ( .A(p_input[1036]), .Z(n7417) );
  XOR U7519 ( .A(n7601), .B(n7602), .Z(n7597) );
  AND U7520 ( .A(n7603), .B(n7604), .Z(n7602) );
  XNOR U7521 ( .A(p_input[1051]), .B(n7601), .Z(n7604) );
  XNOR U7522 ( .A(n7601), .B(n7426), .Z(n7603) );
  IV U7523 ( .A(p_input[1035]), .Z(n7426) );
  XOR U7524 ( .A(n7605), .B(n7606), .Z(n7601) );
  AND U7525 ( .A(n7607), .B(n7608), .Z(n7606) );
  XNOR U7526 ( .A(p_input[1050]), .B(n7605), .Z(n7608) );
  XNOR U7527 ( .A(n7605), .B(n7435), .Z(n7607) );
  IV U7528 ( .A(p_input[1034]), .Z(n7435) );
  XOR U7529 ( .A(n7609), .B(n7610), .Z(n7605) );
  AND U7530 ( .A(n7611), .B(n7612), .Z(n7610) );
  XNOR U7531 ( .A(p_input[1049]), .B(n7609), .Z(n7612) );
  XNOR U7532 ( .A(n7609), .B(n7444), .Z(n7611) );
  IV U7533 ( .A(p_input[1033]), .Z(n7444) );
  XOR U7534 ( .A(n7613), .B(n7614), .Z(n7609) );
  AND U7535 ( .A(n7615), .B(n7616), .Z(n7614) );
  XNOR U7536 ( .A(p_input[1048]), .B(n7613), .Z(n7616) );
  XNOR U7537 ( .A(n7613), .B(n7453), .Z(n7615) );
  IV U7538 ( .A(p_input[1032]), .Z(n7453) );
  XOR U7539 ( .A(n7617), .B(n7618), .Z(n7613) );
  AND U7540 ( .A(n7619), .B(n7620), .Z(n7618) );
  XNOR U7541 ( .A(p_input[1047]), .B(n7617), .Z(n7620) );
  XNOR U7542 ( .A(n7617), .B(n7462), .Z(n7619) );
  IV U7543 ( .A(p_input[1031]), .Z(n7462) );
  XOR U7544 ( .A(n7621), .B(n7622), .Z(n7617) );
  AND U7545 ( .A(n7623), .B(n7624), .Z(n7622) );
  XNOR U7546 ( .A(p_input[1046]), .B(n7621), .Z(n7624) );
  XNOR U7547 ( .A(n7621), .B(n7471), .Z(n7623) );
  IV U7548 ( .A(p_input[1030]), .Z(n7471) );
  XOR U7549 ( .A(n7625), .B(n7626), .Z(n7621) );
  AND U7550 ( .A(n7627), .B(n7628), .Z(n7626) );
  XNOR U7551 ( .A(p_input[1045]), .B(n7625), .Z(n7628) );
  XNOR U7552 ( .A(n7625), .B(n7480), .Z(n7627) );
  IV U7553 ( .A(p_input[1029]), .Z(n7480) );
  XOR U7554 ( .A(n7629), .B(n7630), .Z(n7625) );
  AND U7555 ( .A(n7631), .B(n7632), .Z(n7630) );
  XNOR U7556 ( .A(p_input[1044]), .B(n7629), .Z(n7632) );
  XNOR U7557 ( .A(n7629), .B(n7489), .Z(n7631) );
  IV U7558 ( .A(p_input[1028]), .Z(n7489) );
  XOR U7559 ( .A(n7633), .B(n7634), .Z(n7629) );
  AND U7560 ( .A(n7635), .B(n7636), .Z(n7634) );
  XNOR U7561 ( .A(p_input[1043]), .B(n7633), .Z(n7636) );
  XNOR U7562 ( .A(n7633), .B(n7498), .Z(n7635) );
  IV U7563 ( .A(p_input[1027]), .Z(n7498) );
  XOR U7564 ( .A(n7637), .B(n7638), .Z(n7633) );
  AND U7565 ( .A(n7639), .B(n7640), .Z(n7638) );
  XNOR U7566 ( .A(p_input[1042]), .B(n7637), .Z(n7640) );
  XNOR U7567 ( .A(n7637), .B(n7507), .Z(n7639) );
  IV U7568 ( .A(p_input[1026]), .Z(n7507) );
  XNOR U7569 ( .A(n7641), .B(n7642), .Z(n7637) );
  AND U7570 ( .A(n7643), .B(n7644), .Z(n7642) );
  XOR U7571 ( .A(p_input[1041]), .B(n7641), .Z(n7644) );
  XNOR U7572 ( .A(p_input[1025]), .B(n7641), .Z(n7643) );
  AND U7573 ( .A(p_input[1040]), .B(n7645), .Z(n7641) );
  IV U7574 ( .A(p_input[1024]), .Z(n7645) );
  XOR U7575 ( .A(n7646), .B(n7647), .Z(n11) );
  AND U7576 ( .A(n551), .B(n7648), .Z(n7647) );
  XNOR U7577 ( .A(n7649), .B(n7646), .Z(n7648) );
  XOR U7578 ( .A(n7650), .B(n7651), .Z(n551) );
  AND U7579 ( .A(n7652), .B(n7653), .Z(n7651) );
  XOR U7580 ( .A(n7650), .B(n570), .Z(n7653) );
  XOR U7581 ( .A(n7654), .B(n7655), .Z(n570) );
  AND U7582 ( .A(n542), .B(n7656), .Z(n7655) );
  XOR U7583 ( .A(n7657), .B(n7654), .Z(n7656) );
  XNOR U7584 ( .A(n567), .B(n7650), .Z(n7652) );
  XOR U7585 ( .A(n7658), .B(n7659), .Z(n567) );
  AND U7586 ( .A(n539), .B(n7660), .Z(n7659) );
  XOR U7587 ( .A(n7661), .B(n7658), .Z(n7660) );
  XOR U7588 ( .A(n7662), .B(n7663), .Z(n7650) );
  AND U7589 ( .A(n7664), .B(n7665), .Z(n7663) );
  XOR U7590 ( .A(n7662), .B(n582), .Z(n7665) );
  XOR U7591 ( .A(n7666), .B(n7667), .Z(n582) );
  AND U7592 ( .A(n542), .B(n7668), .Z(n7667) );
  XOR U7593 ( .A(n7669), .B(n7666), .Z(n7668) );
  XNOR U7594 ( .A(n579), .B(n7662), .Z(n7664) );
  XOR U7595 ( .A(n7670), .B(n7671), .Z(n579) );
  AND U7596 ( .A(n539), .B(n7672), .Z(n7671) );
  XOR U7597 ( .A(n7673), .B(n7670), .Z(n7672) );
  XOR U7598 ( .A(n7674), .B(n7675), .Z(n7662) );
  AND U7599 ( .A(n7676), .B(n7677), .Z(n7675) );
  XOR U7600 ( .A(n7674), .B(n594), .Z(n7677) );
  XOR U7601 ( .A(n7678), .B(n7679), .Z(n594) );
  AND U7602 ( .A(n542), .B(n7680), .Z(n7679) );
  XOR U7603 ( .A(n7681), .B(n7678), .Z(n7680) );
  XNOR U7604 ( .A(n591), .B(n7674), .Z(n7676) );
  XOR U7605 ( .A(n7682), .B(n7683), .Z(n591) );
  AND U7606 ( .A(n539), .B(n7684), .Z(n7683) );
  XOR U7607 ( .A(n7685), .B(n7682), .Z(n7684) );
  XOR U7608 ( .A(n7686), .B(n7687), .Z(n7674) );
  AND U7609 ( .A(n7688), .B(n7689), .Z(n7687) );
  XOR U7610 ( .A(n7686), .B(n606), .Z(n7689) );
  XOR U7611 ( .A(n7690), .B(n7691), .Z(n606) );
  AND U7612 ( .A(n542), .B(n7692), .Z(n7691) );
  XOR U7613 ( .A(n7693), .B(n7690), .Z(n7692) );
  XNOR U7614 ( .A(n603), .B(n7686), .Z(n7688) );
  XOR U7615 ( .A(n7694), .B(n7695), .Z(n603) );
  AND U7616 ( .A(n539), .B(n7696), .Z(n7695) );
  XOR U7617 ( .A(n7697), .B(n7694), .Z(n7696) );
  XOR U7618 ( .A(n7698), .B(n7699), .Z(n7686) );
  AND U7619 ( .A(n7700), .B(n7701), .Z(n7699) );
  XOR U7620 ( .A(n7698), .B(n618), .Z(n7701) );
  XOR U7621 ( .A(n7702), .B(n7703), .Z(n618) );
  AND U7622 ( .A(n542), .B(n7704), .Z(n7703) );
  XOR U7623 ( .A(n7705), .B(n7702), .Z(n7704) );
  XNOR U7624 ( .A(n615), .B(n7698), .Z(n7700) );
  XOR U7625 ( .A(n7706), .B(n7707), .Z(n615) );
  AND U7626 ( .A(n539), .B(n7708), .Z(n7707) );
  XOR U7627 ( .A(n7709), .B(n7706), .Z(n7708) );
  XOR U7628 ( .A(n7710), .B(n7711), .Z(n7698) );
  AND U7629 ( .A(n7712), .B(n7713), .Z(n7711) );
  XOR U7630 ( .A(n7710), .B(n630), .Z(n7713) );
  XOR U7631 ( .A(n7714), .B(n7715), .Z(n630) );
  AND U7632 ( .A(n542), .B(n7716), .Z(n7715) );
  XOR U7633 ( .A(n7717), .B(n7714), .Z(n7716) );
  XNOR U7634 ( .A(n627), .B(n7710), .Z(n7712) );
  XOR U7635 ( .A(n7718), .B(n7719), .Z(n627) );
  AND U7636 ( .A(n539), .B(n7720), .Z(n7719) );
  XOR U7637 ( .A(n7721), .B(n7718), .Z(n7720) );
  XOR U7638 ( .A(n7722), .B(n7723), .Z(n7710) );
  AND U7639 ( .A(n7724), .B(n7725), .Z(n7723) );
  XOR U7640 ( .A(n7722), .B(n642), .Z(n7725) );
  XOR U7641 ( .A(n7726), .B(n7727), .Z(n642) );
  AND U7642 ( .A(n542), .B(n7728), .Z(n7727) );
  XOR U7643 ( .A(n7729), .B(n7726), .Z(n7728) );
  XNOR U7644 ( .A(n639), .B(n7722), .Z(n7724) );
  XOR U7645 ( .A(n7730), .B(n7731), .Z(n639) );
  AND U7646 ( .A(n539), .B(n7732), .Z(n7731) );
  XOR U7647 ( .A(n7733), .B(n7730), .Z(n7732) );
  XOR U7648 ( .A(n7734), .B(n7735), .Z(n7722) );
  AND U7649 ( .A(n7736), .B(n7737), .Z(n7735) );
  XOR U7650 ( .A(n7734), .B(n654), .Z(n7737) );
  XOR U7651 ( .A(n7738), .B(n7739), .Z(n654) );
  AND U7652 ( .A(n542), .B(n7740), .Z(n7739) );
  XOR U7653 ( .A(n7741), .B(n7738), .Z(n7740) );
  XNOR U7654 ( .A(n651), .B(n7734), .Z(n7736) );
  XOR U7655 ( .A(n7742), .B(n7743), .Z(n651) );
  AND U7656 ( .A(n539), .B(n7744), .Z(n7743) );
  XOR U7657 ( .A(n7745), .B(n7742), .Z(n7744) );
  XOR U7658 ( .A(n7746), .B(n7747), .Z(n7734) );
  AND U7659 ( .A(n7748), .B(n7749), .Z(n7747) );
  XOR U7660 ( .A(n7746), .B(n666), .Z(n7749) );
  XOR U7661 ( .A(n7750), .B(n7751), .Z(n666) );
  AND U7662 ( .A(n542), .B(n7752), .Z(n7751) );
  XOR U7663 ( .A(n7753), .B(n7750), .Z(n7752) );
  XNOR U7664 ( .A(n663), .B(n7746), .Z(n7748) );
  XOR U7665 ( .A(n7754), .B(n7755), .Z(n663) );
  AND U7666 ( .A(n539), .B(n7756), .Z(n7755) );
  XOR U7667 ( .A(n7757), .B(n7754), .Z(n7756) );
  XOR U7668 ( .A(n7758), .B(n7759), .Z(n7746) );
  AND U7669 ( .A(n7760), .B(n7761), .Z(n7759) );
  XOR U7670 ( .A(n7758), .B(n678), .Z(n7761) );
  XOR U7671 ( .A(n7762), .B(n7763), .Z(n678) );
  AND U7672 ( .A(n542), .B(n7764), .Z(n7763) );
  XOR U7673 ( .A(n7765), .B(n7762), .Z(n7764) );
  XNOR U7674 ( .A(n675), .B(n7758), .Z(n7760) );
  XOR U7675 ( .A(n7766), .B(n7767), .Z(n675) );
  AND U7676 ( .A(n539), .B(n7768), .Z(n7767) );
  XOR U7677 ( .A(n7769), .B(n7766), .Z(n7768) );
  XOR U7678 ( .A(n7770), .B(n7771), .Z(n7758) );
  AND U7679 ( .A(n7772), .B(n7773), .Z(n7771) );
  XOR U7680 ( .A(n7770), .B(n690), .Z(n7773) );
  XOR U7681 ( .A(n7774), .B(n7775), .Z(n690) );
  AND U7682 ( .A(n542), .B(n7776), .Z(n7775) );
  XOR U7683 ( .A(n7777), .B(n7774), .Z(n7776) );
  XNOR U7684 ( .A(n687), .B(n7770), .Z(n7772) );
  XOR U7685 ( .A(n7778), .B(n7779), .Z(n687) );
  AND U7686 ( .A(n539), .B(n7780), .Z(n7779) );
  XOR U7687 ( .A(n7781), .B(n7778), .Z(n7780) );
  XOR U7688 ( .A(n7782), .B(n7783), .Z(n7770) );
  AND U7689 ( .A(n7784), .B(n7785), .Z(n7783) );
  XOR U7690 ( .A(n7782), .B(n702), .Z(n7785) );
  XOR U7691 ( .A(n7786), .B(n7787), .Z(n702) );
  AND U7692 ( .A(n542), .B(n7788), .Z(n7787) );
  XOR U7693 ( .A(n7789), .B(n7786), .Z(n7788) );
  XNOR U7694 ( .A(n699), .B(n7782), .Z(n7784) );
  XOR U7695 ( .A(n7790), .B(n7791), .Z(n699) );
  AND U7696 ( .A(n539), .B(n7792), .Z(n7791) );
  XOR U7697 ( .A(n7793), .B(n7790), .Z(n7792) );
  XOR U7698 ( .A(n7794), .B(n7795), .Z(n7782) );
  AND U7699 ( .A(n7796), .B(n7797), .Z(n7795) );
  XOR U7700 ( .A(n7794), .B(n714), .Z(n7797) );
  XOR U7701 ( .A(n7798), .B(n7799), .Z(n714) );
  AND U7702 ( .A(n542), .B(n7800), .Z(n7799) );
  XOR U7703 ( .A(n7801), .B(n7798), .Z(n7800) );
  XNOR U7704 ( .A(n711), .B(n7794), .Z(n7796) );
  XOR U7705 ( .A(n7802), .B(n7803), .Z(n711) );
  AND U7706 ( .A(n539), .B(n7804), .Z(n7803) );
  XOR U7707 ( .A(n7805), .B(n7802), .Z(n7804) );
  XOR U7708 ( .A(n7806), .B(n7807), .Z(n7794) );
  AND U7709 ( .A(n7808), .B(n7809), .Z(n7807) );
  XOR U7710 ( .A(n726), .B(n7806), .Z(n7809) );
  XOR U7711 ( .A(n7810), .B(n7811), .Z(n726) );
  AND U7712 ( .A(n542), .B(n7812), .Z(n7811) );
  XOR U7713 ( .A(n7810), .B(n7813), .Z(n7812) );
  XNOR U7714 ( .A(n7806), .B(n723), .Z(n7808) );
  XOR U7715 ( .A(n7814), .B(n7815), .Z(n723) );
  AND U7716 ( .A(n539), .B(n7816), .Z(n7815) );
  XOR U7717 ( .A(n7814), .B(n7817), .Z(n7816) );
  XOR U7718 ( .A(n7818), .B(n7819), .Z(n7806) );
  AND U7719 ( .A(n7820), .B(n7821), .Z(n7819) );
  XNOR U7720 ( .A(n7822), .B(n738), .Z(n7821) );
  XOR U7721 ( .A(n7823), .B(n7824), .Z(n738) );
  AND U7722 ( .A(n542), .B(n7825), .Z(n7824) );
  XOR U7723 ( .A(n7826), .B(n7823), .Z(n7825) );
  XNOR U7724 ( .A(n735), .B(n7818), .Z(n7820) );
  XOR U7725 ( .A(n7827), .B(n7828), .Z(n735) );
  AND U7726 ( .A(n539), .B(n7829), .Z(n7828) );
  XOR U7727 ( .A(n7830), .B(n7827), .Z(n7829) );
  IV U7728 ( .A(n7822), .Z(n7818) );
  AND U7729 ( .A(n7646), .B(n7649), .Z(n7822) );
  XNOR U7730 ( .A(n7831), .B(n7832), .Z(n7649) );
  AND U7731 ( .A(n542), .B(n7833), .Z(n7832) );
  XNOR U7732 ( .A(n7834), .B(n7831), .Z(n7833) );
  XOR U7733 ( .A(n7835), .B(n7836), .Z(n542) );
  AND U7734 ( .A(n7837), .B(n7838), .Z(n7836) );
  XOR U7735 ( .A(n7835), .B(n7657), .Z(n7838) );
  XNOR U7736 ( .A(n7839), .B(n7840), .Z(n7657) );
  AND U7737 ( .A(n7841), .B(n510), .Z(n7840) );
  AND U7738 ( .A(n7839), .B(n7842), .Z(n7841) );
  XNOR U7739 ( .A(n7654), .B(n7835), .Z(n7837) );
  XOR U7740 ( .A(n7843), .B(n7844), .Z(n7654) );
  AND U7741 ( .A(n7845), .B(n508), .Z(n7844) );
  NOR U7742 ( .A(n7843), .B(n7846), .Z(n7845) );
  XOR U7743 ( .A(n7847), .B(n7848), .Z(n7835) );
  AND U7744 ( .A(n7849), .B(n7850), .Z(n7848) );
  XOR U7745 ( .A(n7847), .B(n7669), .Z(n7850) );
  XOR U7746 ( .A(n7851), .B(n7852), .Z(n7669) );
  AND U7747 ( .A(n510), .B(n7853), .Z(n7852) );
  XOR U7748 ( .A(n7854), .B(n7851), .Z(n7853) );
  XNOR U7749 ( .A(n7666), .B(n7847), .Z(n7849) );
  XOR U7750 ( .A(n7855), .B(n7856), .Z(n7666) );
  AND U7751 ( .A(n508), .B(n7857), .Z(n7856) );
  XOR U7752 ( .A(n7858), .B(n7855), .Z(n7857) );
  XOR U7753 ( .A(n7859), .B(n7860), .Z(n7847) );
  AND U7754 ( .A(n7861), .B(n7862), .Z(n7860) );
  XOR U7755 ( .A(n7859), .B(n7681), .Z(n7862) );
  XOR U7756 ( .A(n7863), .B(n7864), .Z(n7681) );
  AND U7757 ( .A(n510), .B(n7865), .Z(n7864) );
  XOR U7758 ( .A(n7866), .B(n7863), .Z(n7865) );
  XNOR U7759 ( .A(n7678), .B(n7859), .Z(n7861) );
  XOR U7760 ( .A(n7867), .B(n7868), .Z(n7678) );
  AND U7761 ( .A(n508), .B(n7869), .Z(n7868) );
  XOR U7762 ( .A(n7870), .B(n7867), .Z(n7869) );
  XOR U7763 ( .A(n7871), .B(n7872), .Z(n7859) );
  AND U7764 ( .A(n7873), .B(n7874), .Z(n7872) );
  XOR U7765 ( .A(n7871), .B(n7693), .Z(n7874) );
  XOR U7766 ( .A(n7875), .B(n7876), .Z(n7693) );
  AND U7767 ( .A(n510), .B(n7877), .Z(n7876) );
  XOR U7768 ( .A(n7878), .B(n7875), .Z(n7877) );
  XNOR U7769 ( .A(n7690), .B(n7871), .Z(n7873) );
  XOR U7770 ( .A(n7879), .B(n7880), .Z(n7690) );
  AND U7771 ( .A(n508), .B(n7881), .Z(n7880) );
  XOR U7772 ( .A(n7882), .B(n7879), .Z(n7881) );
  XOR U7773 ( .A(n7883), .B(n7884), .Z(n7871) );
  AND U7774 ( .A(n7885), .B(n7886), .Z(n7884) );
  XOR U7775 ( .A(n7883), .B(n7705), .Z(n7886) );
  XOR U7776 ( .A(n7887), .B(n7888), .Z(n7705) );
  AND U7777 ( .A(n510), .B(n7889), .Z(n7888) );
  XOR U7778 ( .A(n7890), .B(n7887), .Z(n7889) );
  XNOR U7779 ( .A(n7702), .B(n7883), .Z(n7885) );
  XOR U7780 ( .A(n7891), .B(n7892), .Z(n7702) );
  AND U7781 ( .A(n508), .B(n7893), .Z(n7892) );
  XOR U7782 ( .A(n7894), .B(n7891), .Z(n7893) );
  XOR U7783 ( .A(n7895), .B(n7896), .Z(n7883) );
  AND U7784 ( .A(n7897), .B(n7898), .Z(n7896) );
  XOR U7785 ( .A(n7895), .B(n7717), .Z(n7898) );
  XOR U7786 ( .A(n7899), .B(n7900), .Z(n7717) );
  AND U7787 ( .A(n510), .B(n7901), .Z(n7900) );
  XOR U7788 ( .A(n7902), .B(n7899), .Z(n7901) );
  XNOR U7789 ( .A(n7714), .B(n7895), .Z(n7897) );
  XOR U7790 ( .A(n7903), .B(n7904), .Z(n7714) );
  AND U7791 ( .A(n508), .B(n7905), .Z(n7904) );
  XOR U7792 ( .A(n7906), .B(n7903), .Z(n7905) );
  XOR U7793 ( .A(n7907), .B(n7908), .Z(n7895) );
  AND U7794 ( .A(n7909), .B(n7910), .Z(n7908) );
  XOR U7795 ( .A(n7907), .B(n7729), .Z(n7910) );
  XOR U7796 ( .A(n7911), .B(n7912), .Z(n7729) );
  AND U7797 ( .A(n510), .B(n7913), .Z(n7912) );
  XOR U7798 ( .A(n7914), .B(n7911), .Z(n7913) );
  XNOR U7799 ( .A(n7726), .B(n7907), .Z(n7909) );
  XOR U7800 ( .A(n7915), .B(n7916), .Z(n7726) );
  AND U7801 ( .A(n508), .B(n7917), .Z(n7916) );
  XOR U7802 ( .A(n7918), .B(n7915), .Z(n7917) );
  XOR U7803 ( .A(n7919), .B(n7920), .Z(n7907) );
  AND U7804 ( .A(n7921), .B(n7922), .Z(n7920) );
  XOR U7805 ( .A(n7919), .B(n7741), .Z(n7922) );
  XOR U7806 ( .A(n7923), .B(n7924), .Z(n7741) );
  AND U7807 ( .A(n510), .B(n7925), .Z(n7924) );
  XOR U7808 ( .A(n7926), .B(n7923), .Z(n7925) );
  XNOR U7809 ( .A(n7738), .B(n7919), .Z(n7921) );
  XOR U7810 ( .A(n7927), .B(n7928), .Z(n7738) );
  AND U7811 ( .A(n508), .B(n7929), .Z(n7928) );
  XOR U7812 ( .A(n7930), .B(n7927), .Z(n7929) );
  XOR U7813 ( .A(n7931), .B(n7932), .Z(n7919) );
  AND U7814 ( .A(n7933), .B(n7934), .Z(n7932) );
  XOR U7815 ( .A(n7931), .B(n7753), .Z(n7934) );
  XOR U7816 ( .A(n7935), .B(n7936), .Z(n7753) );
  AND U7817 ( .A(n510), .B(n7937), .Z(n7936) );
  XOR U7818 ( .A(n7938), .B(n7935), .Z(n7937) );
  XNOR U7819 ( .A(n7750), .B(n7931), .Z(n7933) );
  XOR U7820 ( .A(n7939), .B(n7940), .Z(n7750) );
  AND U7821 ( .A(n508), .B(n7941), .Z(n7940) );
  XOR U7822 ( .A(n7942), .B(n7939), .Z(n7941) );
  XOR U7823 ( .A(n7943), .B(n7944), .Z(n7931) );
  AND U7824 ( .A(n7945), .B(n7946), .Z(n7944) );
  XOR U7825 ( .A(n7943), .B(n7765), .Z(n7946) );
  XOR U7826 ( .A(n7947), .B(n7948), .Z(n7765) );
  AND U7827 ( .A(n510), .B(n7949), .Z(n7948) );
  XOR U7828 ( .A(n7950), .B(n7947), .Z(n7949) );
  XNOR U7829 ( .A(n7762), .B(n7943), .Z(n7945) );
  XOR U7830 ( .A(n7951), .B(n7952), .Z(n7762) );
  AND U7831 ( .A(n508), .B(n7953), .Z(n7952) );
  XOR U7832 ( .A(n7954), .B(n7951), .Z(n7953) );
  XOR U7833 ( .A(n7955), .B(n7956), .Z(n7943) );
  AND U7834 ( .A(n7957), .B(n7958), .Z(n7956) );
  XOR U7835 ( .A(n7955), .B(n7777), .Z(n7958) );
  XOR U7836 ( .A(n7959), .B(n7960), .Z(n7777) );
  AND U7837 ( .A(n510), .B(n7961), .Z(n7960) );
  XOR U7838 ( .A(n7962), .B(n7959), .Z(n7961) );
  XNOR U7839 ( .A(n7774), .B(n7955), .Z(n7957) );
  XOR U7840 ( .A(n7963), .B(n7964), .Z(n7774) );
  AND U7841 ( .A(n508), .B(n7965), .Z(n7964) );
  XOR U7842 ( .A(n7966), .B(n7963), .Z(n7965) );
  XOR U7843 ( .A(n7967), .B(n7968), .Z(n7955) );
  AND U7844 ( .A(n7969), .B(n7970), .Z(n7968) );
  XOR U7845 ( .A(n7967), .B(n7789), .Z(n7970) );
  XOR U7846 ( .A(n7971), .B(n7972), .Z(n7789) );
  AND U7847 ( .A(n510), .B(n7973), .Z(n7972) );
  XOR U7848 ( .A(n7974), .B(n7971), .Z(n7973) );
  XNOR U7849 ( .A(n7786), .B(n7967), .Z(n7969) );
  XOR U7850 ( .A(n7975), .B(n7976), .Z(n7786) );
  AND U7851 ( .A(n508), .B(n7977), .Z(n7976) );
  XOR U7852 ( .A(n7978), .B(n7975), .Z(n7977) );
  XOR U7853 ( .A(n7979), .B(n7980), .Z(n7967) );
  AND U7854 ( .A(n7981), .B(n7982), .Z(n7980) );
  XOR U7855 ( .A(n7979), .B(n7801), .Z(n7982) );
  XOR U7856 ( .A(n7983), .B(n7984), .Z(n7801) );
  AND U7857 ( .A(n510), .B(n7985), .Z(n7984) );
  XOR U7858 ( .A(n7986), .B(n7983), .Z(n7985) );
  XNOR U7859 ( .A(n7798), .B(n7979), .Z(n7981) );
  XOR U7860 ( .A(n7987), .B(n7988), .Z(n7798) );
  AND U7861 ( .A(n508), .B(n7989), .Z(n7988) );
  XOR U7862 ( .A(n7990), .B(n7987), .Z(n7989) );
  XOR U7863 ( .A(n7991), .B(n7992), .Z(n7979) );
  AND U7864 ( .A(n7993), .B(n7994), .Z(n7992) );
  XOR U7865 ( .A(n7813), .B(n7991), .Z(n7994) );
  XOR U7866 ( .A(n7995), .B(n7996), .Z(n7813) );
  AND U7867 ( .A(n510), .B(n7997), .Z(n7996) );
  XOR U7868 ( .A(n7995), .B(n7998), .Z(n7997) );
  XNOR U7869 ( .A(n7991), .B(n7810), .Z(n7993) );
  XOR U7870 ( .A(n7999), .B(n8000), .Z(n7810) );
  AND U7871 ( .A(n508), .B(n8001), .Z(n8000) );
  XOR U7872 ( .A(n7999), .B(n8002), .Z(n8001) );
  XOR U7873 ( .A(n8003), .B(n8004), .Z(n7991) );
  AND U7874 ( .A(n8005), .B(n8006), .Z(n8004) );
  XNOR U7875 ( .A(n8007), .B(n7826), .Z(n8006) );
  XOR U7876 ( .A(n8008), .B(n8009), .Z(n7826) );
  AND U7877 ( .A(n510), .B(n8010), .Z(n8009) );
  XOR U7878 ( .A(n8011), .B(n8008), .Z(n8010) );
  XNOR U7879 ( .A(n7823), .B(n8003), .Z(n8005) );
  XOR U7880 ( .A(n8012), .B(n8013), .Z(n7823) );
  AND U7881 ( .A(n508), .B(n8014), .Z(n8013) );
  XOR U7882 ( .A(n8015), .B(n8012), .Z(n8014) );
  IV U7883 ( .A(n8007), .Z(n8003) );
  AND U7884 ( .A(n7831), .B(n7834), .Z(n8007) );
  XNOR U7885 ( .A(n8016), .B(n8017), .Z(n7834) );
  AND U7886 ( .A(n510), .B(n8018), .Z(n8017) );
  XNOR U7887 ( .A(n8019), .B(n8016), .Z(n8018) );
  XOR U7888 ( .A(n8020), .B(n8021), .Z(n510) );
  AND U7889 ( .A(n8022), .B(n8023), .Z(n8021) );
  XOR U7890 ( .A(n7842), .B(n8020), .Z(n8023) );
  IV U7891 ( .A(n8024), .Z(n7842) );
  AND U7892 ( .A(n8025), .B(n8026), .Z(n8024) );
  XOR U7893 ( .A(n8020), .B(n7839), .Z(n8022) );
  AND U7894 ( .A(n8027), .B(n8028), .Z(n7839) );
  XOR U7895 ( .A(n8029), .B(n8030), .Z(n8020) );
  AND U7896 ( .A(n8031), .B(n8032), .Z(n8030) );
  XOR U7897 ( .A(n8029), .B(n7854), .Z(n8032) );
  XOR U7898 ( .A(n8033), .B(n8034), .Z(n7854) );
  AND U7899 ( .A(n438), .B(n8035), .Z(n8034) );
  XOR U7900 ( .A(n8036), .B(n8033), .Z(n8035) );
  XNOR U7901 ( .A(n7851), .B(n8029), .Z(n8031) );
  XOR U7902 ( .A(n8037), .B(n8038), .Z(n7851) );
  AND U7903 ( .A(n436), .B(n8039), .Z(n8038) );
  XOR U7904 ( .A(n8040), .B(n8037), .Z(n8039) );
  XOR U7905 ( .A(n8041), .B(n8042), .Z(n8029) );
  AND U7906 ( .A(n8043), .B(n8044), .Z(n8042) );
  XOR U7907 ( .A(n8041), .B(n7866), .Z(n8044) );
  XOR U7908 ( .A(n8045), .B(n8046), .Z(n7866) );
  AND U7909 ( .A(n438), .B(n8047), .Z(n8046) );
  XOR U7910 ( .A(n8048), .B(n8045), .Z(n8047) );
  XNOR U7911 ( .A(n7863), .B(n8041), .Z(n8043) );
  XOR U7912 ( .A(n8049), .B(n8050), .Z(n7863) );
  AND U7913 ( .A(n436), .B(n8051), .Z(n8050) );
  XOR U7914 ( .A(n8052), .B(n8049), .Z(n8051) );
  XOR U7915 ( .A(n8053), .B(n8054), .Z(n8041) );
  AND U7916 ( .A(n8055), .B(n8056), .Z(n8054) );
  XOR U7917 ( .A(n8053), .B(n7878), .Z(n8056) );
  XOR U7918 ( .A(n8057), .B(n8058), .Z(n7878) );
  AND U7919 ( .A(n438), .B(n8059), .Z(n8058) );
  XOR U7920 ( .A(n8060), .B(n8057), .Z(n8059) );
  XNOR U7921 ( .A(n7875), .B(n8053), .Z(n8055) );
  XOR U7922 ( .A(n8061), .B(n8062), .Z(n7875) );
  AND U7923 ( .A(n436), .B(n8063), .Z(n8062) );
  XOR U7924 ( .A(n8064), .B(n8061), .Z(n8063) );
  XOR U7925 ( .A(n8065), .B(n8066), .Z(n8053) );
  AND U7926 ( .A(n8067), .B(n8068), .Z(n8066) );
  XOR U7927 ( .A(n8065), .B(n7890), .Z(n8068) );
  XOR U7928 ( .A(n8069), .B(n8070), .Z(n7890) );
  AND U7929 ( .A(n438), .B(n8071), .Z(n8070) );
  XOR U7930 ( .A(n8072), .B(n8069), .Z(n8071) );
  XNOR U7931 ( .A(n7887), .B(n8065), .Z(n8067) );
  XOR U7932 ( .A(n8073), .B(n8074), .Z(n7887) );
  AND U7933 ( .A(n436), .B(n8075), .Z(n8074) );
  XOR U7934 ( .A(n8076), .B(n8073), .Z(n8075) );
  XOR U7935 ( .A(n8077), .B(n8078), .Z(n8065) );
  AND U7936 ( .A(n8079), .B(n8080), .Z(n8078) );
  XOR U7937 ( .A(n8077), .B(n7902), .Z(n8080) );
  XOR U7938 ( .A(n8081), .B(n8082), .Z(n7902) );
  AND U7939 ( .A(n438), .B(n8083), .Z(n8082) );
  XOR U7940 ( .A(n8084), .B(n8081), .Z(n8083) );
  XNOR U7941 ( .A(n7899), .B(n8077), .Z(n8079) );
  XOR U7942 ( .A(n8085), .B(n8086), .Z(n7899) );
  AND U7943 ( .A(n436), .B(n8087), .Z(n8086) );
  XOR U7944 ( .A(n8088), .B(n8085), .Z(n8087) );
  XOR U7945 ( .A(n8089), .B(n8090), .Z(n8077) );
  AND U7946 ( .A(n8091), .B(n8092), .Z(n8090) );
  XOR U7947 ( .A(n8089), .B(n7914), .Z(n8092) );
  XOR U7948 ( .A(n8093), .B(n8094), .Z(n7914) );
  AND U7949 ( .A(n438), .B(n8095), .Z(n8094) );
  XOR U7950 ( .A(n8096), .B(n8093), .Z(n8095) );
  XNOR U7951 ( .A(n7911), .B(n8089), .Z(n8091) );
  XOR U7952 ( .A(n8097), .B(n8098), .Z(n7911) );
  AND U7953 ( .A(n436), .B(n8099), .Z(n8098) );
  XOR U7954 ( .A(n8100), .B(n8097), .Z(n8099) );
  XOR U7955 ( .A(n8101), .B(n8102), .Z(n8089) );
  AND U7956 ( .A(n8103), .B(n8104), .Z(n8102) );
  XOR U7957 ( .A(n8101), .B(n7926), .Z(n8104) );
  XOR U7958 ( .A(n8105), .B(n8106), .Z(n7926) );
  AND U7959 ( .A(n438), .B(n8107), .Z(n8106) );
  XOR U7960 ( .A(n8108), .B(n8105), .Z(n8107) );
  XNOR U7961 ( .A(n7923), .B(n8101), .Z(n8103) );
  XOR U7962 ( .A(n8109), .B(n8110), .Z(n7923) );
  AND U7963 ( .A(n436), .B(n8111), .Z(n8110) );
  XOR U7964 ( .A(n8112), .B(n8109), .Z(n8111) );
  XOR U7965 ( .A(n8113), .B(n8114), .Z(n8101) );
  AND U7966 ( .A(n8115), .B(n8116), .Z(n8114) );
  XOR U7967 ( .A(n8113), .B(n7938), .Z(n8116) );
  XOR U7968 ( .A(n8117), .B(n8118), .Z(n7938) );
  AND U7969 ( .A(n438), .B(n8119), .Z(n8118) );
  XOR U7970 ( .A(n8120), .B(n8117), .Z(n8119) );
  XNOR U7971 ( .A(n7935), .B(n8113), .Z(n8115) );
  XOR U7972 ( .A(n8121), .B(n8122), .Z(n7935) );
  AND U7973 ( .A(n436), .B(n8123), .Z(n8122) );
  XOR U7974 ( .A(n8124), .B(n8121), .Z(n8123) );
  XOR U7975 ( .A(n8125), .B(n8126), .Z(n8113) );
  AND U7976 ( .A(n8127), .B(n8128), .Z(n8126) );
  XOR U7977 ( .A(n8125), .B(n7950), .Z(n8128) );
  XOR U7978 ( .A(n8129), .B(n8130), .Z(n7950) );
  AND U7979 ( .A(n438), .B(n8131), .Z(n8130) );
  XOR U7980 ( .A(n8132), .B(n8129), .Z(n8131) );
  XNOR U7981 ( .A(n7947), .B(n8125), .Z(n8127) );
  XOR U7982 ( .A(n8133), .B(n8134), .Z(n7947) );
  AND U7983 ( .A(n436), .B(n8135), .Z(n8134) );
  XOR U7984 ( .A(n8136), .B(n8133), .Z(n8135) );
  XOR U7985 ( .A(n8137), .B(n8138), .Z(n8125) );
  AND U7986 ( .A(n8139), .B(n8140), .Z(n8138) );
  XOR U7987 ( .A(n8137), .B(n7962), .Z(n8140) );
  XOR U7988 ( .A(n8141), .B(n8142), .Z(n7962) );
  AND U7989 ( .A(n438), .B(n8143), .Z(n8142) );
  XOR U7990 ( .A(n8144), .B(n8141), .Z(n8143) );
  XNOR U7991 ( .A(n7959), .B(n8137), .Z(n8139) );
  XOR U7992 ( .A(n8145), .B(n8146), .Z(n7959) );
  AND U7993 ( .A(n436), .B(n8147), .Z(n8146) );
  XOR U7994 ( .A(n8148), .B(n8145), .Z(n8147) );
  XOR U7995 ( .A(n8149), .B(n8150), .Z(n8137) );
  AND U7996 ( .A(n8151), .B(n8152), .Z(n8150) );
  XOR U7997 ( .A(n8149), .B(n7974), .Z(n8152) );
  XOR U7998 ( .A(n8153), .B(n8154), .Z(n7974) );
  AND U7999 ( .A(n438), .B(n8155), .Z(n8154) );
  XOR U8000 ( .A(n8156), .B(n8153), .Z(n8155) );
  XNOR U8001 ( .A(n7971), .B(n8149), .Z(n8151) );
  XOR U8002 ( .A(n8157), .B(n8158), .Z(n7971) );
  AND U8003 ( .A(n436), .B(n8159), .Z(n8158) );
  XOR U8004 ( .A(n8160), .B(n8157), .Z(n8159) );
  XOR U8005 ( .A(n8161), .B(n8162), .Z(n8149) );
  AND U8006 ( .A(n8163), .B(n8164), .Z(n8162) );
  XOR U8007 ( .A(n8161), .B(n7986), .Z(n8164) );
  XOR U8008 ( .A(n8165), .B(n8166), .Z(n7986) );
  AND U8009 ( .A(n438), .B(n8167), .Z(n8166) );
  XOR U8010 ( .A(n8168), .B(n8165), .Z(n8167) );
  XNOR U8011 ( .A(n7983), .B(n8161), .Z(n8163) );
  XOR U8012 ( .A(n8169), .B(n8170), .Z(n7983) );
  AND U8013 ( .A(n436), .B(n8171), .Z(n8170) );
  XOR U8014 ( .A(n8172), .B(n8169), .Z(n8171) );
  XOR U8015 ( .A(n8173), .B(n8174), .Z(n8161) );
  AND U8016 ( .A(n8175), .B(n8176), .Z(n8174) );
  XOR U8017 ( .A(n7998), .B(n8173), .Z(n8176) );
  XOR U8018 ( .A(n8177), .B(n8178), .Z(n7998) );
  AND U8019 ( .A(n438), .B(n8179), .Z(n8178) );
  XOR U8020 ( .A(n8177), .B(n8180), .Z(n8179) );
  XNOR U8021 ( .A(n8173), .B(n7995), .Z(n8175) );
  XOR U8022 ( .A(n8181), .B(n8182), .Z(n7995) );
  AND U8023 ( .A(n436), .B(n8183), .Z(n8182) );
  XOR U8024 ( .A(n8181), .B(n8184), .Z(n8183) );
  XOR U8025 ( .A(n8185), .B(n8186), .Z(n8173) );
  AND U8026 ( .A(n8187), .B(n8188), .Z(n8186) );
  XNOR U8027 ( .A(n8189), .B(n8011), .Z(n8188) );
  XOR U8028 ( .A(n8190), .B(n8191), .Z(n8011) );
  AND U8029 ( .A(n438), .B(n8192), .Z(n8191) );
  XOR U8030 ( .A(n8193), .B(n8190), .Z(n8192) );
  XNOR U8031 ( .A(n8008), .B(n8185), .Z(n8187) );
  XOR U8032 ( .A(n8194), .B(n8195), .Z(n8008) );
  AND U8033 ( .A(n436), .B(n8196), .Z(n8195) );
  XOR U8034 ( .A(n8197), .B(n8194), .Z(n8196) );
  IV U8035 ( .A(n8189), .Z(n8185) );
  AND U8036 ( .A(n8016), .B(n8019), .Z(n8189) );
  XNOR U8037 ( .A(n8198), .B(n8199), .Z(n8019) );
  AND U8038 ( .A(n438), .B(n8200), .Z(n8199) );
  XNOR U8039 ( .A(n8201), .B(n8198), .Z(n8200) );
  XOR U8040 ( .A(n8202), .B(n8203), .Z(n438) );
  AND U8041 ( .A(n8204), .B(n8205), .Z(n8203) );
  XNOR U8042 ( .A(n8025), .B(n8202), .Z(n8205) );
  AND U8043 ( .A(n8206), .B(n8207), .Z(n8025) );
  XOR U8044 ( .A(n8202), .B(n8026), .Z(n8204) );
  AND U8045 ( .A(n8208), .B(n8209), .Z(n8026) );
  XOR U8046 ( .A(n8210), .B(n8211), .Z(n8202) );
  AND U8047 ( .A(n8212), .B(n8213), .Z(n8211) );
  XOR U8048 ( .A(n8210), .B(n8036), .Z(n8213) );
  XOR U8049 ( .A(n8214), .B(n8215), .Z(n8036) );
  AND U8050 ( .A(n286), .B(n8216), .Z(n8215) );
  XOR U8051 ( .A(n8217), .B(n8214), .Z(n8216) );
  XNOR U8052 ( .A(n8033), .B(n8210), .Z(n8212) );
  XOR U8053 ( .A(n8218), .B(n8219), .Z(n8033) );
  AND U8054 ( .A(n284), .B(n8220), .Z(n8219) );
  XOR U8055 ( .A(n8221), .B(n8218), .Z(n8220) );
  XOR U8056 ( .A(n8222), .B(n8223), .Z(n8210) );
  AND U8057 ( .A(n8224), .B(n8225), .Z(n8223) );
  XOR U8058 ( .A(n8222), .B(n8048), .Z(n8225) );
  XOR U8059 ( .A(n8226), .B(n8227), .Z(n8048) );
  AND U8060 ( .A(n286), .B(n8228), .Z(n8227) );
  XOR U8061 ( .A(n8229), .B(n8226), .Z(n8228) );
  XNOR U8062 ( .A(n8045), .B(n8222), .Z(n8224) );
  XOR U8063 ( .A(n8230), .B(n8231), .Z(n8045) );
  AND U8064 ( .A(n284), .B(n8232), .Z(n8231) );
  XOR U8065 ( .A(n8233), .B(n8230), .Z(n8232) );
  XOR U8066 ( .A(n8234), .B(n8235), .Z(n8222) );
  AND U8067 ( .A(n8236), .B(n8237), .Z(n8235) );
  XOR U8068 ( .A(n8234), .B(n8060), .Z(n8237) );
  XOR U8069 ( .A(n8238), .B(n8239), .Z(n8060) );
  AND U8070 ( .A(n286), .B(n8240), .Z(n8239) );
  XOR U8071 ( .A(n8241), .B(n8238), .Z(n8240) );
  XNOR U8072 ( .A(n8057), .B(n8234), .Z(n8236) );
  XOR U8073 ( .A(n8242), .B(n8243), .Z(n8057) );
  AND U8074 ( .A(n284), .B(n8244), .Z(n8243) );
  XOR U8075 ( .A(n8245), .B(n8242), .Z(n8244) );
  XOR U8076 ( .A(n8246), .B(n8247), .Z(n8234) );
  AND U8077 ( .A(n8248), .B(n8249), .Z(n8247) );
  XOR U8078 ( .A(n8246), .B(n8072), .Z(n8249) );
  XOR U8079 ( .A(n8250), .B(n8251), .Z(n8072) );
  AND U8080 ( .A(n286), .B(n8252), .Z(n8251) );
  XOR U8081 ( .A(n8253), .B(n8250), .Z(n8252) );
  XNOR U8082 ( .A(n8069), .B(n8246), .Z(n8248) );
  XOR U8083 ( .A(n8254), .B(n8255), .Z(n8069) );
  AND U8084 ( .A(n284), .B(n8256), .Z(n8255) );
  XOR U8085 ( .A(n8257), .B(n8254), .Z(n8256) );
  XOR U8086 ( .A(n8258), .B(n8259), .Z(n8246) );
  AND U8087 ( .A(n8260), .B(n8261), .Z(n8259) );
  XOR U8088 ( .A(n8258), .B(n8084), .Z(n8261) );
  XOR U8089 ( .A(n8262), .B(n8263), .Z(n8084) );
  AND U8090 ( .A(n286), .B(n8264), .Z(n8263) );
  XOR U8091 ( .A(n8265), .B(n8262), .Z(n8264) );
  XNOR U8092 ( .A(n8081), .B(n8258), .Z(n8260) );
  XOR U8093 ( .A(n8266), .B(n8267), .Z(n8081) );
  AND U8094 ( .A(n284), .B(n8268), .Z(n8267) );
  XOR U8095 ( .A(n8269), .B(n8266), .Z(n8268) );
  XOR U8096 ( .A(n8270), .B(n8271), .Z(n8258) );
  AND U8097 ( .A(n8272), .B(n8273), .Z(n8271) );
  XOR U8098 ( .A(n8270), .B(n8096), .Z(n8273) );
  XOR U8099 ( .A(n8274), .B(n8275), .Z(n8096) );
  AND U8100 ( .A(n286), .B(n8276), .Z(n8275) );
  XOR U8101 ( .A(n8277), .B(n8274), .Z(n8276) );
  XNOR U8102 ( .A(n8093), .B(n8270), .Z(n8272) );
  XOR U8103 ( .A(n8278), .B(n8279), .Z(n8093) );
  AND U8104 ( .A(n284), .B(n8280), .Z(n8279) );
  XOR U8105 ( .A(n8281), .B(n8278), .Z(n8280) );
  XOR U8106 ( .A(n8282), .B(n8283), .Z(n8270) );
  AND U8107 ( .A(n8284), .B(n8285), .Z(n8283) );
  XOR U8108 ( .A(n8282), .B(n8108), .Z(n8285) );
  XOR U8109 ( .A(n8286), .B(n8287), .Z(n8108) );
  AND U8110 ( .A(n286), .B(n8288), .Z(n8287) );
  XOR U8111 ( .A(n8289), .B(n8286), .Z(n8288) );
  XNOR U8112 ( .A(n8105), .B(n8282), .Z(n8284) );
  XOR U8113 ( .A(n8290), .B(n8291), .Z(n8105) );
  AND U8114 ( .A(n284), .B(n8292), .Z(n8291) );
  XOR U8115 ( .A(n8293), .B(n8290), .Z(n8292) );
  XOR U8116 ( .A(n8294), .B(n8295), .Z(n8282) );
  AND U8117 ( .A(n8296), .B(n8297), .Z(n8295) );
  XOR U8118 ( .A(n8294), .B(n8120), .Z(n8297) );
  XOR U8119 ( .A(n8298), .B(n8299), .Z(n8120) );
  AND U8120 ( .A(n286), .B(n8300), .Z(n8299) );
  XOR U8121 ( .A(n8301), .B(n8298), .Z(n8300) );
  XNOR U8122 ( .A(n8117), .B(n8294), .Z(n8296) );
  XOR U8123 ( .A(n8302), .B(n8303), .Z(n8117) );
  AND U8124 ( .A(n284), .B(n8304), .Z(n8303) );
  XOR U8125 ( .A(n8305), .B(n8302), .Z(n8304) );
  XOR U8126 ( .A(n8306), .B(n8307), .Z(n8294) );
  AND U8127 ( .A(n8308), .B(n8309), .Z(n8307) );
  XOR U8128 ( .A(n8306), .B(n8132), .Z(n8309) );
  XOR U8129 ( .A(n8310), .B(n8311), .Z(n8132) );
  AND U8130 ( .A(n286), .B(n8312), .Z(n8311) );
  XOR U8131 ( .A(n8313), .B(n8310), .Z(n8312) );
  XNOR U8132 ( .A(n8129), .B(n8306), .Z(n8308) );
  XOR U8133 ( .A(n8314), .B(n8315), .Z(n8129) );
  AND U8134 ( .A(n284), .B(n8316), .Z(n8315) );
  XOR U8135 ( .A(n8317), .B(n8314), .Z(n8316) );
  XOR U8136 ( .A(n8318), .B(n8319), .Z(n8306) );
  AND U8137 ( .A(n8320), .B(n8321), .Z(n8319) );
  XOR U8138 ( .A(n8318), .B(n8144), .Z(n8321) );
  XOR U8139 ( .A(n8322), .B(n8323), .Z(n8144) );
  AND U8140 ( .A(n286), .B(n8324), .Z(n8323) );
  XOR U8141 ( .A(n8325), .B(n8322), .Z(n8324) );
  XNOR U8142 ( .A(n8141), .B(n8318), .Z(n8320) );
  XOR U8143 ( .A(n8326), .B(n8327), .Z(n8141) );
  AND U8144 ( .A(n284), .B(n8328), .Z(n8327) );
  XOR U8145 ( .A(n8329), .B(n8326), .Z(n8328) );
  XOR U8146 ( .A(n8330), .B(n8331), .Z(n8318) );
  AND U8147 ( .A(n8332), .B(n8333), .Z(n8331) );
  XOR U8148 ( .A(n8330), .B(n8156), .Z(n8333) );
  XOR U8149 ( .A(n8334), .B(n8335), .Z(n8156) );
  AND U8150 ( .A(n286), .B(n8336), .Z(n8335) );
  XOR U8151 ( .A(n8337), .B(n8334), .Z(n8336) );
  XNOR U8152 ( .A(n8153), .B(n8330), .Z(n8332) );
  XOR U8153 ( .A(n8338), .B(n8339), .Z(n8153) );
  AND U8154 ( .A(n284), .B(n8340), .Z(n8339) );
  XOR U8155 ( .A(n8341), .B(n8338), .Z(n8340) );
  XOR U8156 ( .A(n8342), .B(n8343), .Z(n8330) );
  AND U8157 ( .A(n8344), .B(n8345), .Z(n8343) );
  XOR U8158 ( .A(n8342), .B(n8168), .Z(n8345) );
  XOR U8159 ( .A(n8346), .B(n8347), .Z(n8168) );
  AND U8160 ( .A(n286), .B(n8348), .Z(n8347) );
  XOR U8161 ( .A(n8349), .B(n8346), .Z(n8348) );
  XNOR U8162 ( .A(n8165), .B(n8342), .Z(n8344) );
  XOR U8163 ( .A(n8350), .B(n8351), .Z(n8165) );
  AND U8164 ( .A(n284), .B(n8352), .Z(n8351) );
  XOR U8165 ( .A(n8353), .B(n8350), .Z(n8352) );
  XOR U8166 ( .A(n8354), .B(n8355), .Z(n8342) );
  AND U8167 ( .A(n8356), .B(n8357), .Z(n8355) );
  XOR U8168 ( .A(n8180), .B(n8354), .Z(n8357) );
  XOR U8169 ( .A(n8358), .B(n8359), .Z(n8180) );
  AND U8170 ( .A(n286), .B(n8360), .Z(n8359) );
  XOR U8171 ( .A(n8358), .B(n8361), .Z(n8360) );
  XNOR U8172 ( .A(n8354), .B(n8177), .Z(n8356) );
  XOR U8173 ( .A(n8362), .B(n8363), .Z(n8177) );
  AND U8174 ( .A(n284), .B(n8364), .Z(n8363) );
  XOR U8175 ( .A(n8362), .B(n8365), .Z(n8364) );
  XOR U8176 ( .A(n8366), .B(n8367), .Z(n8354) );
  AND U8177 ( .A(n8368), .B(n8369), .Z(n8367) );
  XNOR U8178 ( .A(n8370), .B(n8193), .Z(n8369) );
  XOR U8179 ( .A(n8371), .B(n8372), .Z(n8193) );
  AND U8180 ( .A(n286), .B(n8373), .Z(n8372) );
  XOR U8181 ( .A(n8374), .B(n8371), .Z(n8373) );
  XNOR U8182 ( .A(n8190), .B(n8366), .Z(n8368) );
  XOR U8183 ( .A(n8375), .B(n8376), .Z(n8190) );
  AND U8184 ( .A(n284), .B(n8377), .Z(n8376) );
  XOR U8185 ( .A(n8378), .B(n8375), .Z(n8377) );
  IV U8186 ( .A(n8370), .Z(n8366) );
  AND U8187 ( .A(n8198), .B(n8201), .Z(n8370) );
  XNOR U8188 ( .A(n8379), .B(n8380), .Z(n8201) );
  AND U8189 ( .A(n286), .B(n8381), .Z(n8380) );
  XNOR U8190 ( .A(n8382), .B(n8379), .Z(n8381) );
  XOR U8191 ( .A(n8383), .B(n8384), .Z(n286) );
  AND U8192 ( .A(n8385), .B(n8386), .Z(n8384) );
  XNOR U8193 ( .A(n8206), .B(n8383), .Z(n8386) );
  AND U8194 ( .A(p_input[1023]), .B(p_input[1007]), .Z(n8206) );
  XOR U8195 ( .A(n8383), .B(n8207), .Z(n8385) );
  AND U8196 ( .A(p_input[991]), .B(p_input[975]), .Z(n8207) );
  XOR U8197 ( .A(n8387), .B(n8388), .Z(n8383) );
  AND U8198 ( .A(n8389), .B(n8390), .Z(n8388) );
  XOR U8199 ( .A(n8387), .B(n8217), .Z(n8390) );
  XNOR U8200 ( .A(p_input[1006]), .B(n8391), .Z(n8217) );
  AND U8201 ( .A(n350), .B(n8392), .Z(n8391) );
  XOR U8202 ( .A(p_input[1022]), .B(p_input[1006]), .Z(n8392) );
  XNOR U8203 ( .A(n8214), .B(n8387), .Z(n8389) );
  XOR U8204 ( .A(n8393), .B(n8394), .Z(n8214) );
  AND U8205 ( .A(n348), .B(n8395), .Z(n8394) );
  XOR U8206 ( .A(p_input[990]), .B(p_input[974]), .Z(n8395) );
  XOR U8207 ( .A(n8396), .B(n8397), .Z(n8387) );
  AND U8208 ( .A(n8398), .B(n8399), .Z(n8397) );
  XOR U8209 ( .A(n8396), .B(n8229), .Z(n8399) );
  XNOR U8210 ( .A(p_input[1005]), .B(n8400), .Z(n8229) );
  AND U8211 ( .A(n350), .B(n8401), .Z(n8400) );
  XOR U8212 ( .A(p_input[1021]), .B(p_input[1005]), .Z(n8401) );
  XNOR U8213 ( .A(n8226), .B(n8396), .Z(n8398) );
  XOR U8214 ( .A(n8402), .B(n8403), .Z(n8226) );
  AND U8215 ( .A(n348), .B(n8404), .Z(n8403) );
  XOR U8216 ( .A(p_input[989]), .B(p_input[973]), .Z(n8404) );
  XOR U8217 ( .A(n8405), .B(n8406), .Z(n8396) );
  AND U8218 ( .A(n8407), .B(n8408), .Z(n8406) );
  XOR U8219 ( .A(n8405), .B(n8241), .Z(n8408) );
  XNOR U8220 ( .A(p_input[1004]), .B(n8409), .Z(n8241) );
  AND U8221 ( .A(n350), .B(n8410), .Z(n8409) );
  XOR U8222 ( .A(p_input[1020]), .B(p_input[1004]), .Z(n8410) );
  XNOR U8223 ( .A(n8238), .B(n8405), .Z(n8407) );
  XOR U8224 ( .A(n8411), .B(n8412), .Z(n8238) );
  AND U8225 ( .A(n348), .B(n8413), .Z(n8412) );
  XOR U8226 ( .A(p_input[988]), .B(p_input[972]), .Z(n8413) );
  XOR U8227 ( .A(n8414), .B(n8415), .Z(n8405) );
  AND U8228 ( .A(n8416), .B(n8417), .Z(n8415) );
  XOR U8229 ( .A(n8414), .B(n8253), .Z(n8417) );
  XNOR U8230 ( .A(p_input[1003]), .B(n8418), .Z(n8253) );
  AND U8231 ( .A(n350), .B(n8419), .Z(n8418) );
  XOR U8232 ( .A(p_input[1019]), .B(p_input[1003]), .Z(n8419) );
  XNOR U8233 ( .A(n8250), .B(n8414), .Z(n8416) );
  XOR U8234 ( .A(n8420), .B(n8421), .Z(n8250) );
  AND U8235 ( .A(n348), .B(n8422), .Z(n8421) );
  XOR U8236 ( .A(p_input[987]), .B(p_input[971]), .Z(n8422) );
  XOR U8237 ( .A(n8423), .B(n8424), .Z(n8414) );
  AND U8238 ( .A(n8425), .B(n8426), .Z(n8424) );
  XOR U8239 ( .A(n8423), .B(n8265), .Z(n8426) );
  XNOR U8240 ( .A(p_input[1002]), .B(n8427), .Z(n8265) );
  AND U8241 ( .A(n350), .B(n8428), .Z(n8427) );
  XOR U8242 ( .A(p_input[1018]), .B(p_input[1002]), .Z(n8428) );
  XNOR U8243 ( .A(n8262), .B(n8423), .Z(n8425) );
  XOR U8244 ( .A(n8429), .B(n8430), .Z(n8262) );
  AND U8245 ( .A(n348), .B(n8431), .Z(n8430) );
  XOR U8246 ( .A(p_input[986]), .B(p_input[970]), .Z(n8431) );
  XOR U8247 ( .A(n8432), .B(n8433), .Z(n8423) );
  AND U8248 ( .A(n8434), .B(n8435), .Z(n8433) );
  XOR U8249 ( .A(n8432), .B(n8277), .Z(n8435) );
  XNOR U8250 ( .A(p_input[1001]), .B(n8436), .Z(n8277) );
  AND U8251 ( .A(n350), .B(n8437), .Z(n8436) );
  XOR U8252 ( .A(p_input[1017]), .B(p_input[1001]), .Z(n8437) );
  XNOR U8253 ( .A(n8274), .B(n8432), .Z(n8434) );
  XOR U8254 ( .A(n8438), .B(n8439), .Z(n8274) );
  AND U8255 ( .A(n348), .B(n8440), .Z(n8439) );
  XOR U8256 ( .A(p_input[985]), .B(p_input[969]), .Z(n8440) );
  XOR U8257 ( .A(n8441), .B(n8442), .Z(n8432) );
  AND U8258 ( .A(n8443), .B(n8444), .Z(n8442) );
  XOR U8259 ( .A(n8441), .B(n8289), .Z(n8444) );
  XNOR U8260 ( .A(p_input[1000]), .B(n8445), .Z(n8289) );
  AND U8261 ( .A(n350), .B(n8446), .Z(n8445) );
  XOR U8262 ( .A(p_input[1016]), .B(p_input[1000]), .Z(n8446) );
  XNOR U8263 ( .A(n8286), .B(n8441), .Z(n8443) );
  XOR U8264 ( .A(n8447), .B(n8448), .Z(n8286) );
  AND U8265 ( .A(n348), .B(n8449), .Z(n8448) );
  XOR U8266 ( .A(p_input[984]), .B(p_input[968]), .Z(n8449) );
  XOR U8267 ( .A(n8450), .B(n8451), .Z(n8441) );
  AND U8268 ( .A(n8452), .B(n8453), .Z(n8451) );
  XOR U8269 ( .A(n8450), .B(n8301), .Z(n8453) );
  XNOR U8270 ( .A(p_input[999]), .B(n8454), .Z(n8301) );
  AND U8271 ( .A(n350), .B(n8455), .Z(n8454) );
  XOR U8272 ( .A(p_input[999]), .B(p_input[1015]), .Z(n8455) );
  XNOR U8273 ( .A(n8298), .B(n8450), .Z(n8452) );
  XOR U8274 ( .A(n8456), .B(n8457), .Z(n8298) );
  AND U8275 ( .A(n348), .B(n8458), .Z(n8457) );
  XOR U8276 ( .A(p_input[983]), .B(p_input[967]), .Z(n8458) );
  XOR U8277 ( .A(n8459), .B(n8460), .Z(n8450) );
  AND U8278 ( .A(n8461), .B(n8462), .Z(n8460) );
  XOR U8279 ( .A(n8459), .B(n8313), .Z(n8462) );
  XNOR U8280 ( .A(p_input[998]), .B(n8463), .Z(n8313) );
  AND U8281 ( .A(n350), .B(n8464), .Z(n8463) );
  XOR U8282 ( .A(p_input[998]), .B(p_input[1014]), .Z(n8464) );
  XNOR U8283 ( .A(n8310), .B(n8459), .Z(n8461) );
  XOR U8284 ( .A(n8465), .B(n8466), .Z(n8310) );
  AND U8285 ( .A(n348), .B(n8467), .Z(n8466) );
  XOR U8286 ( .A(p_input[982]), .B(p_input[966]), .Z(n8467) );
  XOR U8287 ( .A(n8468), .B(n8469), .Z(n8459) );
  AND U8288 ( .A(n8470), .B(n8471), .Z(n8469) );
  XOR U8289 ( .A(n8468), .B(n8325), .Z(n8471) );
  XNOR U8290 ( .A(p_input[997]), .B(n8472), .Z(n8325) );
  AND U8291 ( .A(n350), .B(n8473), .Z(n8472) );
  XOR U8292 ( .A(p_input[997]), .B(p_input[1013]), .Z(n8473) );
  XNOR U8293 ( .A(n8322), .B(n8468), .Z(n8470) );
  XOR U8294 ( .A(n8474), .B(n8475), .Z(n8322) );
  AND U8295 ( .A(n348), .B(n8476), .Z(n8475) );
  XOR U8296 ( .A(p_input[981]), .B(p_input[965]), .Z(n8476) );
  XOR U8297 ( .A(n8477), .B(n8478), .Z(n8468) );
  AND U8298 ( .A(n8479), .B(n8480), .Z(n8478) );
  XOR U8299 ( .A(n8477), .B(n8337), .Z(n8480) );
  XNOR U8300 ( .A(p_input[996]), .B(n8481), .Z(n8337) );
  AND U8301 ( .A(n350), .B(n8482), .Z(n8481) );
  XOR U8302 ( .A(p_input[996]), .B(p_input[1012]), .Z(n8482) );
  XNOR U8303 ( .A(n8334), .B(n8477), .Z(n8479) );
  XOR U8304 ( .A(n8483), .B(n8484), .Z(n8334) );
  AND U8305 ( .A(n348), .B(n8485), .Z(n8484) );
  XOR U8306 ( .A(p_input[980]), .B(p_input[964]), .Z(n8485) );
  XOR U8307 ( .A(n8486), .B(n8487), .Z(n8477) );
  AND U8308 ( .A(n8488), .B(n8489), .Z(n8487) );
  XOR U8309 ( .A(n8486), .B(n8349), .Z(n8489) );
  XNOR U8310 ( .A(p_input[995]), .B(n8490), .Z(n8349) );
  AND U8311 ( .A(n350), .B(n8491), .Z(n8490) );
  XOR U8312 ( .A(p_input[995]), .B(p_input[1011]), .Z(n8491) );
  XNOR U8313 ( .A(n8346), .B(n8486), .Z(n8488) );
  XOR U8314 ( .A(n8492), .B(n8493), .Z(n8346) );
  AND U8315 ( .A(n348), .B(n8494), .Z(n8493) );
  XOR U8316 ( .A(p_input[979]), .B(p_input[963]), .Z(n8494) );
  XOR U8317 ( .A(n8495), .B(n8496), .Z(n8486) );
  AND U8318 ( .A(n8497), .B(n8498), .Z(n8496) );
  XOR U8319 ( .A(n8361), .B(n8495), .Z(n8498) );
  XNOR U8320 ( .A(p_input[994]), .B(n8499), .Z(n8361) );
  AND U8321 ( .A(n350), .B(n8500), .Z(n8499) );
  XOR U8322 ( .A(p_input[994]), .B(p_input[1010]), .Z(n8500) );
  XNOR U8323 ( .A(n8495), .B(n8358), .Z(n8497) );
  XOR U8324 ( .A(n8501), .B(n8502), .Z(n8358) );
  AND U8325 ( .A(n348), .B(n8503), .Z(n8502) );
  XOR U8326 ( .A(p_input[978]), .B(p_input[962]), .Z(n8503) );
  XOR U8327 ( .A(n8504), .B(n8505), .Z(n8495) );
  AND U8328 ( .A(n8506), .B(n8507), .Z(n8505) );
  XNOR U8329 ( .A(n8508), .B(n8374), .Z(n8507) );
  XNOR U8330 ( .A(p_input[993]), .B(n8509), .Z(n8374) );
  AND U8331 ( .A(n350), .B(n8510), .Z(n8509) );
  XNOR U8332 ( .A(n8511), .B(p_input[1009]), .Z(n8510) );
  IV U8333 ( .A(p_input[993]), .Z(n8511) );
  XNOR U8334 ( .A(n8371), .B(n8504), .Z(n8506) );
  XNOR U8335 ( .A(p_input[961]), .B(n8512), .Z(n8371) );
  AND U8336 ( .A(n348), .B(n8513), .Z(n8512) );
  XOR U8337 ( .A(p_input[977]), .B(p_input[961]), .Z(n8513) );
  IV U8338 ( .A(n8508), .Z(n8504) );
  AND U8339 ( .A(n8379), .B(n8382), .Z(n8508) );
  XOR U8340 ( .A(p_input[992]), .B(n8514), .Z(n8382) );
  AND U8341 ( .A(n350), .B(n8515), .Z(n8514) );
  XOR U8342 ( .A(p_input[992]), .B(p_input[1008]), .Z(n8515) );
  XOR U8343 ( .A(n8516), .B(n8517), .Z(n350) );
  AND U8344 ( .A(n8518), .B(n8519), .Z(n8517) );
  XNOR U8345 ( .A(p_input[1023]), .B(n8516), .Z(n8519) );
  XOR U8346 ( .A(n8516), .B(p_input[1007]), .Z(n8518) );
  XOR U8347 ( .A(n8520), .B(n8521), .Z(n8516) );
  AND U8348 ( .A(n8522), .B(n8523), .Z(n8521) );
  XNOR U8349 ( .A(p_input[1022]), .B(n8520), .Z(n8523) );
  XOR U8350 ( .A(n8520), .B(p_input[1006]), .Z(n8522) );
  XOR U8351 ( .A(n8524), .B(n8525), .Z(n8520) );
  AND U8352 ( .A(n8526), .B(n8527), .Z(n8525) );
  XNOR U8353 ( .A(p_input[1021]), .B(n8524), .Z(n8527) );
  XOR U8354 ( .A(n8524), .B(p_input[1005]), .Z(n8526) );
  XOR U8355 ( .A(n8528), .B(n8529), .Z(n8524) );
  AND U8356 ( .A(n8530), .B(n8531), .Z(n8529) );
  XNOR U8357 ( .A(p_input[1020]), .B(n8528), .Z(n8531) );
  XOR U8358 ( .A(n8528), .B(p_input[1004]), .Z(n8530) );
  XOR U8359 ( .A(n8532), .B(n8533), .Z(n8528) );
  AND U8360 ( .A(n8534), .B(n8535), .Z(n8533) );
  XNOR U8361 ( .A(p_input[1019]), .B(n8532), .Z(n8535) );
  XOR U8362 ( .A(n8532), .B(p_input[1003]), .Z(n8534) );
  XOR U8363 ( .A(n8536), .B(n8537), .Z(n8532) );
  AND U8364 ( .A(n8538), .B(n8539), .Z(n8537) );
  XNOR U8365 ( .A(p_input[1018]), .B(n8536), .Z(n8539) );
  XOR U8366 ( .A(n8536), .B(p_input[1002]), .Z(n8538) );
  XOR U8367 ( .A(n8540), .B(n8541), .Z(n8536) );
  AND U8368 ( .A(n8542), .B(n8543), .Z(n8541) );
  XNOR U8369 ( .A(p_input[1017]), .B(n8540), .Z(n8543) );
  XOR U8370 ( .A(n8540), .B(p_input[1001]), .Z(n8542) );
  XOR U8371 ( .A(n8544), .B(n8545), .Z(n8540) );
  AND U8372 ( .A(n8546), .B(n8547), .Z(n8545) );
  XNOR U8373 ( .A(p_input[1016]), .B(n8544), .Z(n8547) );
  XOR U8374 ( .A(n8544), .B(p_input[1000]), .Z(n8546) );
  XOR U8375 ( .A(n8548), .B(n8549), .Z(n8544) );
  AND U8376 ( .A(n8550), .B(n8551), .Z(n8549) );
  XNOR U8377 ( .A(p_input[1015]), .B(n8548), .Z(n8551) );
  XOR U8378 ( .A(n8548), .B(p_input[999]), .Z(n8550) );
  XOR U8379 ( .A(n8552), .B(n8553), .Z(n8548) );
  AND U8380 ( .A(n8554), .B(n8555), .Z(n8553) );
  XNOR U8381 ( .A(p_input[1014]), .B(n8552), .Z(n8555) );
  XOR U8382 ( .A(n8552), .B(p_input[998]), .Z(n8554) );
  XOR U8383 ( .A(n8556), .B(n8557), .Z(n8552) );
  AND U8384 ( .A(n8558), .B(n8559), .Z(n8557) );
  XNOR U8385 ( .A(p_input[1013]), .B(n8556), .Z(n8559) );
  XOR U8386 ( .A(n8556), .B(p_input[997]), .Z(n8558) );
  XOR U8387 ( .A(n8560), .B(n8561), .Z(n8556) );
  AND U8388 ( .A(n8562), .B(n8563), .Z(n8561) );
  XNOR U8389 ( .A(p_input[1012]), .B(n8560), .Z(n8563) );
  XOR U8390 ( .A(n8560), .B(p_input[996]), .Z(n8562) );
  XOR U8391 ( .A(n8564), .B(n8565), .Z(n8560) );
  AND U8392 ( .A(n8566), .B(n8567), .Z(n8565) );
  XNOR U8393 ( .A(p_input[1011]), .B(n8564), .Z(n8567) );
  XOR U8394 ( .A(n8564), .B(p_input[995]), .Z(n8566) );
  XOR U8395 ( .A(n8568), .B(n8569), .Z(n8564) );
  AND U8396 ( .A(n8570), .B(n8571), .Z(n8569) );
  XNOR U8397 ( .A(p_input[1010]), .B(n8568), .Z(n8571) );
  XOR U8398 ( .A(n8568), .B(p_input[994]), .Z(n8570) );
  XNOR U8399 ( .A(n8572), .B(n8573), .Z(n8568) );
  AND U8400 ( .A(n8574), .B(n8575), .Z(n8573) );
  XOR U8401 ( .A(p_input[1009]), .B(n8572), .Z(n8575) );
  XNOR U8402 ( .A(p_input[993]), .B(n8572), .Z(n8574) );
  AND U8403 ( .A(p_input[1008]), .B(n8576), .Z(n8572) );
  IV U8404 ( .A(p_input[992]), .Z(n8576) );
  XNOR U8405 ( .A(p_input[960]), .B(n8577), .Z(n8379) );
  AND U8406 ( .A(n348), .B(n8578), .Z(n8577) );
  XOR U8407 ( .A(p_input[976]), .B(p_input[960]), .Z(n8578) );
  XOR U8408 ( .A(n8579), .B(n8580), .Z(n348) );
  AND U8409 ( .A(n8581), .B(n8582), .Z(n8580) );
  XNOR U8410 ( .A(p_input[991]), .B(n8579), .Z(n8582) );
  XOR U8411 ( .A(n8579), .B(p_input[975]), .Z(n8581) );
  XOR U8412 ( .A(n8583), .B(n8584), .Z(n8579) );
  AND U8413 ( .A(n8585), .B(n8586), .Z(n8584) );
  XNOR U8414 ( .A(p_input[990]), .B(n8583), .Z(n8586) );
  XNOR U8415 ( .A(n8583), .B(n8393), .Z(n8585) );
  IV U8416 ( .A(p_input[974]), .Z(n8393) );
  XOR U8417 ( .A(n8587), .B(n8588), .Z(n8583) );
  AND U8418 ( .A(n8589), .B(n8590), .Z(n8588) );
  XNOR U8419 ( .A(p_input[989]), .B(n8587), .Z(n8590) );
  XNOR U8420 ( .A(n8587), .B(n8402), .Z(n8589) );
  IV U8421 ( .A(p_input[973]), .Z(n8402) );
  XOR U8422 ( .A(n8591), .B(n8592), .Z(n8587) );
  AND U8423 ( .A(n8593), .B(n8594), .Z(n8592) );
  XNOR U8424 ( .A(p_input[988]), .B(n8591), .Z(n8594) );
  XNOR U8425 ( .A(n8591), .B(n8411), .Z(n8593) );
  IV U8426 ( .A(p_input[972]), .Z(n8411) );
  XOR U8427 ( .A(n8595), .B(n8596), .Z(n8591) );
  AND U8428 ( .A(n8597), .B(n8598), .Z(n8596) );
  XNOR U8429 ( .A(p_input[987]), .B(n8595), .Z(n8598) );
  XNOR U8430 ( .A(n8595), .B(n8420), .Z(n8597) );
  IV U8431 ( .A(p_input[971]), .Z(n8420) );
  XOR U8432 ( .A(n8599), .B(n8600), .Z(n8595) );
  AND U8433 ( .A(n8601), .B(n8602), .Z(n8600) );
  XNOR U8434 ( .A(p_input[986]), .B(n8599), .Z(n8602) );
  XNOR U8435 ( .A(n8599), .B(n8429), .Z(n8601) );
  IV U8436 ( .A(p_input[970]), .Z(n8429) );
  XOR U8437 ( .A(n8603), .B(n8604), .Z(n8599) );
  AND U8438 ( .A(n8605), .B(n8606), .Z(n8604) );
  XNOR U8439 ( .A(p_input[985]), .B(n8603), .Z(n8606) );
  XNOR U8440 ( .A(n8603), .B(n8438), .Z(n8605) );
  IV U8441 ( .A(p_input[969]), .Z(n8438) );
  XOR U8442 ( .A(n8607), .B(n8608), .Z(n8603) );
  AND U8443 ( .A(n8609), .B(n8610), .Z(n8608) );
  XNOR U8444 ( .A(p_input[984]), .B(n8607), .Z(n8610) );
  XNOR U8445 ( .A(n8607), .B(n8447), .Z(n8609) );
  IV U8446 ( .A(p_input[968]), .Z(n8447) );
  XOR U8447 ( .A(n8611), .B(n8612), .Z(n8607) );
  AND U8448 ( .A(n8613), .B(n8614), .Z(n8612) );
  XNOR U8449 ( .A(p_input[983]), .B(n8611), .Z(n8614) );
  XNOR U8450 ( .A(n8611), .B(n8456), .Z(n8613) );
  IV U8451 ( .A(p_input[967]), .Z(n8456) );
  XOR U8452 ( .A(n8615), .B(n8616), .Z(n8611) );
  AND U8453 ( .A(n8617), .B(n8618), .Z(n8616) );
  XNOR U8454 ( .A(p_input[982]), .B(n8615), .Z(n8618) );
  XNOR U8455 ( .A(n8615), .B(n8465), .Z(n8617) );
  IV U8456 ( .A(p_input[966]), .Z(n8465) );
  XOR U8457 ( .A(n8619), .B(n8620), .Z(n8615) );
  AND U8458 ( .A(n8621), .B(n8622), .Z(n8620) );
  XNOR U8459 ( .A(p_input[981]), .B(n8619), .Z(n8622) );
  XNOR U8460 ( .A(n8619), .B(n8474), .Z(n8621) );
  IV U8461 ( .A(p_input[965]), .Z(n8474) );
  XOR U8462 ( .A(n8623), .B(n8624), .Z(n8619) );
  AND U8463 ( .A(n8625), .B(n8626), .Z(n8624) );
  XNOR U8464 ( .A(p_input[980]), .B(n8623), .Z(n8626) );
  XNOR U8465 ( .A(n8623), .B(n8483), .Z(n8625) );
  IV U8466 ( .A(p_input[964]), .Z(n8483) );
  XOR U8467 ( .A(n8627), .B(n8628), .Z(n8623) );
  AND U8468 ( .A(n8629), .B(n8630), .Z(n8628) );
  XNOR U8469 ( .A(p_input[979]), .B(n8627), .Z(n8630) );
  XNOR U8470 ( .A(n8627), .B(n8492), .Z(n8629) );
  IV U8471 ( .A(p_input[963]), .Z(n8492) );
  XOR U8472 ( .A(n8631), .B(n8632), .Z(n8627) );
  AND U8473 ( .A(n8633), .B(n8634), .Z(n8632) );
  XNOR U8474 ( .A(p_input[978]), .B(n8631), .Z(n8634) );
  XNOR U8475 ( .A(n8631), .B(n8501), .Z(n8633) );
  IV U8476 ( .A(p_input[962]), .Z(n8501) );
  XNOR U8477 ( .A(n8635), .B(n8636), .Z(n8631) );
  AND U8478 ( .A(n8637), .B(n8638), .Z(n8636) );
  XOR U8479 ( .A(p_input[977]), .B(n8635), .Z(n8638) );
  XNOR U8480 ( .A(p_input[961]), .B(n8635), .Z(n8637) );
  AND U8481 ( .A(p_input[976]), .B(n8639), .Z(n8635) );
  IV U8482 ( .A(p_input[960]), .Z(n8639) );
  XOR U8483 ( .A(n8640), .B(n8641), .Z(n8198) );
  AND U8484 ( .A(n284), .B(n8642), .Z(n8641) );
  XNOR U8485 ( .A(n8643), .B(n8640), .Z(n8642) );
  XOR U8486 ( .A(n8644), .B(n8645), .Z(n284) );
  AND U8487 ( .A(n8646), .B(n8647), .Z(n8645) );
  XNOR U8488 ( .A(n8208), .B(n8644), .Z(n8647) );
  AND U8489 ( .A(p_input[959]), .B(p_input[943]), .Z(n8208) );
  XOR U8490 ( .A(n8644), .B(n8209), .Z(n8646) );
  AND U8491 ( .A(p_input[927]), .B(p_input[911]), .Z(n8209) );
  XOR U8492 ( .A(n8648), .B(n8649), .Z(n8644) );
  AND U8493 ( .A(n8650), .B(n8651), .Z(n8649) );
  XOR U8494 ( .A(n8648), .B(n8221), .Z(n8651) );
  XNOR U8495 ( .A(p_input[942]), .B(n8652), .Z(n8221) );
  AND U8496 ( .A(n354), .B(n8653), .Z(n8652) );
  XOR U8497 ( .A(p_input[958]), .B(p_input[942]), .Z(n8653) );
  XNOR U8498 ( .A(n8218), .B(n8648), .Z(n8650) );
  XOR U8499 ( .A(n8654), .B(n8655), .Z(n8218) );
  AND U8500 ( .A(n351), .B(n8656), .Z(n8655) );
  XOR U8501 ( .A(p_input[926]), .B(p_input[910]), .Z(n8656) );
  XOR U8502 ( .A(n8657), .B(n8658), .Z(n8648) );
  AND U8503 ( .A(n8659), .B(n8660), .Z(n8658) );
  XOR U8504 ( .A(n8657), .B(n8233), .Z(n8660) );
  XNOR U8505 ( .A(p_input[941]), .B(n8661), .Z(n8233) );
  AND U8506 ( .A(n354), .B(n8662), .Z(n8661) );
  XOR U8507 ( .A(p_input[957]), .B(p_input[941]), .Z(n8662) );
  XNOR U8508 ( .A(n8230), .B(n8657), .Z(n8659) );
  XOR U8509 ( .A(n8663), .B(n8664), .Z(n8230) );
  AND U8510 ( .A(n351), .B(n8665), .Z(n8664) );
  XOR U8511 ( .A(p_input[925]), .B(p_input[909]), .Z(n8665) );
  XOR U8512 ( .A(n8666), .B(n8667), .Z(n8657) );
  AND U8513 ( .A(n8668), .B(n8669), .Z(n8667) );
  XOR U8514 ( .A(n8666), .B(n8245), .Z(n8669) );
  XNOR U8515 ( .A(p_input[940]), .B(n8670), .Z(n8245) );
  AND U8516 ( .A(n354), .B(n8671), .Z(n8670) );
  XOR U8517 ( .A(p_input[956]), .B(p_input[940]), .Z(n8671) );
  XNOR U8518 ( .A(n8242), .B(n8666), .Z(n8668) );
  XOR U8519 ( .A(n8672), .B(n8673), .Z(n8242) );
  AND U8520 ( .A(n351), .B(n8674), .Z(n8673) );
  XOR U8521 ( .A(p_input[924]), .B(p_input[908]), .Z(n8674) );
  XOR U8522 ( .A(n8675), .B(n8676), .Z(n8666) );
  AND U8523 ( .A(n8677), .B(n8678), .Z(n8676) );
  XOR U8524 ( .A(n8675), .B(n8257), .Z(n8678) );
  XNOR U8525 ( .A(p_input[939]), .B(n8679), .Z(n8257) );
  AND U8526 ( .A(n354), .B(n8680), .Z(n8679) );
  XOR U8527 ( .A(p_input[955]), .B(p_input[939]), .Z(n8680) );
  XNOR U8528 ( .A(n8254), .B(n8675), .Z(n8677) );
  XOR U8529 ( .A(n8681), .B(n8682), .Z(n8254) );
  AND U8530 ( .A(n351), .B(n8683), .Z(n8682) );
  XOR U8531 ( .A(p_input[923]), .B(p_input[907]), .Z(n8683) );
  XOR U8532 ( .A(n8684), .B(n8685), .Z(n8675) );
  AND U8533 ( .A(n8686), .B(n8687), .Z(n8685) );
  XOR U8534 ( .A(n8684), .B(n8269), .Z(n8687) );
  XNOR U8535 ( .A(p_input[938]), .B(n8688), .Z(n8269) );
  AND U8536 ( .A(n354), .B(n8689), .Z(n8688) );
  XOR U8537 ( .A(p_input[954]), .B(p_input[938]), .Z(n8689) );
  XNOR U8538 ( .A(n8266), .B(n8684), .Z(n8686) );
  XOR U8539 ( .A(n8690), .B(n8691), .Z(n8266) );
  AND U8540 ( .A(n351), .B(n8692), .Z(n8691) );
  XOR U8541 ( .A(p_input[922]), .B(p_input[906]), .Z(n8692) );
  XOR U8542 ( .A(n8693), .B(n8694), .Z(n8684) );
  AND U8543 ( .A(n8695), .B(n8696), .Z(n8694) );
  XOR U8544 ( .A(n8693), .B(n8281), .Z(n8696) );
  XNOR U8545 ( .A(p_input[937]), .B(n8697), .Z(n8281) );
  AND U8546 ( .A(n354), .B(n8698), .Z(n8697) );
  XOR U8547 ( .A(p_input[953]), .B(p_input[937]), .Z(n8698) );
  XNOR U8548 ( .A(n8278), .B(n8693), .Z(n8695) );
  XOR U8549 ( .A(n8699), .B(n8700), .Z(n8278) );
  AND U8550 ( .A(n351), .B(n8701), .Z(n8700) );
  XOR U8551 ( .A(p_input[921]), .B(p_input[905]), .Z(n8701) );
  XOR U8552 ( .A(n8702), .B(n8703), .Z(n8693) );
  AND U8553 ( .A(n8704), .B(n8705), .Z(n8703) );
  XOR U8554 ( .A(n8702), .B(n8293), .Z(n8705) );
  XNOR U8555 ( .A(p_input[936]), .B(n8706), .Z(n8293) );
  AND U8556 ( .A(n354), .B(n8707), .Z(n8706) );
  XOR U8557 ( .A(p_input[952]), .B(p_input[936]), .Z(n8707) );
  XNOR U8558 ( .A(n8290), .B(n8702), .Z(n8704) );
  XOR U8559 ( .A(n8708), .B(n8709), .Z(n8290) );
  AND U8560 ( .A(n351), .B(n8710), .Z(n8709) );
  XOR U8561 ( .A(p_input[920]), .B(p_input[904]), .Z(n8710) );
  XOR U8562 ( .A(n8711), .B(n8712), .Z(n8702) );
  AND U8563 ( .A(n8713), .B(n8714), .Z(n8712) );
  XOR U8564 ( .A(n8711), .B(n8305), .Z(n8714) );
  XNOR U8565 ( .A(p_input[935]), .B(n8715), .Z(n8305) );
  AND U8566 ( .A(n354), .B(n8716), .Z(n8715) );
  XOR U8567 ( .A(p_input[951]), .B(p_input[935]), .Z(n8716) );
  XNOR U8568 ( .A(n8302), .B(n8711), .Z(n8713) );
  XOR U8569 ( .A(n8717), .B(n8718), .Z(n8302) );
  AND U8570 ( .A(n351), .B(n8719), .Z(n8718) );
  XOR U8571 ( .A(p_input[919]), .B(p_input[903]), .Z(n8719) );
  XOR U8572 ( .A(n8720), .B(n8721), .Z(n8711) );
  AND U8573 ( .A(n8722), .B(n8723), .Z(n8721) );
  XOR U8574 ( .A(n8720), .B(n8317), .Z(n8723) );
  XNOR U8575 ( .A(p_input[934]), .B(n8724), .Z(n8317) );
  AND U8576 ( .A(n354), .B(n8725), .Z(n8724) );
  XOR U8577 ( .A(p_input[950]), .B(p_input[934]), .Z(n8725) );
  XNOR U8578 ( .A(n8314), .B(n8720), .Z(n8722) );
  XOR U8579 ( .A(n8726), .B(n8727), .Z(n8314) );
  AND U8580 ( .A(n351), .B(n8728), .Z(n8727) );
  XOR U8581 ( .A(p_input[918]), .B(p_input[902]), .Z(n8728) );
  XOR U8582 ( .A(n8729), .B(n8730), .Z(n8720) );
  AND U8583 ( .A(n8731), .B(n8732), .Z(n8730) );
  XOR U8584 ( .A(n8729), .B(n8329), .Z(n8732) );
  XNOR U8585 ( .A(p_input[933]), .B(n8733), .Z(n8329) );
  AND U8586 ( .A(n354), .B(n8734), .Z(n8733) );
  XOR U8587 ( .A(p_input[949]), .B(p_input[933]), .Z(n8734) );
  XNOR U8588 ( .A(n8326), .B(n8729), .Z(n8731) );
  XOR U8589 ( .A(n8735), .B(n8736), .Z(n8326) );
  AND U8590 ( .A(n351), .B(n8737), .Z(n8736) );
  XOR U8591 ( .A(p_input[917]), .B(p_input[901]), .Z(n8737) );
  XOR U8592 ( .A(n8738), .B(n8739), .Z(n8729) );
  AND U8593 ( .A(n8740), .B(n8741), .Z(n8739) );
  XOR U8594 ( .A(n8738), .B(n8341), .Z(n8741) );
  XNOR U8595 ( .A(p_input[932]), .B(n8742), .Z(n8341) );
  AND U8596 ( .A(n354), .B(n8743), .Z(n8742) );
  XOR U8597 ( .A(p_input[948]), .B(p_input[932]), .Z(n8743) );
  XNOR U8598 ( .A(n8338), .B(n8738), .Z(n8740) );
  XOR U8599 ( .A(n8744), .B(n8745), .Z(n8338) );
  AND U8600 ( .A(n351), .B(n8746), .Z(n8745) );
  XOR U8601 ( .A(p_input[916]), .B(p_input[900]), .Z(n8746) );
  XOR U8602 ( .A(n8747), .B(n8748), .Z(n8738) );
  AND U8603 ( .A(n8749), .B(n8750), .Z(n8748) );
  XOR U8604 ( .A(n8747), .B(n8353), .Z(n8750) );
  XNOR U8605 ( .A(p_input[931]), .B(n8751), .Z(n8353) );
  AND U8606 ( .A(n354), .B(n8752), .Z(n8751) );
  XOR U8607 ( .A(p_input[947]), .B(p_input[931]), .Z(n8752) );
  XNOR U8608 ( .A(n8350), .B(n8747), .Z(n8749) );
  XOR U8609 ( .A(n8753), .B(n8754), .Z(n8350) );
  AND U8610 ( .A(n351), .B(n8755), .Z(n8754) );
  XOR U8611 ( .A(p_input[915]), .B(p_input[899]), .Z(n8755) );
  XOR U8612 ( .A(n8756), .B(n8757), .Z(n8747) );
  AND U8613 ( .A(n8758), .B(n8759), .Z(n8757) );
  XOR U8614 ( .A(n8365), .B(n8756), .Z(n8759) );
  XNOR U8615 ( .A(p_input[930]), .B(n8760), .Z(n8365) );
  AND U8616 ( .A(n354), .B(n8761), .Z(n8760) );
  XOR U8617 ( .A(p_input[946]), .B(p_input[930]), .Z(n8761) );
  XNOR U8618 ( .A(n8756), .B(n8362), .Z(n8758) );
  XOR U8619 ( .A(n8762), .B(n8763), .Z(n8362) );
  AND U8620 ( .A(n351), .B(n8764), .Z(n8763) );
  XOR U8621 ( .A(p_input[914]), .B(p_input[898]), .Z(n8764) );
  XOR U8622 ( .A(n8765), .B(n8766), .Z(n8756) );
  AND U8623 ( .A(n8767), .B(n8768), .Z(n8766) );
  XNOR U8624 ( .A(n8769), .B(n8378), .Z(n8768) );
  XNOR U8625 ( .A(p_input[929]), .B(n8770), .Z(n8378) );
  AND U8626 ( .A(n354), .B(n8771), .Z(n8770) );
  XNOR U8627 ( .A(p_input[945]), .B(n8772), .Z(n8771) );
  IV U8628 ( .A(p_input[929]), .Z(n8772) );
  XNOR U8629 ( .A(n8375), .B(n8765), .Z(n8767) );
  XNOR U8630 ( .A(p_input[897]), .B(n8773), .Z(n8375) );
  AND U8631 ( .A(n351), .B(n8774), .Z(n8773) );
  XOR U8632 ( .A(p_input[913]), .B(p_input[897]), .Z(n8774) );
  IV U8633 ( .A(n8769), .Z(n8765) );
  AND U8634 ( .A(n8640), .B(n8643), .Z(n8769) );
  XOR U8635 ( .A(p_input[928]), .B(n8775), .Z(n8643) );
  AND U8636 ( .A(n354), .B(n8776), .Z(n8775) );
  XOR U8637 ( .A(p_input[944]), .B(p_input[928]), .Z(n8776) );
  XOR U8638 ( .A(n8777), .B(n8778), .Z(n354) );
  AND U8639 ( .A(n8779), .B(n8780), .Z(n8778) );
  XNOR U8640 ( .A(p_input[959]), .B(n8777), .Z(n8780) );
  XOR U8641 ( .A(n8777), .B(p_input[943]), .Z(n8779) );
  XOR U8642 ( .A(n8781), .B(n8782), .Z(n8777) );
  AND U8643 ( .A(n8783), .B(n8784), .Z(n8782) );
  XNOR U8644 ( .A(p_input[958]), .B(n8781), .Z(n8784) );
  XOR U8645 ( .A(n8781), .B(p_input[942]), .Z(n8783) );
  XOR U8646 ( .A(n8785), .B(n8786), .Z(n8781) );
  AND U8647 ( .A(n8787), .B(n8788), .Z(n8786) );
  XNOR U8648 ( .A(p_input[957]), .B(n8785), .Z(n8788) );
  XOR U8649 ( .A(n8785), .B(p_input[941]), .Z(n8787) );
  XOR U8650 ( .A(n8789), .B(n8790), .Z(n8785) );
  AND U8651 ( .A(n8791), .B(n8792), .Z(n8790) );
  XNOR U8652 ( .A(p_input[956]), .B(n8789), .Z(n8792) );
  XOR U8653 ( .A(n8789), .B(p_input[940]), .Z(n8791) );
  XOR U8654 ( .A(n8793), .B(n8794), .Z(n8789) );
  AND U8655 ( .A(n8795), .B(n8796), .Z(n8794) );
  XNOR U8656 ( .A(p_input[955]), .B(n8793), .Z(n8796) );
  XOR U8657 ( .A(n8793), .B(p_input[939]), .Z(n8795) );
  XOR U8658 ( .A(n8797), .B(n8798), .Z(n8793) );
  AND U8659 ( .A(n8799), .B(n8800), .Z(n8798) );
  XNOR U8660 ( .A(p_input[954]), .B(n8797), .Z(n8800) );
  XOR U8661 ( .A(n8797), .B(p_input[938]), .Z(n8799) );
  XOR U8662 ( .A(n8801), .B(n8802), .Z(n8797) );
  AND U8663 ( .A(n8803), .B(n8804), .Z(n8802) );
  XNOR U8664 ( .A(p_input[953]), .B(n8801), .Z(n8804) );
  XOR U8665 ( .A(n8801), .B(p_input[937]), .Z(n8803) );
  XOR U8666 ( .A(n8805), .B(n8806), .Z(n8801) );
  AND U8667 ( .A(n8807), .B(n8808), .Z(n8806) );
  XNOR U8668 ( .A(p_input[952]), .B(n8805), .Z(n8808) );
  XOR U8669 ( .A(n8805), .B(p_input[936]), .Z(n8807) );
  XOR U8670 ( .A(n8809), .B(n8810), .Z(n8805) );
  AND U8671 ( .A(n8811), .B(n8812), .Z(n8810) );
  XNOR U8672 ( .A(p_input[951]), .B(n8809), .Z(n8812) );
  XOR U8673 ( .A(n8809), .B(p_input[935]), .Z(n8811) );
  XOR U8674 ( .A(n8813), .B(n8814), .Z(n8809) );
  AND U8675 ( .A(n8815), .B(n8816), .Z(n8814) );
  XNOR U8676 ( .A(p_input[950]), .B(n8813), .Z(n8816) );
  XOR U8677 ( .A(n8813), .B(p_input[934]), .Z(n8815) );
  XOR U8678 ( .A(n8817), .B(n8818), .Z(n8813) );
  AND U8679 ( .A(n8819), .B(n8820), .Z(n8818) );
  XNOR U8680 ( .A(p_input[949]), .B(n8817), .Z(n8820) );
  XOR U8681 ( .A(n8817), .B(p_input[933]), .Z(n8819) );
  XOR U8682 ( .A(n8821), .B(n8822), .Z(n8817) );
  AND U8683 ( .A(n8823), .B(n8824), .Z(n8822) );
  XNOR U8684 ( .A(p_input[948]), .B(n8821), .Z(n8824) );
  XOR U8685 ( .A(n8821), .B(p_input[932]), .Z(n8823) );
  XOR U8686 ( .A(n8825), .B(n8826), .Z(n8821) );
  AND U8687 ( .A(n8827), .B(n8828), .Z(n8826) );
  XNOR U8688 ( .A(p_input[947]), .B(n8825), .Z(n8828) );
  XOR U8689 ( .A(n8825), .B(p_input[931]), .Z(n8827) );
  XOR U8690 ( .A(n8829), .B(n8830), .Z(n8825) );
  AND U8691 ( .A(n8831), .B(n8832), .Z(n8830) );
  XNOR U8692 ( .A(p_input[946]), .B(n8829), .Z(n8832) );
  XOR U8693 ( .A(n8829), .B(p_input[930]), .Z(n8831) );
  XNOR U8694 ( .A(n8833), .B(n8834), .Z(n8829) );
  AND U8695 ( .A(n8835), .B(n8836), .Z(n8834) );
  XOR U8696 ( .A(p_input[945]), .B(n8833), .Z(n8836) );
  XNOR U8697 ( .A(p_input[929]), .B(n8833), .Z(n8835) );
  AND U8698 ( .A(p_input[944]), .B(n8837), .Z(n8833) );
  IV U8699 ( .A(p_input[928]), .Z(n8837) );
  XNOR U8700 ( .A(p_input[896]), .B(n8838), .Z(n8640) );
  AND U8701 ( .A(n351), .B(n8839), .Z(n8838) );
  XOR U8702 ( .A(p_input[912]), .B(p_input[896]), .Z(n8839) );
  XOR U8703 ( .A(n8840), .B(n8841), .Z(n351) );
  AND U8704 ( .A(n8842), .B(n8843), .Z(n8841) );
  XNOR U8705 ( .A(p_input[927]), .B(n8840), .Z(n8843) );
  XOR U8706 ( .A(n8840), .B(p_input[911]), .Z(n8842) );
  XOR U8707 ( .A(n8844), .B(n8845), .Z(n8840) );
  AND U8708 ( .A(n8846), .B(n8847), .Z(n8845) );
  XNOR U8709 ( .A(p_input[926]), .B(n8844), .Z(n8847) );
  XNOR U8710 ( .A(n8844), .B(n8654), .Z(n8846) );
  IV U8711 ( .A(p_input[910]), .Z(n8654) );
  XOR U8712 ( .A(n8848), .B(n8849), .Z(n8844) );
  AND U8713 ( .A(n8850), .B(n8851), .Z(n8849) );
  XNOR U8714 ( .A(p_input[925]), .B(n8848), .Z(n8851) );
  XNOR U8715 ( .A(n8848), .B(n8663), .Z(n8850) );
  IV U8716 ( .A(p_input[909]), .Z(n8663) );
  XOR U8717 ( .A(n8852), .B(n8853), .Z(n8848) );
  AND U8718 ( .A(n8854), .B(n8855), .Z(n8853) );
  XNOR U8719 ( .A(p_input[924]), .B(n8852), .Z(n8855) );
  XNOR U8720 ( .A(n8852), .B(n8672), .Z(n8854) );
  IV U8721 ( .A(p_input[908]), .Z(n8672) );
  XOR U8722 ( .A(n8856), .B(n8857), .Z(n8852) );
  AND U8723 ( .A(n8858), .B(n8859), .Z(n8857) );
  XNOR U8724 ( .A(p_input[923]), .B(n8856), .Z(n8859) );
  XNOR U8725 ( .A(n8856), .B(n8681), .Z(n8858) );
  IV U8726 ( .A(p_input[907]), .Z(n8681) );
  XOR U8727 ( .A(n8860), .B(n8861), .Z(n8856) );
  AND U8728 ( .A(n8862), .B(n8863), .Z(n8861) );
  XNOR U8729 ( .A(p_input[922]), .B(n8860), .Z(n8863) );
  XNOR U8730 ( .A(n8860), .B(n8690), .Z(n8862) );
  IV U8731 ( .A(p_input[906]), .Z(n8690) );
  XOR U8732 ( .A(n8864), .B(n8865), .Z(n8860) );
  AND U8733 ( .A(n8866), .B(n8867), .Z(n8865) );
  XNOR U8734 ( .A(p_input[921]), .B(n8864), .Z(n8867) );
  XNOR U8735 ( .A(n8864), .B(n8699), .Z(n8866) );
  IV U8736 ( .A(p_input[905]), .Z(n8699) );
  XOR U8737 ( .A(n8868), .B(n8869), .Z(n8864) );
  AND U8738 ( .A(n8870), .B(n8871), .Z(n8869) );
  XNOR U8739 ( .A(p_input[920]), .B(n8868), .Z(n8871) );
  XNOR U8740 ( .A(n8868), .B(n8708), .Z(n8870) );
  IV U8741 ( .A(p_input[904]), .Z(n8708) );
  XOR U8742 ( .A(n8872), .B(n8873), .Z(n8868) );
  AND U8743 ( .A(n8874), .B(n8875), .Z(n8873) );
  XNOR U8744 ( .A(p_input[919]), .B(n8872), .Z(n8875) );
  XNOR U8745 ( .A(n8872), .B(n8717), .Z(n8874) );
  IV U8746 ( .A(p_input[903]), .Z(n8717) );
  XOR U8747 ( .A(n8876), .B(n8877), .Z(n8872) );
  AND U8748 ( .A(n8878), .B(n8879), .Z(n8877) );
  XNOR U8749 ( .A(p_input[918]), .B(n8876), .Z(n8879) );
  XNOR U8750 ( .A(n8876), .B(n8726), .Z(n8878) );
  IV U8751 ( .A(p_input[902]), .Z(n8726) );
  XOR U8752 ( .A(n8880), .B(n8881), .Z(n8876) );
  AND U8753 ( .A(n8882), .B(n8883), .Z(n8881) );
  XNOR U8754 ( .A(p_input[917]), .B(n8880), .Z(n8883) );
  XNOR U8755 ( .A(n8880), .B(n8735), .Z(n8882) );
  IV U8756 ( .A(p_input[901]), .Z(n8735) );
  XOR U8757 ( .A(n8884), .B(n8885), .Z(n8880) );
  AND U8758 ( .A(n8886), .B(n8887), .Z(n8885) );
  XNOR U8759 ( .A(p_input[916]), .B(n8884), .Z(n8887) );
  XNOR U8760 ( .A(n8884), .B(n8744), .Z(n8886) );
  IV U8761 ( .A(p_input[900]), .Z(n8744) );
  XOR U8762 ( .A(n8888), .B(n8889), .Z(n8884) );
  AND U8763 ( .A(n8890), .B(n8891), .Z(n8889) );
  XNOR U8764 ( .A(p_input[915]), .B(n8888), .Z(n8891) );
  XNOR U8765 ( .A(n8888), .B(n8753), .Z(n8890) );
  IV U8766 ( .A(p_input[899]), .Z(n8753) );
  XOR U8767 ( .A(n8892), .B(n8893), .Z(n8888) );
  AND U8768 ( .A(n8894), .B(n8895), .Z(n8893) );
  XNOR U8769 ( .A(p_input[914]), .B(n8892), .Z(n8895) );
  XNOR U8770 ( .A(n8892), .B(n8762), .Z(n8894) );
  IV U8771 ( .A(p_input[898]), .Z(n8762) );
  XNOR U8772 ( .A(n8896), .B(n8897), .Z(n8892) );
  AND U8773 ( .A(n8898), .B(n8899), .Z(n8897) );
  XOR U8774 ( .A(p_input[913]), .B(n8896), .Z(n8899) );
  XNOR U8775 ( .A(p_input[897]), .B(n8896), .Z(n8898) );
  AND U8776 ( .A(p_input[912]), .B(n8900), .Z(n8896) );
  IV U8777 ( .A(p_input[896]), .Z(n8900) );
  XOR U8778 ( .A(n8901), .B(n8902), .Z(n8016) );
  AND U8779 ( .A(n436), .B(n8903), .Z(n8902) );
  XNOR U8780 ( .A(n8904), .B(n8901), .Z(n8903) );
  XOR U8781 ( .A(n8905), .B(n8906), .Z(n436) );
  AND U8782 ( .A(n8907), .B(n8908), .Z(n8906) );
  XNOR U8783 ( .A(n8028), .B(n8905), .Z(n8908) );
  AND U8784 ( .A(n8909), .B(n8910), .Z(n8028) );
  XOR U8785 ( .A(n8905), .B(n8027), .Z(n8907) );
  AND U8786 ( .A(n8911), .B(n8912), .Z(n8027) );
  XOR U8787 ( .A(n8913), .B(n8914), .Z(n8905) );
  AND U8788 ( .A(n8915), .B(n8916), .Z(n8914) );
  XOR U8789 ( .A(n8913), .B(n8040), .Z(n8916) );
  XOR U8790 ( .A(n8917), .B(n8918), .Z(n8040) );
  AND U8791 ( .A(n290), .B(n8919), .Z(n8918) );
  XOR U8792 ( .A(n8920), .B(n8917), .Z(n8919) );
  XNOR U8793 ( .A(n8037), .B(n8913), .Z(n8915) );
  XOR U8794 ( .A(n8921), .B(n8922), .Z(n8037) );
  AND U8795 ( .A(n287), .B(n8923), .Z(n8922) );
  XOR U8796 ( .A(n8924), .B(n8921), .Z(n8923) );
  XOR U8797 ( .A(n8925), .B(n8926), .Z(n8913) );
  AND U8798 ( .A(n8927), .B(n8928), .Z(n8926) );
  XOR U8799 ( .A(n8925), .B(n8052), .Z(n8928) );
  XOR U8800 ( .A(n8929), .B(n8930), .Z(n8052) );
  AND U8801 ( .A(n290), .B(n8931), .Z(n8930) );
  XOR U8802 ( .A(n8932), .B(n8929), .Z(n8931) );
  XNOR U8803 ( .A(n8049), .B(n8925), .Z(n8927) );
  XOR U8804 ( .A(n8933), .B(n8934), .Z(n8049) );
  AND U8805 ( .A(n287), .B(n8935), .Z(n8934) );
  XOR U8806 ( .A(n8936), .B(n8933), .Z(n8935) );
  XOR U8807 ( .A(n8937), .B(n8938), .Z(n8925) );
  AND U8808 ( .A(n8939), .B(n8940), .Z(n8938) );
  XOR U8809 ( .A(n8937), .B(n8064), .Z(n8940) );
  XOR U8810 ( .A(n8941), .B(n8942), .Z(n8064) );
  AND U8811 ( .A(n290), .B(n8943), .Z(n8942) );
  XOR U8812 ( .A(n8944), .B(n8941), .Z(n8943) );
  XNOR U8813 ( .A(n8061), .B(n8937), .Z(n8939) );
  XOR U8814 ( .A(n8945), .B(n8946), .Z(n8061) );
  AND U8815 ( .A(n287), .B(n8947), .Z(n8946) );
  XOR U8816 ( .A(n8948), .B(n8945), .Z(n8947) );
  XOR U8817 ( .A(n8949), .B(n8950), .Z(n8937) );
  AND U8818 ( .A(n8951), .B(n8952), .Z(n8950) );
  XOR U8819 ( .A(n8949), .B(n8076), .Z(n8952) );
  XOR U8820 ( .A(n8953), .B(n8954), .Z(n8076) );
  AND U8821 ( .A(n290), .B(n8955), .Z(n8954) );
  XOR U8822 ( .A(n8956), .B(n8953), .Z(n8955) );
  XNOR U8823 ( .A(n8073), .B(n8949), .Z(n8951) );
  XOR U8824 ( .A(n8957), .B(n8958), .Z(n8073) );
  AND U8825 ( .A(n287), .B(n8959), .Z(n8958) );
  XOR U8826 ( .A(n8960), .B(n8957), .Z(n8959) );
  XOR U8827 ( .A(n8961), .B(n8962), .Z(n8949) );
  AND U8828 ( .A(n8963), .B(n8964), .Z(n8962) );
  XOR U8829 ( .A(n8961), .B(n8088), .Z(n8964) );
  XOR U8830 ( .A(n8965), .B(n8966), .Z(n8088) );
  AND U8831 ( .A(n290), .B(n8967), .Z(n8966) );
  XOR U8832 ( .A(n8968), .B(n8965), .Z(n8967) );
  XNOR U8833 ( .A(n8085), .B(n8961), .Z(n8963) );
  XOR U8834 ( .A(n8969), .B(n8970), .Z(n8085) );
  AND U8835 ( .A(n287), .B(n8971), .Z(n8970) );
  XOR U8836 ( .A(n8972), .B(n8969), .Z(n8971) );
  XOR U8837 ( .A(n8973), .B(n8974), .Z(n8961) );
  AND U8838 ( .A(n8975), .B(n8976), .Z(n8974) );
  XOR U8839 ( .A(n8973), .B(n8100), .Z(n8976) );
  XOR U8840 ( .A(n8977), .B(n8978), .Z(n8100) );
  AND U8841 ( .A(n290), .B(n8979), .Z(n8978) );
  XOR U8842 ( .A(n8980), .B(n8977), .Z(n8979) );
  XNOR U8843 ( .A(n8097), .B(n8973), .Z(n8975) );
  XOR U8844 ( .A(n8981), .B(n8982), .Z(n8097) );
  AND U8845 ( .A(n287), .B(n8983), .Z(n8982) );
  XOR U8846 ( .A(n8984), .B(n8981), .Z(n8983) );
  XOR U8847 ( .A(n8985), .B(n8986), .Z(n8973) );
  AND U8848 ( .A(n8987), .B(n8988), .Z(n8986) );
  XOR U8849 ( .A(n8985), .B(n8112), .Z(n8988) );
  XOR U8850 ( .A(n8989), .B(n8990), .Z(n8112) );
  AND U8851 ( .A(n290), .B(n8991), .Z(n8990) );
  XOR U8852 ( .A(n8992), .B(n8989), .Z(n8991) );
  XNOR U8853 ( .A(n8109), .B(n8985), .Z(n8987) );
  XOR U8854 ( .A(n8993), .B(n8994), .Z(n8109) );
  AND U8855 ( .A(n287), .B(n8995), .Z(n8994) );
  XOR U8856 ( .A(n8996), .B(n8993), .Z(n8995) );
  XOR U8857 ( .A(n8997), .B(n8998), .Z(n8985) );
  AND U8858 ( .A(n8999), .B(n9000), .Z(n8998) );
  XOR U8859 ( .A(n8997), .B(n8124), .Z(n9000) );
  XOR U8860 ( .A(n9001), .B(n9002), .Z(n8124) );
  AND U8861 ( .A(n290), .B(n9003), .Z(n9002) );
  XOR U8862 ( .A(n9004), .B(n9001), .Z(n9003) );
  XNOR U8863 ( .A(n8121), .B(n8997), .Z(n8999) );
  XOR U8864 ( .A(n9005), .B(n9006), .Z(n8121) );
  AND U8865 ( .A(n287), .B(n9007), .Z(n9006) );
  XOR U8866 ( .A(n9008), .B(n9005), .Z(n9007) );
  XOR U8867 ( .A(n9009), .B(n9010), .Z(n8997) );
  AND U8868 ( .A(n9011), .B(n9012), .Z(n9010) );
  XOR U8869 ( .A(n9009), .B(n8136), .Z(n9012) );
  XOR U8870 ( .A(n9013), .B(n9014), .Z(n8136) );
  AND U8871 ( .A(n290), .B(n9015), .Z(n9014) );
  XOR U8872 ( .A(n9016), .B(n9013), .Z(n9015) );
  XNOR U8873 ( .A(n8133), .B(n9009), .Z(n9011) );
  XOR U8874 ( .A(n9017), .B(n9018), .Z(n8133) );
  AND U8875 ( .A(n287), .B(n9019), .Z(n9018) );
  XOR U8876 ( .A(n9020), .B(n9017), .Z(n9019) );
  XOR U8877 ( .A(n9021), .B(n9022), .Z(n9009) );
  AND U8878 ( .A(n9023), .B(n9024), .Z(n9022) );
  XOR U8879 ( .A(n9021), .B(n8148), .Z(n9024) );
  XOR U8880 ( .A(n9025), .B(n9026), .Z(n8148) );
  AND U8881 ( .A(n290), .B(n9027), .Z(n9026) );
  XOR U8882 ( .A(n9028), .B(n9025), .Z(n9027) );
  XNOR U8883 ( .A(n8145), .B(n9021), .Z(n9023) );
  XOR U8884 ( .A(n9029), .B(n9030), .Z(n8145) );
  AND U8885 ( .A(n287), .B(n9031), .Z(n9030) );
  XOR U8886 ( .A(n9032), .B(n9029), .Z(n9031) );
  XOR U8887 ( .A(n9033), .B(n9034), .Z(n9021) );
  AND U8888 ( .A(n9035), .B(n9036), .Z(n9034) );
  XOR U8889 ( .A(n9033), .B(n8160), .Z(n9036) );
  XOR U8890 ( .A(n9037), .B(n9038), .Z(n8160) );
  AND U8891 ( .A(n290), .B(n9039), .Z(n9038) );
  XOR U8892 ( .A(n9040), .B(n9037), .Z(n9039) );
  XNOR U8893 ( .A(n8157), .B(n9033), .Z(n9035) );
  XOR U8894 ( .A(n9041), .B(n9042), .Z(n8157) );
  AND U8895 ( .A(n287), .B(n9043), .Z(n9042) );
  XOR U8896 ( .A(n9044), .B(n9041), .Z(n9043) );
  XOR U8897 ( .A(n9045), .B(n9046), .Z(n9033) );
  AND U8898 ( .A(n9047), .B(n9048), .Z(n9046) );
  XOR U8899 ( .A(n9045), .B(n8172), .Z(n9048) );
  XOR U8900 ( .A(n9049), .B(n9050), .Z(n8172) );
  AND U8901 ( .A(n290), .B(n9051), .Z(n9050) );
  XOR U8902 ( .A(n9052), .B(n9049), .Z(n9051) );
  XNOR U8903 ( .A(n8169), .B(n9045), .Z(n9047) );
  XOR U8904 ( .A(n9053), .B(n9054), .Z(n8169) );
  AND U8905 ( .A(n287), .B(n9055), .Z(n9054) );
  XOR U8906 ( .A(n9056), .B(n9053), .Z(n9055) );
  XOR U8907 ( .A(n9057), .B(n9058), .Z(n9045) );
  AND U8908 ( .A(n9059), .B(n9060), .Z(n9058) );
  XOR U8909 ( .A(n8184), .B(n9057), .Z(n9060) );
  XOR U8910 ( .A(n9061), .B(n9062), .Z(n8184) );
  AND U8911 ( .A(n290), .B(n9063), .Z(n9062) );
  XOR U8912 ( .A(n9061), .B(n9064), .Z(n9063) );
  XNOR U8913 ( .A(n9057), .B(n8181), .Z(n9059) );
  XOR U8914 ( .A(n9065), .B(n9066), .Z(n8181) );
  AND U8915 ( .A(n287), .B(n9067), .Z(n9066) );
  XOR U8916 ( .A(n9065), .B(n9068), .Z(n9067) );
  XOR U8917 ( .A(n9069), .B(n9070), .Z(n9057) );
  AND U8918 ( .A(n9071), .B(n9072), .Z(n9070) );
  XNOR U8919 ( .A(n9073), .B(n8197), .Z(n9072) );
  XOR U8920 ( .A(n9074), .B(n9075), .Z(n8197) );
  AND U8921 ( .A(n290), .B(n9076), .Z(n9075) );
  XOR U8922 ( .A(n9077), .B(n9074), .Z(n9076) );
  XNOR U8923 ( .A(n8194), .B(n9069), .Z(n9071) );
  XOR U8924 ( .A(n9078), .B(n9079), .Z(n8194) );
  AND U8925 ( .A(n287), .B(n9080), .Z(n9079) );
  XOR U8926 ( .A(n9081), .B(n9078), .Z(n9080) );
  IV U8927 ( .A(n9073), .Z(n9069) );
  AND U8928 ( .A(n8901), .B(n8904), .Z(n9073) );
  XNOR U8929 ( .A(n9082), .B(n9083), .Z(n8904) );
  AND U8930 ( .A(n290), .B(n9084), .Z(n9083) );
  XNOR U8931 ( .A(n9085), .B(n9082), .Z(n9084) );
  XOR U8932 ( .A(n9086), .B(n9087), .Z(n290) );
  AND U8933 ( .A(n9088), .B(n9089), .Z(n9087) );
  XNOR U8934 ( .A(n8909), .B(n9086), .Z(n9089) );
  AND U8935 ( .A(p_input[895]), .B(p_input[879]), .Z(n8909) );
  XOR U8936 ( .A(n9086), .B(n8910), .Z(n9088) );
  AND U8937 ( .A(p_input[863]), .B(p_input[847]), .Z(n8910) );
  XOR U8938 ( .A(n9090), .B(n9091), .Z(n9086) );
  AND U8939 ( .A(n9092), .B(n9093), .Z(n9091) );
  XOR U8940 ( .A(n9090), .B(n8920), .Z(n9093) );
  XNOR U8941 ( .A(p_input[878]), .B(n9094), .Z(n8920) );
  AND U8942 ( .A(n362), .B(n9095), .Z(n9094) );
  XOR U8943 ( .A(p_input[894]), .B(p_input[878]), .Z(n9095) );
  XNOR U8944 ( .A(n8917), .B(n9090), .Z(n9092) );
  XOR U8945 ( .A(n9096), .B(n9097), .Z(n8917) );
  AND U8946 ( .A(n360), .B(n9098), .Z(n9097) );
  XOR U8947 ( .A(p_input[862]), .B(p_input[846]), .Z(n9098) );
  XOR U8948 ( .A(n9099), .B(n9100), .Z(n9090) );
  AND U8949 ( .A(n9101), .B(n9102), .Z(n9100) );
  XOR U8950 ( .A(n9099), .B(n8932), .Z(n9102) );
  XNOR U8951 ( .A(p_input[877]), .B(n9103), .Z(n8932) );
  AND U8952 ( .A(n362), .B(n9104), .Z(n9103) );
  XOR U8953 ( .A(p_input[893]), .B(p_input[877]), .Z(n9104) );
  XNOR U8954 ( .A(n8929), .B(n9099), .Z(n9101) );
  XOR U8955 ( .A(n9105), .B(n9106), .Z(n8929) );
  AND U8956 ( .A(n360), .B(n9107), .Z(n9106) );
  XOR U8957 ( .A(p_input[861]), .B(p_input[845]), .Z(n9107) );
  XOR U8958 ( .A(n9108), .B(n9109), .Z(n9099) );
  AND U8959 ( .A(n9110), .B(n9111), .Z(n9109) );
  XOR U8960 ( .A(n9108), .B(n8944), .Z(n9111) );
  XNOR U8961 ( .A(p_input[876]), .B(n9112), .Z(n8944) );
  AND U8962 ( .A(n362), .B(n9113), .Z(n9112) );
  XOR U8963 ( .A(p_input[892]), .B(p_input[876]), .Z(n9113) );
  XNOR U8964 ( .A(n8941), .B(n9108), .Z(n9110) );
  XOR U8965 ( .A(n9114), .B(n9115), .Z(n8941) );
  AND U8966 ( .A(n360), .B(n9116), .Z(n9115) );
  XOR U8967 ( .A(p_input[860]), .B(p_input[844]), .Z(n9116) );
  XOR U8968 ( .A(n9117), .B(n9118), .Z(n9108) );
  AND U8969 ( .A(n9119), .B(n9120), .Z(n9118) );
  XOR U8970 ( .A(n9117), .B(n8956), .Z(n9120) );
  XNOR U8971 ( .A(p_input[875]), .B(n9121), .Z(n8956) );
  AND U8972 ( .A(n362), .B(n9122), .Z(n9121) );
  XOR U8973 ( .A(p_input[891]), .B(p_input[875]), .Z(n9122) );
  XNOR U8974 ( .A(n8953), .B(n9117), .Z(n9119) );
  XOR U8975 ( .A(n9123), .B(n9124), .Z(n8953) );
  AND U8976 ( .A(n360), .B(n9125), .Z(n9124) );
  XOR U8977 ( .A(p_input[859]), .B(p_input[843]), .Z(n9125) );
  XOR U8978 ( .A(n9126), .B(n9127), .Z(n9117) );
  AND U8979 ( .A(n9128), .B(n9129), .Z(n9127) );
  XOR U8980 ( .A(n9126), .B(n8968), .Z(n9129) );
  XNOR U8981 ( .A(p_input[874]), .B(n9130), .Z(n8968) );
  AND U8982 ( .A(n362), .B(n9131), .Z(n9130) );
  XOR U8983 ( .A(p_input[890]), .B(p_input[874]), .Z(n9131) );
  XNOR U8984 ( .A(n8965), .B(n9126), .Z(n9128) );
  XOR U8985 ( .A(n9132), .B(n9133), .Z(n8965) );
  AND U8986 ( .A(n360), .B(n9134), .Z(n9133) );
  XOR U8987 ( .A(p_input[858]), .B(p_input[842]), .Z(n9134) );
  XOR U8988 ( .A(n9135), .B(n9136), .Z(n9126) );
  AND U8989 ( .A(n9137), .B(n9138), .Z(n9136) );
  XOR U8990 ( .A(n9135), .B(n8980), .Z(n9138) );
  XNOR U8991 ( .A(p_input[873]), .B(n9139), .Z(n8980) );
  AND U8992 ( .A(n362), .B(n9140), .Z(n9139) );
  XOR U8993 ( .A(p_input[889]), .B(p_input[873]), .Z(n9140) );
  XNOR U8994 ( .A(n8977), .B(n9135), .Z(n9137) );
  XOR U8995 ( .A(n9141), .B(n9142), .Z(n8977) );
  AND U8996 ( .A(n360), .B(n9143), .Z(n9142) );
  XOR U8997 ( .A(p_input[857]), .B(p_input[841]), .Z(n9143) );
  XOR U8998 ( .A(n9144), .B(n9145), .Z(n9135) );
  AND U8999 ( .A(n9146), .B(n9147), .Z(n9145) );
  XOR U9000 ( .A(n9144), .B(n8992), .Z(n9147) );
  XNOR U9001 ( .A(p_input[872]), .B(n9148), .Z(n8992) );
  AND U9002 ( .A(n362), .B(n9149), .Z(n9148) );
  XOR U9003 ( .A(p_input[888]), .B(p_input[872]), .Z(n9149) );
  XNOR U9004 ( .A(n8989), .B(n9144), .Z(n9146) );
  XOR U9005 ( .A(n9150), .B(n9151), .Z(n8989) );
  AND U9006 ( .A(n360), .B(n9152), .Z(n9151) );
  XOR U9007 ( .A(p_input[856]), .B(p_input[840]), .Z(n9152) );
  XOR U9008 ( .A(n9153), .B(n9154), .Z(n9144) );
  AND U9009 ( .A(n9155), .B(n9156), .Z(n9154) );
  XOR U9010 ( .A(n9153), .B(n9004), .Z(n9156) );
  XNOR U9011 ( .A(p_input[871]), .B(n9157), .Z(n9004) );
  AND U9012 ( .A(n362), .B(n9158), .Z(n9157) );
  XOR U9013 ( .A(p_input[887]), .B(p_input[871]), .Z(n9158) );
  XNOR U9014 ( .A(n9001), .B(n9153), .Z(n9155) );
  XOR U9015 ( .A(n9159), .B(n9160), .Z(n9001) );
  AND U9016 ( .A(n360), .B(n9161), .Z(n9160) );
  XOR U9017 ( .A(p_input[855]), .B(p_input[839]), .Z(n9161) );
  XOR U9018 ( .A(n9162), .B(n9163), .Z(n9153) );
  AND U9019 ( .A(n9164), .B(n9165), .Z(n9163) );
  XOR U9020 ( .A(n9162), .B(n9016), .Z(n9165) );
  XNOR U9021 ( .A(p_input[870]), .B(n9166), .Z(n9016) );
  AND U9022 ( .A(n362), .B(n9167), .Z(n9166) );
  XOR U9023 ( .A(p_input[886]), .B(p_input[870]), .Z(n9167) );
  XNOR U9024 ( .A(n9013), .B(n9162), .Z(n9164) );
  XOR U9025 ( .A(n9168), .B(n9169), .Z(n9013) );
  AND U9026 ( .A(n360), .B(n9170), .Z(n9169) );
  XOR U9027 ( .A(p_input[854]), .B(p_input[838]), .Z(n9170) );
  XOR U9028 ( .A(n9171), .B(n9172), .Z(n9162) );
  AND U9029 ( .A(n9173), .B(n9174), .Z(n9172) );
  XOR U9030 ( .A(n9171), .B(n9028), .Z(n9174) );
  XNOR U9031 ( .A(p_input[869]), .B(n9175), .Z(n9028) );
  AND U9032 ( .A(n362), .B(n9176), .Z(n9175) );
  XOR U9033 ( .A(p_input[885]), .B(p_input[869]), .Z(n9176) );
  XNOR U9034 ( .A(n9025), .B(n9171), .Z(n9173) );
  XOR U9035 ( .A(n9177), .B(n9178), .Z(n9025) );
  AND U9036 ( .A(n360), .B(n9179), .Z(n9178) );
  XOR U9037 ( .A(p_input[853]), .B(p_input[837]), .Z(n9179) );
  XOR U9038 ( .A(n9180), .B(n9181), .Z(n9171) );
  AND U9039 ( .A(n9182), .B(n9183), .Z(n9181) );
  XOR U9040 ( .A(n9180), .B(n9040), .Z(n9183) );
  XNOR U9041 ( .A(p_input[868]), .B(n9184), .Z(n9040) );
  AND U9042 ( .A(n362), .B(n9185), .Z(n9184) );
  XOR U9043 ( .A(p_input[884]), .B(p_input[868]), .Z(n9185) );
  XNOR U9044 ( .A(n9037), .B(n9180), .Z(n9182) );
  XOR U9045 ( .A(n9186), .B(n9187), .Z(n9037) );
  AND U9046 ( .A(n360), .B(n9188), .Z(n9187) );
  XOR U9047 ( .A(p_input[852]), .B(p_input[836]), .Z(n9188) );
  XOR U9048 ( .A(n9189), .B(n9190), .Z(n9180) );
  AND U9049 ( .A(n9191), .B(n9192), .Z(n9190) );
  XOR U9050 ( .A(n9189), .B(n9052), .Z(n9192) );
  XNOR U9051 ( .A(p_input[867]), .B(n9193), .Z(n9052) );
  AND U9052 ( .A(n362), .B(n9194), .Z(n9193) );
  XOR U9053 ( .A(p_input[883]), .B(p_input[867]), .Z(n9194) );
  XNOR U9054 ( .A(n9049), .B(n9189), .Z(n9191) );
  XOR U9055 ( .A(n9195), .B(n9196), .Z(n9049) );
  AND U9056 ( .A(n360), .B(n9197), .Z(n9196) );
  XOR U9057 ( .A(p_input[851]), .B(p_input[835]), .Z(n9197) );
  XOR U9058 ( .A(n9198), .B(n9199), .Z(n9189) );
  AND U9059 ( .A(n9200), .B(n9201), .Z(n9199) );
  XOR U9060 ( .A(n9064), .B(n9198), .Z(n9201) );
  XNOR U9061 ( .A(p_input[866]), .B(n9202), .Z(n9064) );
  AND U9062 ( .A(n362), .B(n9203), .Z(n9202) );
  XOR U9063 ( .A(p_input[882]), .B(p_input[866]), .Z(n9203) );
  XNOR U9064 ( .A(n9198), .B(n9061), .Z(n9200) );
  XOR U9065 ( .A(n9204), .B(n9205), .Z(n9061) );
  AND U9066 ( .A(n360), .B(n9206), .Z(n9205) );
  XOR U9067 ( .A(p_input[850]), .B(p_input[834]), .Z(n9206) );
  XOR U9068 ( .A(n9207), .B(n9208), .Z(n9198) );
  AND U9069 ( .A(n9209), .B(n9210), .Z(n9208) );
  XNOR U9070 ( .A(n9211), .B(n9077), .Z(n9210) );
  XNOR U9071 ( .A(p_input[865]), .B(n9212), .Z(n9077) );
  AND U9072 ( .A(n362), .B(n9213), .Z(n9212) );
  XNOR U9073 ( .A(p_input[881]), .B(n9214), .Z(n9213) );
  IV U9074 ( .A(p_input[865]), .Z(n9214) );
  XNOR U9075 ( .A(n9074), .B(n9207), .Z(n9209) );
  XNOR U9076 ( .A(p_input[833]), .B(n9215), .Z(n9074) );
  AND U9077 ( .A(n360), .B(n9216), .Z(n9215) );
  XOR U9078 ( .A(p_input[849]), .B(p_input[833]), .Z(n9216) );
  IV U9079 ( .A(n9211), .Z(n9207) );
  AND U9080 ( .A(n9082), .B(n9085), .Z(n9211) );
  XOR U9081 ( .A(p_input[864]), .B(n9217), .Z(n9085) );
  AND U9082 ( .A(n362), .B(n9218), .Z(n9217) );
  XOR U9083 ( .A(p_input[880]), .B(p_input[864]), .Z(n9218) );
  XOR U9084 ( .A(n9219), .B(n9220), .Z(n362) );
  AND U9085 ( .A(n9221), .B(n9222), .Z(n9220) );
  XNOR U9086 ( .A(p_input[895]), .B(n9219), .Z(n9222) );
  XOR U9087 ( .A(n9219), .B(p_input[879]), .Z(n9221) );
  XOR U9088 ( .A(n9223), .B(n9224), .Z(n9219) );
  AND U9089 ( .A(n9225), .B(n9226), .Z(n9224) );
  XNOR U9090 ( .A(p_input[894]), .B(n9223), .Z(n9226) );
  XOR U9091 ( .A(n9223), .B(p_input[878]), .Z(n9225) );
  XOR U9092 ( .A(n9227), .B(n9228), .Z(n9223) );
  AND U9093 ( .A(n9229), .B(n9230), .Z(n9228) );
  XNOR U9094 ( .A(p_input[893]), .B(n9227), .Z(n9230) );
  XOR U9095 ( .A(n9227), .B(p_input[877]), .Z(n9229) );
  XOR U9096 ( .A(n9231), .B(n9232), .Z(n9227) );
  AND U9097 ( .A(n9233), .B(n9234), .Z(n9232) );
  XNOR U9098 ( .A(p_input[892]), .B(n9231), .Z(n9234) );
  XOR U9099 ( .A(n9231), .B(p_input[876]), .Z(n9233) );
  XOR U9100 ( .A(n9235), .B(n9236), .Z(n9231) );
  AND U9101 ( .A(n9237), .B(n9238), .Z(n9236) );
  XNOR U9102 ( .A(p_input[891]), .B(n9235), .Z(n9238) );
  XOR U9103 ( .A(n9235), .B(p_input[875]), .Z(n9237) );
  XOR U9104 ( .A(n9239), .B(n9240), .Z(n9235) );
  AND U9105 ( .A(n9241), .B(n9242), .Z(n9240) );
  XNOR U9106 ( .A(p_input[890]), .B(n9239), .Z(n9242) );
  XOR U9107 ( .A(n9239), .B(p_input[874]), .Z(n9241) );
  XOR U9108 ( .A(n9243), .B(n9244), .Z(n9239) );
  AND U9109 ( .A(n9245), .B(n9246), .Z(n9244) );
  XNOR U9110 ( .A(p_input[889]), .B(n9243), .Z(n9246) );
  XOR U9111 ( .A(n9243), .B(p_input[873]), .Z(n9245) );
  XOR U9112 ( .A(n9247), .B(n9248), .Z(n9243) );
  AND U9113 ( .A(n9249), .B(n9250), .Z(n9248) );
  XNOR U9114 ( .A(p_input[888]), .B(n9247), .Z(n9250) );
  XOR U9115 ( .A(n9247), .B(p_input[872]), .Z(n9249) );
  XOR U9116 ( .A(n9251), .B(n9252), .Z(n9247) );
  AND U9117 ( .A(n9253), .B(n9254), .Z(n9252) );
  XNOR U9118 ( .A(p_input[887]), .B(n9251), .Z(n9254) );
  XOR U9119 ( .A(n9251), .B(p_input[871]), .Z(n9253) );
  XOR U9120 ( .A(n9255), .B(n9256), .Z(n9251) );
  AND U9121 ( .A(n9257), .B(n9258), .Z(n9256) );
  XNOR U9122 ( .A(p_input[886]), .B(n9255), .Z(n9258) );
  XOR U9123 ( .A(n9255), .B(p_input[870]), .Z(n9257) );
  XOR U9124 ( .A(n9259), .B(n9260), .Z(n9255) );
  AND U9125 ( .A(n9261), .B(n9262), .Z(n9260) );
  XNOR U9126 ( .A(p_input[885]), .B(n9259), .Z(n9262) );
  XOR U9127 ( .A(n9259), .B(p_input[869]), .Z(n9261) );
  XOR U9128 ( .A(n9263), .B(n9264), .Z(n9259) );
  AND U9129 ( .A(n9265), .B(n9266), .Z(n9264) );
  XNOR U9130 ( .A(p_input[884]), .B(n9263), .Z(n9266) );
  XOR U9131 ( .A(n9263), .B(p_input[868]), .Z(n9265) );
  XOR U9132 ( .A(n9267), .B(n9268), .Z(n9263) );
  AND U9133 ( .A(n9269), .B(n9270), .Z(n9268) );
  XNOR U9134 ( .A(p_input[883]), .B(n9267), .Z(n9270) );
  XOR U9135 ( .A(n9267), .B(p_input[867]), .Z(n9269) );
  XOR U9136 ( .A(n9271), .B(n9272), .Z(n9267) );
  AND U9137 ( .A(n9273), .B(n9274), .Z(n9272) );
  XNOR U9138 ( .A(p_input[882]), .B(n9271), .Z(n9274) );
  XOR U9139 ( .A(n9271), .B(p_input[866]), .Z(n9273) );
  XNOR U9140 ( .A(n9275), .B(n9276), .Z(n9271) );
  AND U9141 ( .A(n9277), .B(n9278), .Z(n9276) );
  XOR U9142 ( .A(p_input[881]), .B(n9275), .Z(n9278) );
  XNOR U9143 ( .A(p_input[865]), .B(n9275), .Z(n9277) );
  AND U9144 ( .A(p_input[880]), .B(n9279), .Z(n9275) );
  IV U9145 ( .A(p_input[864]), .Z(n9279) );
  XNOR U9146 ( .A(p_input[832]), .B(n9280), .Z(n9082) );
  AND U9147 ( .A(n360), .B(n9281), .Z(n9280) );
  XOR U9148 ( .A(p_input[848]), .B(p_input[832]), .Z(n9281) );
  XOR U9149 ( .A(n9282), .B(n9283), .Z(n360) );
  AND U9150 ( .A(n9284), .B(n9285), .Z(n9283) );
  XNOR U9151 ( .A(p_input[863]), .B(n9282), .Z(n9285) );
  XOR U9152 ( .A(n9282), .B(p_input[847]), .Z(n9284) );
  XOR U9153 ( .A(n9286), .B(n9287), .Z(n9282) );
  AND U9154 ( .A(n9288), .B(n9289), .Z(n9287) );
  XNOR U9155 ( .A(p_input[862]), .B(n9286), .Z(n9289) );
  XNOR U9156 ( .A(n9286), .B(n9096), .Z(n9288) );
  IV U9157 ( .A(p_input[846]), .Z(n9096) );
  XOR U9158 ( .A(n9290), .B(n9291), .Z(n9286) );
  AND U9159 ( .A(n9292), .B(n9293), .Z(n9291) );
  XNOR U9160 ( .A(p_input[861]), .B(n9290), .Z(n9293) );
  XNOR U9161 ( .A(n9290), .B(n9105), .Z(n9292) );
  IV U9162 ( .A(p_input[845]), .Z(n9105) );
  XOR U9163 ( .A(n9294), .B(n9295), .Z(n9290) );
  AND U9164 ( .A(n9296), .B(n9297), .Z(n9295) );
  XNOR U9165 ( .A(p_input[860]), .B(n9294), .Z(n9297) );
  XNOR U9166 ( .A(n9294), .B(n9114), .Z(n9296) );
  IV U9167 ( .A(p_input[844]), .Z(n9114) );
  XOR U9168 ( .A(n9298), .B(n9299), .Z(n9294) );
  AND U9169 ( .A(n9300), .B(n9301), .Z(n9299) );
  XNOR U9170 ( .A(p_input[859]), .B(n9298), .Z(n9301) );
  XNOR U9171 ( .A(n9298), .B(n9123), .Z(n9300) );
  IV U9172 ( .A(p_input[843]), .Z(n9123) );
  XOR U9173 ( .A(n9302), .B(n9303), .Z(n9298) );
  AND U9174 ( .A(n9304), .B(n9305), .Z(n9303) );
  XNOR U9175 ( .A(p_input[858]), .B(n9302), .Z(n9305) );
  XNOR U9176 ( .A(n9302), .B(n9132), .Z(n9304) );
  IV U9177 ( .A(p_input[842]), .Z(n9132) );
  XOR U9178 ( .A(n9306), .B(n9307), .Z(n9302) );
  AND U9179 ( .A(n9308), .B(n9309), .Z(n9307) );
  XNOR U9180 ( .A(p_input[857]), .B(n9306), .Z(n9309) );
  XNOR U9181 ( .A(n9306), .B(n9141), .Z(n9308) );
  IV U9182 ( .A(p_input[841]), .Z(n9141) );
  XOR U9183 ( .A(n9310), .B(n9311), .Z(n9306) );
  AND U9184 ( .A(n9312), .B(n9313), .Z(n9311) );
  XNOR U9185 ( .A(p_input[856]), .B(n9310), .Z(n9313) );
  XNOR U9186 ( .A(n9310), .B(n9150), .Z(n9312) );
  IV U9187 ( .A(p_input[840]), .Z(n9150) );
  XOR U9188 ( .A(n9314), .B(n9315), .Z(n9310) );
  AND U9189 ( .A(n9316), .B(n9317), .Z(n9315) );
  XNOR U9190 ( .A(p_input[855]), .B(n9314), .Z(n9317) );
  XNOR U9191 ( .A(n9314), .B(n9159), .Z(n9316) );
  IV U9192 ( .A(p_input[839]), .Z(n9159) );
  XOR U9193 ( .A(n9318), .B(n9319), .Z(n9314) );
  AND U9194 ( .A(n9320), .B(n9321), .Z(n9319) );
  XNOR U9195 ( .A(p_input[854]), .B(n9318), .Z(n9321) );
  XNOR U9196 ( .A(n9318), .B(n9168), .Z(n9320) );
  IV U9197 ( .A(p_input[838]), .Z(n9168) );
  XOR U9198 ( .A(n9322), .B(n9323), .Z(n9318) );
  AND U9199 ( .A(n9324), .B(n9325), .Z(n9323) );
  XNOR U9200 ( .A(p_input[853]), .B(n9322), .Z(n9325) );
  XNOR U9201 ( .A(n9322), .B(n9177), .Z(n9324) );
  IV U9202 ( .A(p_input[837]), .Z(n9177) );
  XOR U9203 ( .A(n9326), .B(n9327), .Z(n9322) );
  AND U9204 ( .A(n9328), .B(n9329), .Z(n9327) );
  XNOR U9205 ( .A(p_input[852]), .B(n9326), .Z(n9329) );
  XNOR U9206 ( .A(n9326), .B(n9186), .Z(n9328) );
  IV U9207 ( .A(p_input[836]), .Z(n9186) );
  XOR U9208 ( .A(n9330), .B(n9331), .Z(n9326) );
  AND U9209 ( .A(n9332), .B(n9333), .Z(n9331) );
  XNOR U9210 ( .A(p_input[851]), .B(n9330), .Z(n9333) );
  XNOR U9211 ( .A(n9330), .B(n9195), .Z(n9332) );
  IV U9212 ( .A(p_input[835]), .Z(n9195) );
  XOR U9213 ( .A(n9334), .B(n9335), .Z(n9330) );
  AND U9214 ( .A(n9336), .B(n9337), .Z(n9335) );
  XNOR U9215 ( .A(p_input[850]), .B(n9334), .Z(n9337) );
  XNOR U9216 ( .A(n9334), .B(n9204), .Z(n9336) );
  IV U9217 ( .A(p_input[834]), .Z(n9204) );
  XNOR U9218 ( .A(n9338), .B(n9339), .Z(n9334) );
  AND U9219 ( .A(n9340), .B(n9341), .Z(n9339) );
  XOR U9220 ( .A(p_input[849]), .B(n9338), .Z(n9341) );
  XNOR U9221 ( .A(p_input[833]), .B(n9338), .Z(n9340) );
  AND U9222 ( .A(p_input[848]), .B(n9342), .Z(n9338) );
  IV U9223 ( .A(p_input[832]), .Z(n9342) );
  XOR U9224 ( .A(n9343), .B(n9344), .Z(n8901) );
  AND U9225 ( .A(n287), .B(n9345), .Z(n9344) );
  XNOR U9226 ( .A(n9346), .B(n9343), .Z(n9345) );
  XOR U9227 ( .A(n9347), .B(n9348), .Z(n287) );
  AND U9228 ( .A(n9349), .B(n9350), .Z(n9348) );
  XNOR U9229 ( .A(n8912), .B(n9347), .Z(n9350) );
  AND U9230 ( .A(p_input[831]), .B(p_input[815]), .Z(n8912) );
  XOR U9231 ( .A(n9347), .B(n8911), .Z(n9349) );
  AND U9232 ( .A(p_input[783]), .B(p_input[799]), .Z(n8911) );
  XOR U9233 ( .A(n9351), .B(n9352), .Z(n9347) );
  AND U9234 ( .A(n9353), .B(n9354), .Z(n9352) );
  XOR U9235 ( .A(n9351), .B(n8924), .Z(n9354) );
  XNOR U9236 ( .A(p_input[814]), .B(n9355), .Z(n8924) );
  AND U9237 ( .A(n366), .B(n9356), .Z(n9355) );
  XOR U9238 ( .A(p_input[830]), .B(p_input[814]), .Z(n9356) );
  XNOR U9239 ( .A(n8921), .B(n9351), .Z(n9353) );
  XOR U9240 ( .A(n9357), .B(n9358), .Z(n8921) );
  AND U9241 ( .A(n363), .B(n9359), .Z(n9358) );
  XOR U9242 ( .A(p_input[798]), .B(p_input[782]), .Z(n9359) );
  XOR U9243 ( .A(n9360), .B(n9361), .Z(n9351) );
  AND U9244 ( .A(n9362), .B(n9363), .Z(n9361) );
  XOR U9245 ( .A(n9360), .B(n8936), .Z(n9363) );
  XNOR U9246 ( .A(p_input[813]), .B(n9364), .Z(n8936) );
  AND U9247 ( .A(n366), .B(n9365), .Z(n9364) );
  XOR U9248 ( .A(p_input[829]), .B(p_input[813]), .Z(n9365) );
  XNOR U9249 ( .A(n8933), .B(n9360), .Z(n9362) );
  XOR U9250 ( .A(n9366), .B(n9367), .Z(n8933) );
  AND U9251 ( .A(n363), .B(n9368), .Z(n9367) );
  XOR U9252 ( .A(p_input[797]), .B(p_input[781]), .Z(n9368) );
  XOR U9253 ( .A(n9369), .B(n9370), .Z(n9360) );
  AND U9254 ( .A(n9371), .B(n9372), .Z(n9370) );
  XOR U9255 ( .A(n9369), .B(n8948), .Z(n9372) );
  XNOR U9256 ( .A(p_input[812]), .B(n9373), .Z(n8948) );
  AND U9257 ( .A(n366), .B(n9374), .Z(n9373) );
  XOR U9258 ( .A(p_input[828]), .B(p_input[812]), .Z(n9374) );
  XNOR U9259 ( .A(n8945), .B(n9369), .Z(n9371) );
  XOR U9260 ( .A(n9375), .B(n9376), .Z(n8945) );
  AND U9261 ( .A(n363), .B(n9377), .Z(n9376) );
  XOR U9262 ( .A(p_input[796]), .B(p_input[780]), .Z(n9377) );
  XOR U9263 ( .A(n9378), .B(n9379), .Z(n9369) );
  AND U9264 ( .A(n9380), .B(n9381), .Z(n9379) );
  XOR U9265 ( .A(n9378), .B(n8960), .Z(n9381) );
  XNOR U9266 ( .A(p_input[811]), .B(n9382), .Z(n8960) );
  AND U9267 ( .A(n366), .B(n9383), .Z(n9382) );
  XOR U9268 ( .A(p_input[827]), .B(p_input[811]), .Z(n9383) );
  XNOR U9269 ( .A(n8957), .B(n9378), .Z(n9380) );
  XOR U9270 ( .A(n9384), .B(n9385), .Z(n8957) );
  AND U9271 ( .A(n363), .B(n9386), .Z(n9385) );
  XOR U9272 ( .A(p_input[795]), .B(p_input[779]), .Z(n9386) );
  XOR U9273 ( .A(n9387), .B(n9388), .Z(n9378) );
  AND U9274 ( .A(n9389), .B(n9390), .Z(n9388) );
  XOR U9275 ( .A(n9387), .B(n8972), .Z(n9390) );
  XNOR U9276 ( .A(p_input[810]), .B(n9391), .Z(n8972) );
  AND U9277 ( .A(n366), .B(n9392), .Z(n9391) );
  XOR U9278 ( .A(p_input[826]), .B(p_input[810]), .Z(n9392) );
  XNOR U9279 ( .A(n8969), .B(n9387), .Z(n9389) );
  XOR U9280 ( .A(n9393), .B(n9394), .Z(n8969) );
  AND U9281 ( .A(n363), .B(n9395), .Z(n9394) );
  XOR U9282 ( .A(p_input[794]), .B(p_input[778]), .Z(n9395) );
  XOR U9283 ( .A(n9396), .B(n9397), .Z(n9387) );
  AND U9284 ( .A(n9398), .B(n9399), .Z(n9397) );
  XOR U9285 ( .A(n9396), .B(n8984), .Z(n9399) );
  XNOR U9286 ( .A(p_input[809]), .B(n9400), .Z(n8984) );
  AND U9287 ( .A(n366), .B(n9401), .Z(n9400) );
  XOR U9288 ( .A(p_input[825]), .B(p_input[809]), .Z(n9401) );
  XNOR U9289 ( .A(n8981), .B(n9396), .Z(n9398) );
  XOR U9290 ( .A(n9402), .B(n9403), .Z(n8981) );
  AND U9291 ( .A(n363), .B(n9404), .Z(n9403) );
  XOR U9292 ( .A(p_input[793]), .B(p_input[777]), .Z(n9404) );
  XOR U9293 ( .A(n9405), .B(n9406), .Z(n9396) );
  AND U9294 ( .A(n9407), .B(n9408), .Z(n9406) );
  XOR U9295 ( .A(n9405), .B(n8996), .Z(n9408) );
  XNOR U9296 ( .A(p_input[808]), .B(n9409), .Z(n8996) );
  AND U9297 ( .A(n366), .B(n9410), .Z(n9409) );
  XOR U9298 ( .A(p_input[824]), .B(p_input[808]), .Z(n9410) );
  XNOR U9299 ( .A(n8993), .B(n9405), .Z(n9407) );
  XOR U9300 ( .A(n9411), .B(n9412), .Z(n8993) );
  AND U9301 ( .A(n363), .B(n9413), .Z(n9412) );
  XOR U9302 ( .A(p_input[792]), .B(p_input[776]), .Z(n9413) );
  XOR U9303 ( .A(n9414), .B(n9415), .Z(n9405) );
  AND U9304 ( .A(n9416), .B(n9417), .Z(n9415) );
  XOR U9305 ( .A(n9414), .B(n9008), .Z(n9417) );
  XNOR U9306 ( .A(p_input[807]), .B(n9418), .Z(n9008) );
  AND U9307 ( .A(n366), .B(n9419), .Z(n9418) );
  XOR U9308 ( .A(p_input[823]), .B(p_input[807]), .Z(n9419) );
  XNOR U9309 ( .A(n9005), .B(n9414), .Z(n9416) );
  XOR U9310 ( .A(n9420), .B(n9421), .Z(n9005) );
  AND U9311 ( .A(n363), .B(n9422), .Z(n9421) );
  XOR U9312 ( .A(p_input[791]), .B(p_input[775]), .Z(n9422) );
  XOR U9313 ( .A(n9423), .B(n9424), .Z(n9414) );
  AND U9314 ( .A(n9425), .B(n9426), .Z(n9424) );
  XOR U9315 ( .A(n9423), .B(n9020), .Z(n9426) );
  XNOR U9316 ( .A(p_input[806]), .B(n9427), .Z(n9020) );
  AND U9317 ( .A(n366), .B(n9428), .Z(n9427) );
  XOR U9318 ( .A(p_input[822]), .B(p_input[806]), .Z(n9428) );
  XNOR U9319 ( .A(n9017), .B(n9423), .Z(n9425) );
  XOR U9320 ( .A(n9429), .B(n9430), .Z(n9017) );
  AND U9321 ( .A(n363), .B(n9431), .Z(n9430) );
  XOR U9322 ( .A(p_input[790]), .B(p_input[774]), .Z(n9431) );
  XOR U9323 ( .A(n9432), .B(n9433), .Z(n9423) );
  AND U9324 ( .A(n9434), .B(n9435), .Z(n9433) );
  XOR U9325 ( .A(n9432), .B(n9032), .Z(n9435) );
  XNOR U9326 ( .A(p_input[805]), .B(n9436), .Z(n9032) );
  AND U9327 ( .A(n366), .B(n9437), .Z(n9436) );
  XOR U9328 ( .A(p_input[821]), .B(p_input[805]), .Z(n9437) );
  XNOR U9329 ( .A(n9029), .B(n9432), .Z(n9434) );
  XOR U9330 ( .A(n9438), .B(n9439), .Z(n9029) );
  AND U9331 ( .A(n363), .B(n9440), .Z(n9439) );
  XOR U9332 ( .A(p_input[789]), .B(p_input[773]), .Z(n9440) );
  XOR U9333 ( .A(n9441), .B(n9442), .Z(n9432) );
  AND U9334 ( .A(n9443), .B(n9444), .Z(n9442) );
  XOR U9335 ( .A(n9441), .B(n9044), .Z(n9444) );
  XNOR U9336 ( .A(p_input[804]), .B(n9445), .Z(n9044) );
  AND U9337 ( .A(n366), .B(n9446), .Z(n9445) );
  XOR U9338 ( .A(p_input[820]), .B(p_input[804]), .Z(n9446) );
  XNOR U9339 ( .A(n9041), .B(n9441), .Z(n9443) );
  XOR U9340 ( .A(n9447), .B(n9448), .Z(n9041) );
  AND U9341 ( .A(n363), .B(n9449), .Z(n9448) );
  XOR U9342 ( .A(p_input[788]), .B(p_input[772]), .Z(n9449) );
  XOR U9343 ( .A(n9450), .B(n9451), .Z(n9441) );
  AND U9344 ( .A(n9452), .B(n9453), .Z(n9451) );
  XOR U9345 ( .A(n9450), .B(n9056), .Z(n9453) );
  XNOR U9346 ( .A(p_input[803]), .B(n9454), .Z(n9056) );
  AND U9347 ( .A(n366), .B(n9455), .Z(n9454) );
  XOR U9348 ( .A(p_input[819]), .B(p_input[803]), .Z(n9455) );
  XNOR U9349 ( .A(n9053), .B(n9450), .Z(n9452) );
  XOR U9350 ( .A(n9456), .B(n9457), .Z(n9053) );
  AND U9351 ( .A(n363), .B(n9458), .Z(n9457) );
  XOR U9352 ( .A(p_input[787]), .B(p_input[771]), .Z(n9458) );
  XOR U9353 ( .A(n9459), .B(n9460), .Z(n9450) );
  AND U9354 ( .A(n9461), .B(n9462), .Z(n9460) );
  XOR U9355 ( .A(n9068), .B(n9459), .Z(n9462) );
  XNOR U9356 ( .A(p_input[802]), .B(n9463), .Z(n9068) );
  AND U9357 ( .A(n366), .B(n9464), .Z(n9463) );
  XOR U9358 ( .A(p_input[818]), .B(p_input[802]), .Z(n9464) );
  XNOR U9359 ( .A(n9459), .B(n9065), .Z(n9461) );
  XOR U9360 ( .A(n9465), .B(n9466), .Z(n9065) );
  AND U9361 ( .A(n363), .B(n9467), .Z(n9466) );
  XOR U9362 ( .A(p_input[786]), .B(p_input[770]), .Z(n9467) );
  XOR U9363 ( .A(n9468), .B(n9469), .Z(n9459) );
  AND U9364 ( .A(n9470), .B(n9471), .Z(n9469) );
  XNOR U9365 ( .A(n9472), .B(n9081), .Z(n9471) );
  XNOR U9366 ( .A(p_input[801]), .B(n9473), .Z(n9081) );
  AND U9367 ( .A(n366), .B(n9474), .Z(n9473) );
  XNOR U9368 ( .A(p_input[817]), .B(n9475), .Z(n9474) );
  IV U9369 ( .A(p_input[801]), .Z(n9475) );
  XNOR U9370 ( .A(n9078), .B(n9468), .Z(n9470) );
  XNOR U9371 ( .A(p_input[769]), .B(n9476), .Z(n9078) );
  AND U9372 ( .A(n363), .B(n9477), .Z(n9476) );
  XOR U9373 ( .A(p_input[785]), .B(p_input[769]), .Z(n9477) );
  IV U9374 ( .A(n9472), .Z(n9468) );
  AND U9375 ( .A(n9343), .B(n9346), .Z(n9472) );
  XOR U9376 ( .A(p_input[800]), .B(n9478), .Z(n9346) );
  AND U9377 ( .A(n366), .B(n9479), .Z(n9478) );
  XOR U9378 ( .A(p_input[816]), .B(p_input[800]), .Z(n9479) );
  XOR U9379 ( .A(n9480), .B(n9481), .Z(n366) );
  AND U9380 ( .A(n9482), .B(n9483), .Z(n9481) );
  XNOR U9381 ( .A(p_input[831]), .B(n9480), .Z(n9483) );
  XOR U9382 ( .A(n9480), .B(p_input[815]), .Z(n9482) );
  XOR U9383 ( .A(n9484), .B(n9485), .Z(n9480) );
  AND U9384 ( .A(n9486), .B(n9487), .Z(n9485) );
  XNOR U9385 ( .A(p_input[830]), .B(n9484), .Z(n9487) );
  XOR U9386 ( .A(n9484), .B(p_input[814]), .Z(n9486) );
  XOR U9387 ( .A(n9488), .B(n9489), .Z(n9484) );
  AND U9388 ( .A(n9490), .B(n9491), .Z(n9489) );
  XNOR U9389 ( .A(p_input[829]), .B(n9488), .Z(n9491) );
  XOR U9390 ( .A(n9488), .B(p_input[813]), .Z(n9490) );
  XOR U9391 ( .A(n9492), .B(n9493), .Z(n9488) );
  AND U9392 ( .A(n9494), .B(n9495), .Z(n9493) );
  XNOR U9393 ( .A(p_input[828]), .B(n9492), .Z(n9495) );
  XOR U9394 ( .A(n9492), .B(p_input[812]), .Z(n9494) );
  XOR U9395 ( .A(n9496), .B(n9497), .Z(n9492) );
  AND U9396 ( .A(n9498), .B(n9499), .Z(n9497) );
  XNOR U9397 ( .A(p_input[827]), .B(n9496), .Z(n9499) );
  XOR U9398 ( .A(n9496), .B(p_input[811]), .Z(n9498) );
  XOR U9399 ( .A(n9500), .B(n9501), .Z(n9496) );
  AND U9400 ( .A(n9502), .B(n9503), .Z(n9501) );
  XNOR U9401 ( .A(p_input[826]), .B(n9500), .Z(n9503) );
  XOR U9402 ( .A(n9500), .B(p_input[810]), .Z(n9502) );
  XOR U9403 ( .A(n9504), .B(n9505), .Z(n9500) );
  AND U9404 ( .A(n9506), .B(n9507), .Z(n9505) );
  XNOR U9405 ( .A(p_input[825]), .B(n9504), .Z(n9507) );
  XOR U9406 ( .A(n9504), .B(p_input[809]), .Z(n9506) );
  XOR U9407 ( .A(n9508), .B(n9509), .Z(n9504) );
  AND U9408 ( .A(n9510), .B(n9511), .Z(n9509) );
  XNOR U9409 ( .A(p_input[824]), .B(n9508), .Z(n9511) );
  XOR U9410 ( .A(n9508), .B(p_input[808]), .Z(n9510) );
  XOR U9411 ( .A(n9512), .B(n9513), .Z(n9508) );
  AND U9412 ( .A(n9514), .B(n9515), .Z(n9513) );
  XNOR U9413 ( .A(p_input[823]), .B(n9512), .Z(n9515) );
  XOR U9414 ( .A(n9512), .B(p_input[807]), .Z(n9514) );
  XOR U9415 ( .A(n9516), .B(n9517), .Z(n9512) );
  AND U9416 ( .A(n9518), .B(n9519), .Z(n9517) );
  XNOR U9417 ( .A(p_input[822]), .B(n9516), .Z(n9519) );
  XOR U9418 ( .A(n9516), .B(p_input[806]), .Z(n9518) );
  XOR U9419 ( .A(n9520), .B(n9521), .Z(n9516) );
  AND U9420 ( .A(n9522), .B(n9523), .Z(n9521) );
  XNOR U9421 ( .A(p_input[821]), .B(n9520), .Z(n9523) );
  XOR U9422 ( .A(n9520), .B(p_input[805]), .Z(n9522) );
  XOR U9423 ( .A(n9524), .B(n9525), .Z(n9520) );
  AND U9424 ( .A(n9526), .B(n9527), .Z(n9525) );
  XNOR U9425 ( .A(p_input[820]), .B(n9524), .Z(n9527) );
  XOR U9426 ( .A(n9524), .B(p_input[804]), .Z(n9526) );
  XOR U9427 ( .A(n9528), .B(n9529), .Z(n9524) );
  AND U9428 ( .A(n9530), .B(n9531), .Z(n9529) );
  XNOR U9429 ( .A(p_input[819]), .B(n9528), .Z(n9531) );
  XOR U9430 ( .A(n9528), .B(p_input[803]), .Z(n9530) );
  XOR U9431 ( .A(n9532), .B(n9533), .Z(n9528) );
  AND U9432 ( .A(n9534), .B(n9535), .Z(n9533) );
  XNOR U9433 ( .A(p_input[818]), .B(n9532), .Z(n9535) );
  XOR U9434 ( .A(n9532), .B(p_input[802]), .Z(n9534) );
  XNOR U9435 ( .A(n9536), .B(n9537), .Z(n9532) );
  AND U9436 ( .A(n9538), .B(n9539), .Z(n9537) );
  XOR U9437 ( .A(p_input[817]), .B(n9536), .Z(n9539) );
  XNOR U9438 ( .A(p_input[801]), .B(n9536), .Z(n9538) );
  AND U9439 ( .A(p_input[816]), .B(n9540), .Z(n9536) );
  IV U9440 ( .A(p_input[800]), .Z(n9540) );
  XNOR U9441 ( .A(p_input[768]), .B(n9541), .Z(n9343) );
  AND U9442 ( .A(n363), .B(n9542), .Z(n9541) );
  XOR U9443 ( .A(p_input[784]), .B(p_input[768]), .Z(n9542) );
  XOR U9444 ( .A(n9543), .B(n9544), .Z(n363) );
  AND U9445 ( .A(n9545), .B(n9546), .Z(n9544) );
  XNOR U9446 ( .A(p_input[799]), .B(n9543), .Z(n9546) );
  XOR U9447 ( .A(n9543), .B(p_input[783]), .Z(n9545) );
  XOR U9448 ( .A(n9547), .B(n9548), .Z(n9543) );
  AND U9449 ( .A(n9549), .B(n9550), .Z(n9548) );
  XNOR U9450 ( .A(p_input[798]), .B(n9547), .Z(n9550) );
  XNOR U9451 ( .A(n9547), .B(n9357), .Z(n9549) );
  IV U9452 ( .A(p_input[782]), .Z(n9357) );
  XOR U9453 ( .A(n9551), .B(n9552), .Z(n9547) );
  AND U9454 ( .A(n9553), .B(n9554), .Z(n9552) );
  XNOR U9455 ( .A(p_input[797]), .B(n9551), .Z(n9554) );
  XNOR U9456 ( .A(n9551), .B(n9366), .Z(n9553) );
  IV U9457 ( .A(p_input[781]), .Z(n9366) );
  XOR U9458 ( .A(n9555), .B(n9556), .Z(n9551) );
  AND U9459 ( .A(n9557), .B(n9558), .Z(n9556) );
  XNOR U9460 ( .A(p_input[796]), .B(n9555), .Z(n9558) );
  XNOR U9461 ( .A(n9555), .B(n9375), .Z(n9557) );
  IV U9462 ( .A(p_input[780]), .Z(n9375) );
  XOR U9463 ( .A(n9559), .B(n9560), .Z(n9555) );
  AND U9464 ( .A(n9561), .B(n9562), .Z(n9560) );
  XNOR U9465 ( .A(p_input[795]), .B(n9559), .Z(n9562) );
  XNOR U9466 ( .A(n9559), .B(n9384), .Z(n9561) );
  IV U9467 ( .A(p_input[779]), .Z(n9384) );
  XOR U9468 ( .A(n9563), .B(n9564), .Z(n9559) );
  AND U9469 ( .A(n9565), .B(n9566), .Z(n9564) );
  XNOR U9470 ( .A(p_input[794]), .B(n9563), .Z(n9566) );
  XNOR U9471 ( .A(n9563), .B(n9393), .Z(n9565) );
  IV U9472 ( .A(p_input[778]), .Z(n9393) );
  XOR U9473 ( .A(n9567), .B(n9568), .Z(n9563) );
  AND U9474 ( .A(n9569), .B(n9570), .Z(n9568) );
  XNOR U9475 ( .A(p_input[793]), .B(n9567), .Z(n9570) );
  XNOR U9476 ( .A(n9567), .B(n9402), .Z(n9569) );
  IV U9477 ( .A(p_input[777]), .Z(n9402) );
  XOR U9478 ( .A(n9571), .B(n9572), .Z(n9567) );
  AND U9479 ( .A(n9573), .B(n9574), .Z(n9572) );
  XNOR U9480 ( .A(p_input[792]), .B(n9571), .Z(n9574) );
  XNOR U9481 ( .A(n9571), .B(n9411), .Z(n9573) );
  IV U9482 ( .A(p_input[776]), .Z(n9411) );
  XOR U9483 ( .A(n9575), .B(n9576), .Z(n9571) );
  AND U9484 ( .A(n9577), .B(n9578), .Z(n9576) );
  XNOR U9485 ( .A(p_input[791]), .B(n9575), .Z(n9578) );
  XNOR U9486 ( .A(n9575), .B(n9420), .Z(n9577) );
  IV U9487 ( .A(p_input[775]), .Z(n9420) );
  XOR U9488 ( .A(n9579), .B(n9580), .Z(n9575) );
  AND U9489 ( .A(n9581), .B(n9582), .Z(n9580) );
  XNOR U9490 ( .A(p_input[790]), .B(n9579), .Z(n9582) );
  XNOR U9491 ( .A(n9579), .B(n9429), .Z(n9581) );
  IV U9492 ( .A(p_input[774]), .Z(n9429) );
  XOR U9493 ( .A(n9583), .B(n9584), .Z(n9579) );
  AND U9494 ( .A(n9585), .B(n9586), .Z(n9584) );
  XNOR U9495 ( .A(p_input[789]), .B(n9583), .Z(n9586) );
  XNOR U9496 ( .A(n9583), .B(n9438), .Z(n9585) );
  IV U9497 ( .A(p_input[773]), .Z(n9438) );
  XOR U9498 ( .A(n9587), .B(n9588), .Z(n9583) );
  AND U9499 ( .A(n9589), .B(n9590), .Z(n9588) );
  XNOR U9500 ( .A(p_input[788]), .B(n9587), .Z(n9590) );
  XNOR U9501 ( .A(n9587), .B(n9447), .Z(n9589) );
  IV U9502 ( .A(p_input[772]), .Z(n9447) );
  XOR U9503 ( .A(n9591), .B(n9592), .Z(n9587) );
  AND U9504 ( .A(n9593), .B(n9594), .Z(n9592) );
  XNOR U9505 ( .A(p_input[787]), .B(n9591), .Z(n9594) );
  XNOR U9506 ( .A(n9591), .B(n9456), .Z(n9593) );
  IV U9507 ( .A(p_input[771]), .Z(n9456) );
  XOR U9508 ( .A(n9595), .B(n9596), .Z(n9591) );
  AND U9509 ( .A(n9597), .B(n9598), .Z(n9596) );
  XNOR U9510 ( .A(p_input[786]), .B(n9595), .Z(n9598) );
  XNOR U9511 ( .A(n9595), .B(n9465), .Z(n9597) );
  IV U9512 ( .A(p_input[770]), .Z(n9465) );
  XNOR U9513 ( .A(n9599), .B(n9600), .Z(n9595) );
  AND U9514 ( .A(n9601), .B(n9602), .Z(n9600) );
  XOR U9515 ( .A(p_input[785]), .B(n9599), .Z(n9602) );
  XNOR U9516 ( .A(p_input[769]), .B(n9599), .Z(n9601) );
  AND U9517 ( .A(p_input[784]), .B(n9603), .Z(n9599) );
  IV U9518 ( .A(p_input[768]), .Z(n9603) );
  XOR U9519 ( .A(n9604), .B(n9605), .Z(n7831) );
  AND U9520 ( .A(n508), .B(n9606), .Z(n9605) );
  XNOR U9521 ( .A(n9607), .B(n9604), .Z(n9606) );
  XOR U9522 ( .A(n9608), .B(n9609), .Z(n508) );
  AND U9523 ( .A(n9610), .B(n9611), .Z(n9609) );
  XNOR U9524 ( .A(n7846), .B(n9608), .Z(n9611) );
  AND U9525 ( .A(n9612), .B(n9613), .Z(n7846) );
  XNOR U9526 ( .A(n9608), .B(n7843), .Z(n9610) );
  IV U9527 ( .A(n9614), .Z(n7843) );
  AND U9528 ( .A(n9615), .B(n9616), .Z(n9614) );
  XOR U9529 ( .A(n9617), .B(n9618), .Z(n9608) );
  AND U9530 ( .A(n9619), .B(n9620), .Z(n9618) );
  XOR U9531 ( .A(n9617), .B(n7858), .Z(n9620) );
  XOR U9532 ( .A(n9621), .B(n9622), .Z(n7858) );
  AND U9533 ( .A(n442), .B(n9623), .Z(n9622) );
  XOR U9534 ( .A(n9624), .B(n9621), .Z(n9623) );
  XNOR U9535 ( .A(n7855), .B(n9617), .Z(n9619) );
  XOR U9536 ( .A(n9625), .B(n9626), .Z(n7855) );
  AND U9537 ( .A(n439), .B(n9627), .Z(n9626) );
  XOR U9538 ( .A(n9628), .B(n9625), .Z(n9627) );
  XOR U9539 ( .A(n9629), .B(n9630), .Z(n9617) );
  AND U9540 ( .A(n9631), .B(n9632), .Z(n9630) );
  XOR U9541 ( .A(n9629), .B(n7870), .Z(n9632) );
  XOR U9542 ( .A(n9633), .B(n9634), .Z(n7870) );
  AND U9543 ( .A(n442), .B(n9635), .Z(n9634) );
  XOR U9544 ( .A(n9636), .B(n9633), .Z(n9635) );
  XNOR U9545 ( .A(n7867), .B(n9629), .Z(n9631) );
  XOR U9546 ( .A(n9637), .B(n9638), .Z(n7867) );
  AND U9547 ( .A(n439), .B(n9639), .Z(n9638) );
  XOR U9548 ( .A(n9640), .B(n9637), .Z(n9639) );
  XOR U9549 ( .A(n9641), .B(n9642), .Z(n9629) );
  AND U9550 ( .A(n9643), .B(n9644), .Z(n9642) );
  XOR U9551 ( .A(n9641), .B(n7882), .Z(n9644) );
  XOR U9552 ( .A(n9645), .B(n9646), .Z(n7882) );
  AND U9553 ( .A(n442), .B(n9647), .Z(n9646) );
  XOR U9554 ( .A(n9648), .B(n9645), .Z(n9647) );
  XNOR U9555 ( .A(n7879), .B(n9641), .Z(n9643) );
  XOR U9556 ( .A(n9649), .B(n9650), .Z(n7879) );
  AND U9557 ( .A(n439), .B(n9651), .Z(n9650) );
  XOR U9558 ( .A(n9652), .B(n9649), .Z(n9651) );
  XOR U9559 ( .A(n9653), .B(n9654), .Z(n9641) );
  AND U9560 ( .A(n9655), .B(n9656), .Z(n9654) );
  XOR U9561 ( .A(n9653), .B(n7894), .Z(n9656) );
  XOR U9562 ( .A(n9657), .B(n9658), .Z(n7894) );
  AND U9563 ( .A(n442), .B(n9659), .Z(n9658) );
  XOR U9564 ( .A(n9660), .B(n9657), .Z(n9659) );
  XNOR U9565 ( .A(n7891), .B(n9653), .Z(n9655) );
  XOR U9566 ( .A(n9661), .B(n9662), .Z(n7891) );
  AND U9567 ( .A(n439), .B(n9663), .Z(n9662) );
  XOR U9568 ( .A(n9664), .B(n9661), .Z(n9663) );
  XOR U9569 ( .A(n9665), .B(n9666), .Z(n9653) );
  AND U9570 ( .A(n9667), .B(n9668), .Z(n9666) );
  XOR U9571 ( .A(n9665), .B(n7906), .Z(n9668) );
  XOR U9572 ( .A(n9669), .B(n9670), .Z(n7906) );
  AND U9573 ( .A(n442), .B(n9671), .Z(n9670) );
  XOR U9574 ( .A(n9672), .B(n9669), .Z(n9671) );
  XNOR U9575 ( .A(n7903), .B(n9665), .Z(n9667) );
  XOR U9576 ( .A(n9673), .B(n9674), .Z(n7903) );
  AND U9577 ( .A(n439), .B(n9675), .Z(n9674) );
  XOR U9578 ( .A(n9676), .B(n9673), .Z(n9675) );
  XOR U9579 ( .A(n9677), .B(n9678), .Z(n9665) );
  AND U9580 ( .A(n9679), .B(n9680), .Z(n9678) );
  XOR U9581 ( .A(n9677), .B(n7918), .Z(n9680) );
  XOR U9582 ( .A(n9681), .B(n9682), .Z(n7918) );
  AND U9583 ( .A(n442), .B(n9683), .Z(n9682) );
  XOR U9584 ( .A(n9684), .B(n9681), .Z(n9683) );
  XNOR U9585 ( .A(n7915), .B(n9677), .Z(n9679) );
  XOR U9586 ( .A(n9685), .B(n9686), .Z(n7915) );
  AND U9587 ( .A(n439), .B(n9687), .Z(n9686) );
  XOR U9588 ( .A(n9688), .B(n9685), .Z(n9687) );
  XOR U9589 ( .A(n9689), .B(n9690), .Z(n9677) );
  AND U9590 ( .A(n9691), .B(n9692), .Z(n9690) );
  XOR U9591 ( .A(n9689), .B(n7930), .Z(n9692) );
  XOR U9592 ( .A(n9693), .B(n9694), .Z(n7930) );
  AND U9593 ( .A(n442), .B(n9695), .Z(n9694) );
  XOR U9594 ( .A(n9696), .B(n9693), .Z(n9695) );
  XNOR U9595 ( .A(n7927), .B(n9689), .Z(n9691) );
  XOR U9596 ( .A(n9697), .B(n9698), .Z(n7927) );
  AND U9597 ( .A(n439), .B(n9699), .Z(n9698) );
  XOR U9598 ( .A(n9700), .B(n9697), .Z(n9699) );
  XOR U9599 ( .A(n9701), .B(n9702), .Z(n9689) );
  AND U9600 ( .A(n9703), .B(n9704), .Z(n9702) );
  XOR U9601 ( .A(n9701), .B(n7942), .Z(n9704) );
  XOR U9602 ( .A(n9705), .B(n9706), .Z(n7942) );
  AND U9603 ( .A(n442), .B(n9707), .Z(n9706) );
  XOR U9604 ( .A(n9708), .B(n9705), .Z(n9707) );
  XNOR U9605 ( .A(n7939), .B(n9701), .Z(n9703) );
  XOR U9606 ( .A(n9709), .B(n9710), .Z(n7939) );
  AND U9607 ( .A(n439), .B(n9711), .Z(n9710) );
  XOR U9608 ( .A(n9712), .B(n9709), .Z(n9711) );
  XOR U9609 ( .A(n9713), .B(n9714), .Z(n9701) );
  AND U9610 ( .A(n9715), .B(n9716), .Z(n9714) );
  XOR U9611 ( .A(n9713), .B(n7954), .Z(n9716) );
  XOR U9612 ( .A(n9717), .B(n9718), .Z(n7954) );
  AND U9613 ( .A(n442), .B(n9719), .Z(n9718) );
  XOR U9614 ( .A(n9720), .B(n9717), .Z(n9719) );
  XNOR U9615 ( .A(n7951), .B(n9713), .Z(n9715) );
  XOR U9616 ( .A(n9721), .B(n9722), .Z(n7951) );
  AND U9617 ( .A(n439), .B(n9723), .Z(n9722) );
  XOR U9618 ( .A(n9724), .B(n9721), .Z(n9723) );
  XOR U9619 ( .A(n9725), .B(n9726), .Z(n9713) );
  AND U9620 ( .A(n9727), .B(n9728), .Z(n9726) );
  XOR U9621 ( .A(n9725), .B(n7966), .Z(n9728) );
  XOR U9622 ( .A(n9729), .B(n9730), .Z(n7966) );
  AND U9623 ( .A(n442), .B(n9731), .Z(n9730) );
  XOR U9624 ( .A(n9732), .B(n9729), .Z(n9731) );
  XNOR U9625 ( .A(n7963), .B(n9725), .Z(n9727) );
  XOR U9626 ( .A(n9733), .B(n9734), .Z(n7963) );
  AND U9627 ( .A(n439), .B(n9735), .Z(n9734) );
  XOR U9628 ( .A(n9736), .B(n9733), .Z(n9735) );
  XOR U9629 ( .A(n9737), .B(n9738), .Z(n9725) );
  AND U9630 ( .A(n9739), .B(n9740), .Z(n9738) );
  XOR U9631 ( .A(n9737), .B(n7978), .Z(n9740) );
  XOR U9632 ( .A(n9741), .B(n9742), .Z(n7978) );
  AND U9633 ( .A(n442), .B(n9743), .Z(n9742) );
  XOR U9634 ( .A(n9744), .B(n9741), .Z(n9743) );
  XNOR U9635 ( .A(n7975), .B(n9737), .Z(n9739) );
  XOR U9636 ( .A(n9745), .B(n9746), .Z(n7975) );
  AND U9637 ( .A(n439), .B(n9747), .Z(n9746) );
  XOR U9638 ( .A(n9748), .B(n9745), .Z(n9747) );
  XOR U9639 ( .A(n9749), .B(n9750), .Z(n9737) );
  AND U9640 ( .A(n9751), .B(n9752), .Z(n9750) );
  XOR U9641 ( .A(n9749), .B(n7990), .Z(n9752) );
  XOR U9642 ( .A(n9753), .B(n9754), .Z(n7990) );
  AND U9643 ( .A(n442), .B(n9755), .Z(n9754) );
  XOR U9644 ( .A(n9756), .B(n9753), .Z(n9755) );
  XNOR U9645 ( .A(n7987), .B(n9749), .Z(n9751) );
  XOR U9646 ( .A(n9757), .B(n9758), .Z(n7987) );
  AND U9647 ( .A(n439), .B(n9759), .Z(n9758) );
  XOR U9648 ( .A(n9760), .B(n9757), .Z(n9759) );
  XOR U9649 ( .A(n9761), .B(n9762), .Z(n9749) );
  AND U9650 ( .A(n9763), .B(n9764), .Z(n9762) );
  XOR U9651 ( .A(n8002), .B(n9761), .Z(n9764) );
  XOR U9652 ( .A(n9765), .B(n9766), .Z(n8002) );
  AND U9653 ( .A(n442), .B(n9767), .Z(n9766) );
  XOR U9654 ( .A(n9765), .B(n9768), .Z(n9767) );
  XNOR U9655 ( .A(n9761), .B(n7999), .Z(n9763) );
  XOR U9656 ( .A(n9769), .B(n9770), .Z(n7999) );
  AND U9657 ( .A(n439), .B(n9771), .Z(n9770) );
  XOR U9658 ( .A(n9769), .B(n9772), .Z(n9771) );
  XOR U9659 ( .A(n9773), .B(n9774), .Z(n9761) );
  AND U9660 ( .A(n9775), .B(n9776), .Z(n9774) );
  XNOR U9661 ( .A(n9777), .B(n8015), .Z(n9776) );
  XOR U9662 ( .A(n9778), .B(n9779), .Z(n8015) );
  AND U9663 ( .A(n442), .B(n9780), .Z(n9779) );
  XOR U9664 ( .A(n9781), .B(n9778), .Z(n9780) );
  XNOR U9665 ( .A(n8012), .B(n9773), .Z(n9775) );
  XOR U9666 ( .A(n9782), .B(n9783), .Z(n8012) );
  AND U9667 ( .A(n439), .B(n9784), .Z(n9783) );
  XOR U9668 ( .A(n9785), .B(n9782), .Z(n9784) );
  IV U9669 ( .A(n9777), .Z(n9773) );
  AND U9670 ( .A(n9604), .B(n9607), .Z(n9777) );
  XNOR U9671 ( .A(n9786), .B(n9787), .Z(n9607) );
  AND U9672 ( .A(n442), .B(n9788), .Z(n9787) );
  XNOR U9673 ( .A(n9789), .B(n9786), .Z(n9788) );
  XOR U9674 ( .A(n9790), .B(n9791), .Z(n442) );
  AND U9675 ( .A(n9792), .B(n9793), .Z(n9791) );
  XNOR U9676 ( .A(n9612), .B(n9790), .Z(n9793) );
  AND U9677 ( .A(n9794), .B(n9795), .Z(n9612) );
  XOR U9678 ( .A(n9790), .B(n9613), .Z(n9792) );
  AND U9679 ( .A(n9796), .B(n9797), .Z(n9613) );
  XOR U9680 ( .A(n9798), .B(n9799), .Z(n9790) );
  AND U9681 ( .A(n9800), .B(n9801), .Z(n9799) );
  XOR U9682 ( .A(n9798), .B(n9624), .Z(n9801) );
  XOR U9683 ( .A(n9802), .B(n9803), .Z(n9624) );
  AND U9684 ( .A(n298), .B(n9804), .Z(n9803) );
  XOR U9685 ( .A(n9805), .B(n9802), .Z(n9804) );
  XNOR U9686 ( .A(n9621), .B(n9798), .Z(n9800) );
  XOR U9687 ( .A(n9806), .B(n9807), .Z(n9621) );
  AND U9688 ( .A(n296), .B(n9808), .Z(n9807) );
  XOR U9689 ( .A(n9809), .B(n9806), .Z(n9808) );
  XOR U9690 ( .A(n9810), .B(n9811), .Z(n9798) );
  AND U9691 ( .A(n9812), .B(n9813), .Z(n9811) );
  XOR U9692 ( .A(n9810), .B(n9636), .Z(n9813) );
  XOR U9693 ( .A(n9814), .B(n9815), .Z(n9636) );
  AND U9694 ( .A(n298), .B(n9816), .Z(n9815) );
  XOR U9695 ( .A(n9817), .B(n9814), .Z(n9816) );
  XNOR U9696 ( .A(n9633), .B(n9810), .Z(n9812) );
  XOR U9697 ( .A(n9818), .B(n9819), .Z(n9633) );
  AND U9698 ( .A(n296), .B(n9820), .Z(n9819) );
  XOR U9699 ( .A(n9821), .B(n9818), .Z(n9820) );
  XOR U9700 ( .A(n9822), .B(n9823), .Z(n9810) );
  AND U9701 ( .A(n9824), .B(n9825), .Z(n9823) );
  XOR U9702 ( .A(n9822), .B(n9648), .Z(n9825) );
  XOR U9703 ( .A(n9826), .B(n9827), .Z(n9648) );
  AND U9704 ( .A(n298), .B(n9828), .Z(n9827) );
  XOR U9705 ( .A(n9829), .B(n9826), .Z(n9828) );
  XNOR U9706 ( .A(n9645), .B(n9822), .Z(n9824) );
  XOR U9707 ( .A(n9830), .B(n9831), .Z(n9645) );
  AND U9708 ( .A(n296), .B(n9832), .Z(n9831) );
  XOR U9709 ( .A(n9833), .B(n9830), .Z(n9832) );
  XOR U9710 ( .A(n9834), .B(n9835), .Z(n9822) );
  AND U9711 ( .A(n9836), .B(n9837), .Z(n9835) );
  XOR U9712 ( .A(n9834), .B(n9660), .Z(n9837) );
  XOR U9713 ( .A(n9838), .B(n9839), .Z(n9660) );
  AND U9714 ( .A(n298), .B(n9840), .Z(n9839) );
  XOR U9715 ( .A(n9841), .B(n9838), .Z(n9840) );
  XNOR U9716 ( .A(n9657), .B(n9834), .Z(n9836) );
  XOR U9717 ( .A(n9842), .B(n9843), .Z(n9657) );
  AND U9718 ( .A(n296), .B(n9844), .Z(n9843) );
  XOR U9719 ( .A(n9845), .B(n9842), .Z(n9844) );
  XOR U9720 ( .A(n9846), .B(n9847), .Z(n9834) );
  AND U9721 ( .A(n9848), .B(n9849), .Z(n9847) );
  XOR U9722 ( .A(n9846), .B(n9672), .Z(n9849) );
  XOR U9723 ( .A(n9850), .B(n9851), .Z(n9672) );
  AND U9724 ( .A(n298), .B(n9852), .Z(n9851) );
  XOR U9725 ( .A(n9853), .B(n9850), .Z(n9852) );
  XNOR U9726 ( .A(n9669), .B(n9846), .Z(n9848) );
  XOR U9727 ( .A(n9854), .B(n9855), .Z(n9669) );
  AND U9728 ( .A(n296), .B(n9856), .Z(n9855) );
  XOR U9729 ( .A(n9857), .B(n9854), .Z(n9856) );
  XOR U9730 ( .A(n9858), .B(n9859), .Z(n9846) );
  AND U9731 ( .A(n9860), .B(n9861), .Z(n9859) );
  XOR U9732 ( .A(n9858), .B(n9684), .Z(n9861) );
  XOR U9733 ( .A(n9862), .B(n9863), .Z(n9684) );
  AND U9734 ( .A(n298), .B(n9864), .Z(n9863) );
  XOR U9735 ( .A(n9865), .B(n9862), .Z(n9864) );
  XNOR U9736 ( .A(n9681), .B(n9858), .Z(n9860) );
  XOR U9737 ( .A(n9866), .B(n9867), .Z(n9681) );
  AND U9738 ( .A(n296), .B(n9868), .Z(n9867) );
  XOR U9739 ( .A(n9869), .B(n9866), .Z(n9868) );
  XOR U9740 ( .A(n9870), .B(n9871), .Z(n9858) );
  AND U9741 ( .A(n9872), .B(n9873), .Z(n9871) );
  XOR U9742 ( .A(n9870), .B(n9696), .Z(n9873) );
  XOR U9743 ( .A(n9874), .B(n9875), .Z(n9696) );
  AND U9744 ( .A(n298), .B(n9876), .Z(n9875) );
  XOR U9745 ( .A(n9877), .B(n9874), .Z(n9876) );
  XNOR U9746 ( .A(n9693), .B(n9870), .Z(n9872) );
  XOR U9747 ( .A(n9878), .B(n9879), .Z(n9693) );
  AND U9748 ( .A(n296), .B(n9880), .Z(n9879) );
  XOR U9749 ( .A(n9881), .B(n9878), .Z(n9880) );
  XOR U9750 ( .A(n9882), .B(n9883), .Z(n9870) );
  AND U9751 ( .A(n9884), .B(n9885), .Z(n9883) );
  XOR U9752 ( .A(n9882), .B(n9708), .Z(n9885) );
  XOR U9753 ( .A(n9886), .B(n9887), .Z(n9708) );
  AND U9754 ( .A(n298), .B(n9888), .Z(n9887) );
  XOR U9755 ( .A(n9889), .B(n9886), .Z(n9888) );
  XNOR U9756 ( .A(n9705), .B(n9882), .Z(n9884) );
  XOR U9757 ( .A(n9890), .B(n9891), .Z(n9705) );
  AND U9758 ( .A(n296), .B(n9892), .Z(n9891) );
  XOR U9759 ( .A(n9893), .B(n9890), .Z(n9892) );
  XOR U9760 ( .A(n9894), .B(n9895), .Z(n9882) );
  AND U9761 ( .A(n9896), .B(n9897), .Z(n9895) );
  XOR U9762 ( .A(n9894), .B(n9720), .Z(n9897) );
  XOR U9763 ( .A(n9898), .B(n9899), .Z(n9720) );
  AND U9764 ( .A(n298), .B(n9900), .Z(n9899) );
  XOR U9765 ( .A(n9901), .B(n9898), .Z(n9900) );
  XNOR U9766 ( .A(n9717), .B(n9894), .Z(n9896) );
  XOR U9767 ( .A(n9902), .B(n9903), .Z(n9717) );
  AND U9768 ( .A(n296), .B(n9904), .Z(n9903) );
  XOR U9769 ( .A(n9905), .B(n9902), .Z(n9904) );
  XOR U9770 ( .A(n9906), .B(n9907), .Z(n9894) );
  AND U9771 ( .A(n9908), .B(n9909), .Z(n9907) );
  XOR U9772 ( .A(n9906), .B(n9732), .Z(n9909) );
  XOR U9773 ( .A(n9910), .B(n9911), .Z(n9732) );
  AND U9774 ( .A(n298), .B(n9912), .Z(n9911) );
  XOR U9775 ( .A(n9913), .B(n9910), .Z(n9912) );
  XNOR U9776 ( .A(n9729), .B(n9906), .Z(n9908) );
  XOR U9777 ( .A(n9914), .B(n9915), .Z(n9729) );
  AND U9778 ( .A(n296), .B(n9916), .Z(n9915) );
  XOR U9779 ( .A(n9917), .B(n9914), .Z(n9916) );
  XOR U9780 ( .A(n9918), .B(n9919), .Z(n9906) );
  AND U9781 ( .A(n9920), .B(n9921), .Z(n9919) );
  XOR U9782 ( .A(n9918), .B(n9744), .Z(n9921) );
  XOR U9783 ( .A(n9922), .B(n9923), .Z(n9744) );
  AND U9784 ( .A(n298), .B(n9924), .Z(n9923) );
  XOR U9785 ( .A(n9925), .B(n9922), .Z(n9924) );
  XNOR U9786 ( .A(n9741), .B(n9918), .Z(n9920) );
  XOR U9787 ( .A(n9926), .B(n9927), .Z(n9741) );
  AND U9788 ( .A(n296), .B(n9928), .Z(n9927) );
  XOR U9789 ( .A(n9929), .B(n9926), .Z(n9928) );
  XOR U9790 ( .A(n9930), .B(n9931), .Z(n9918) );
  AND U9791 ( .A(n9932), .B(n9933), .Z(n9931) );
  XOR U9792 ( .A(n9930), .B(n9756), .Z(n9933) );
  XOR U9793 ( .A(n9934), .B(n9935), .Z(n9756) );
  AND U9794 ( .A(n298), .B(n9936), .Z(n9935) );
  XOR U9795 ( .A(n9937), .B(n9934), .Z(n9936) );
  XNOR U9796 ( .A(n9753), .B(n9930), .Z(n9932) );
  XOR U9797 ( .A(n9938), .B(n9939), .Z(n9753) );
  AND U9798 ( .A(n296), .B(n9940), .Z(n9939) );
  XOR U9799 ( .A(n9941), .B(n9938), .Z(n9940) );
  XOR U9800 ( .A(n9942), .B(n9943), .Z(n9930) );
  AND U9801 ( .A(n9944), .B(n9945), .Z(n9943) );
  XOR U9802 ( .A(n9768), .B(n9942), .Z(n9945) );
  XOR U9803 ( .A(n9946), .B(n9947), .Z(n9768) );
  AND U9804 ( .A(n298), .B(n9948), .Z(n9947) );
  XOR U9805 ( .A(n9946), .B(n9949), .Z(n9948) );
  XNOR U9806 ( .A(n9942), .B(n9765), .Z(n9944) );
  XOR U9807 ( .A(n9950), .B(n9951), .Z(n9765) );
  AND U9808 ( .A(n296), .B(n9952), .Z(n9951) );
  XOR U9809 ( .A(n9950), .B(n9953), .Z(n9952) );
  XOR U9810 ( .A(n9954), .B(n9955), .Z(n9942) );
  AND U9811 ( .A(n9956), .B(n9957), .Z(n9955) );
  XNOR U9812 ( .A(n9958), .B(n9781), .Z(n9957) );
  XOR U9813 ( .A(n9959), .B(n9960), .Z(n9781) );
  AND U9814 ( .A(n298), .B(n9961), .Z(n9960) );
  XOR U9815 ( .A(n9962), .B(n9959), .Z(n9961) );
  XNOR U9816 ( .A(n9778), .B(n9954), .Z(n9956) );
  XOR U9817 ( .A(n9963), .B(n9964), .Z(n9778) );
  AND U9818 ( .A(n296), .B(n9965), .Z(n9964) );
  XOR U9819 ( .A(n9966), .B(n9963), .Z(n9965) );
  IV U9820 ( .A(n9958), .Z(n9954) );
  AND U9821 ( .A(n9786), .B(n9789), .Z(n9958) );
  XNOR U9822 ( .A(n9967), .B(n9968), .Z(n9789) );
  AND U9823 ( .A(n298), .B(n9969), .Z(n9968) );
  XNOR U9824 ( .A(n9970), .B(n9967), .Z(n9969) );
  XOR U9825 ( .A(n9971), .B(n9972), .Z(n298) );
  AND U9826 ( .A(n9973), .B(n9974), .Z(n9972) );
  XNOR U9827 ( .A(n9794), .B(n9971), .Z(n9974) );
  AND U9828 ( .A(p_input[767]), .B(p_input[751]), .Z(n9794) );
  XOR U9829 ( .A(n9971), .B(n9795), .Z(n9973) );
  AND U9830 ( .A(p_input[735]), .B(p_input[719]), .Z(n9795) );
  XOR U9831 ( .A(n9975), .B(n9976), .Z(n9971) );
  AND U9832 ( .A(n9977), .B(n9978), .Z(n9976) );
  XOR U9833 ( .A(n9975), .B(n9805), .Z(n9978) );
  XNOR U9834 ( .A(p_input[750]), .B(n9979), .Z(n9805) );
  AND U9835 ( .A(n378), .B(n9980), .Z(n9979) );
  XOR U9836 ( .A(p_input[766]), .B(p_input[750]), .Z(n9980) );
  XNOR U9837 ( .A(n9802), .B(n9975), .Z(n9977) );
  XOR U9838 ( .A(n9981), .B(n9982), .Z(n9802) );
  AND U9839 ( .A(n376), .B(n9983), .Z(n9982) );
  XOR U9840 ( .A(p_input[734]), .B(p_input[718]), .Z(n9983) );
  XOR U9841 ( .A(n9984), .B(n9985), .Z(n9975) );
  AND U9842 ( .A(n9986), .B(n9987), .Z(n9985) );
  XOR U9843 ( .A(n9984), .B(n9817), .Z(n9987) );
  XNOR U9844 ( .A(p_input[749]), .B(n9988), .Z(n9817) );
  AND U9845 ( .A(n378), .B(n9989), .Z(n9988) );
  XOR U9846 ( .A(p_input[765]), .B(p_input[749]), .Z(n9989) );
  XNOR U9847 ( .A(n9814), .B(n9984), .Z(n9986) );
  XOR U9848 ( .A(n9990), .B(n9991), .Z(n9814) );
  AND U9849 ( .A(n376), .B(n9992), .Z(n9991) );
  XOR U9850 ( .A(p_input[733]), .B(p_input[717]), .Z(n9992) );
  XOR U9851 ( .A(n9993), .B(n9994), .Z(n9984) );
  AND U9852 ( .A(n9995), .B(n9996), .Z(n9994) );
  XOR U9853 ( .A(n9993), .B(n9829), .Z(n9996) );
  XNOR U9854 ( .A(p_input[748]), .B(n9997), .Z(n9829) );
  AND U9855 ( .A(n378), .B(n9998), .Z(n9997) );
  XOR U9856 ( .A(p_input[764]), .B(p_input[748]), .Z(n9998) );
  XNOR U9857 ( .A(n9826), .B(n9993), .Z(n9995) );
  XOR U9858 ( .A(n9999), .B(n10000), .Z(n9826) );
  AND U9859 ( .A(n376), .B(n10001), .Z(n10000) );
  XOR U9860 ( .A(p_input[732]), .B(p_input[716]), .Z(n10001) );
  XOR U9861 ( .A(n10002), .B(n10003), .Z(n9993) );
  AND U9862 ( .A(n10004), .B(n10005), .Z(n10003) );
  XOR U9863 ( .A(n10002), .B(n9841), .Z(n10005) );
  XNOR U9864 ( .A(p_input[747]), .B(n10006), .Z(n9841) );
  AND U9865 ( .A(n378), .B(n10007), .Z(n10006) );
  XOR U9866 ( .A(p_input[763]), .B(p_input[747]), .Z(n10007) );
  XNOR U9867 ( .A(n9838), .B(n10002), .Z(n10004) );
  XOR U9868 ( .A(n10008), .B(n10009), .Z(n9838) );
  AND U9869 ( .A(n376), .B(n10010), .Z(n10009) );
  XOR U9870 ( .A(p_input[731]), .B(p_input[715]), .Z(n10010) );
  XOR U9871 ( .A(n10011), .B(n10012), .Z(n10002) );
  AND U9872 ( .A(n10013), .B(n10014), .Z(n10012) );
  XOR U9873 ( .A(n10011), .B(n9853), .Z(n10014) );
  XNOR U9874 ( .A(p_input[746]), .B(n10015), .Z(n9853) );
  AND U9875 ( .A(n378), .B(n10016), .Z(n10015) );
  XOR U9876 ( .A(p_input[762]), .B(p_input[746]), .Z(n10016) );
  XNOR U9877 ( .A(n9850), .B(n10011), .Z(n10013) );
  XOR U9878 ( .A(n10017), .B(n10018), .Z(n9850) );
  AND U9879 ( .A(n376), .B(n10019), .Z(n10018) );
  XOR U9880 ( .A(p_input[730]), .B(p_input[714]), .Z(n10019) );
  XOR U9881 ( .A(n10020), .B(n10021), .Z(n10011) );
  AND U9882 ( .A(n10022), .B(n10023), .Z(n10021) );
  XOR U9883 ( .A(n10020), .B(n9865), .Z(n10023) );
  XNOR U9884 ( .A(p_input[745]), .B(n10024), .Z(n9865) );
  AND U9885 ( .A(n378), .B(n10025), .Z(n10024) );
  XOR U9886 ( .A(p_input[761]), .B(p_input[745]), .Z(n10025) );
  XNOR U9887 ( .A(n9862), .B(n10020), .Z(n10022) );
  XOR U9888 ( .A(n10026), .B(n10027), .Z(n9862) );
  AND U9889 ( .A(n376), .B(n10028), .Z(n10027) );
  XOR U9890 ( .A(p_input[729]), .B(p_input[713]), .Z(n10028) );
  XOR U9891 ( .A(n10029), .B(n10030), .Z(n10020) );
  AND U9892 ( .A(n10031), .B(n10032), .Z(n10030) );
  XOR U9893 ( .A(n10029), .B(n9877), .Z(n10032) );
  XNOR U9894 ( .A(p_input[744]), .B(n10033), .Z(n9877) );
  AND U9895 ( .A(n378), .B(n10034), .Z(n10033) );
  XOR U9896 ( .A(p_input[760]), .B(p_input[744]), .Z(n10034) );
  XNOR U9897 ( .A(n9874), .B(n10029), .Z(n10031) );
  XOR U9898 ( .A(n10035), .B(n10036), .Z(n9874) );
  AND U9899 ( .A(n376), .B(n10037), .Z(n10036) );
  XOR U9900 ( .A(p_input[728]), .B(p_input[712]), .Z(n10037) );
  XOR U9901 ( .A(n10038), .B(n10039), .Z(n10029) );
  AND U9902 ( .A(n10040), .B(n10041), .Z(n10039) );
  XOR U9903 ( .A(n10038), .B(n9889), .Z(n10041) );
  XNOR U9904 ( .A(p_input[743]), .B(n10042), .Z(n9889) );
  AND U9905 ( .A(n378), .B(n10043), .Z(n10042) );
  XOR U9906 ( .A(p_input[759]), .B(p_input[743]), .Z(n10043) );
  XNOR U9907 ( .A(n9886), .B(n10038), .Z(n10040) );
  XOR U9908 ( .A(n10044), .B(n10045), .Z(n9886) );
  AND U9909 ( .A(n376), .B(n10046), .Z(n10045) );
  XOR U9910 ( .A(p_input[727]), .B(p_input[711]), .Z(n10046) );
  XOR U9911 ( .A(n10047), .B(n10048), .Z(n10038) );
  AND U9912 ( .A(n10049), .B(n10050), .Z(n10048) );
  XOR U9913 ( .A(n10047), .B(n9901), .Z(n10050) );
  XNOR U9914 ( .A(p_input[742]), .B(n10051), .Z(n9901) );
  AND U9915 ( .A(n378), .B(n10052), .Z(n10051) );
  XOR U9916 ( .A(p_input[758]), .B(p_input[742]), .Z(n10052) );
  XNOR U9917 ( .A(n9898), .B(n10047), .Z(n10049) );
  XOR U9918 ( .A(n10053), .B(n10054), .Z(n9898) );
  AND U9919 ( .A(n376), .B(n10055), .Z(n10054) );
  XOR U9920 ( .A(p_input[726]), .B(p_input[710]), .Z(n10055) );
  XOR U9921 ( .A(n10056), .B(n10057), .Z(n10047) );
  AND U9922 ( .A(n10058), .B(n10059), .Z(n10057) );
  XOR U9923 ( .A(n10056), .B(n9913), .Z(n10059) );
  XNOR U9924 ( .A(p_input[741]), .B(n10060), .Z(n9913) );
  AND U9925 ( .A(n378), .B(n10061), .Z(n10060) );
  XOR U9926 ( .A(p_input[757]), .B(p_input[741]), .Z(n10061) );
  XNOR U9927 ( .A(n9910), .B(n10056), .Z(n10058) );
  XOR U9928 ( .A(n10062), .B(n10063), .Z(n9910) );
  AND U9929 ( .A(n376), .B(n10064), .Z(n10063) );
  XOR U9930 ( .A(p_input[725]), .B(p_input[709]), .Z(n10064) );
  XOR U9931 ( .A(n10065), .B(n10066), .Z(n10056) );
  AND U9932 ( .A(n10067), .B(n10068), .Z(n10066) );
  XOR U9933 ( .A(n10065), .B(n9925), .Z(n10068) );
  XNOR U9934 ( .A(p_input[740]), .B(n10069), .Z(n9925) );
  AND U9935 ( .A(n378), .B(n10070), .Z(n10069) );
  XOR U9936 ( .A(p_input[756]), .B(p_input[740]), .Z(n10070) );
  XNOR U9937 ( .A(n9922), .B(n10065), .Z(n10067) );
  XOR U9938 ( .A(n10071), .B(n10072), .Z(n9922) );
  AND U9939 ( .A(n376), .B(n10073), .Z(n10072) );
  XOR U9940 ( .A(p_input[724]), .B(p_input[708]), .Z(n10073) );
  XOR U9941 ( .A(n10074), .B(n10075), .Z(n10065) );
  AND U9942 ( .A(n10076), .B(n10077), .Z(n10075) );
  XOR U9943 ( .A(n10074), .B(n9937), .Z(n10077) );
  XNOR U9944 ( .A(p_input[739]), .B(n10078), .Z(n9937) );
  AND U9945 ( .A(n378), .B(n10079), .Z(n10078) );
  XOR U9946 ( .A(p_input[755]), .B(p_input[739]), .Z(n10079) );
  XNOR U9947 ( .A(n9934), .B(n10074), .Z(n10076) );
  XOR U9948 ( .A(n10080), .B(n10081), .Z(n9934) );
  AND U9949 ( .A(n376), .B(n10082), .Z(n10081) );
  XOR U9950 ( .A(p_input[723]), .B(p_input[707]), .Z(n10082) );
  XOR U9951 ( .A(n10083), .B(n10084), .Z(n10074) );
  AND U9952 ( .A(n10085), .B(n10086), .Z(n10084) );
  XOR U9953 ( .A(n9949), .B(n10083), .Z(n10086) );
  XNOR U9954 ( .A(p_input[738]), .B(n10087), .Z(n9949) );
  AND U9955 ( .A(n378), .B(n10088), .Z(n10087) );
  XOR U9956 ( .A(p_input[754]), .B(p_input[738]), .Z(n10088) );
  XNOR U9957 ( .A(n10083), .B(n9946), .Z(n10085) );
  XOR U9958 ( .A(n10089), .B(n10090), .Z(n9946) );
  AND U9959 ( .A(n376), .B(n10091), .Z(n10090) );
  XOR U9960 ( .A(p_input[722]), .B(p_input[706]), .Z(n10091) );
  XOR U9961 ( .A(n10092), .B(n10093), .Z(n10083) );
  AND U9962 ( .A(n10094), .B(n10095), .Z(n10093) );
  XNOR U9963 ( .A(n10096), .B(n9962), .Z(n10095) );
  XNOR U9964 ( .A(p_input[737]), .B(n10097), .Z(n9962) );
  AND U9965 ( .A(n378), .B(n10098), .Z(n10097) );
  XNOR U9966 ( .A(p_input[753]), .B(n10099), .Z(n10098) );
  IV U9967 ( .A(p_input[737]), .Z(n10099) );
  XNOR U9968 ( .A(n9959), .B(n10092), .Z(n10094) );
  XNOR U9969 ( .A(p_input[705]), .B(n10100), .Z(n9959) );
  AND U9970 ( .A(n376), .B(n10101), .Z(n10100) );
  XOR U9971 ( .A(p_input[721]), .B(p_input[705]), .Z(n10101) );
  IV U9972 ( .A(n10096), .Z(n10092) );
  AND U9973 ( .A(n9967), .B(n9970), .Z(n10096) );
  XOR U9974 ( .A(p_input[736]), .B(n10102), .Z(n9970) );
  AND U9975 ( .A(n378), .B(n10103), .Z(n10102) );
  XOR U9976 ( .A(p_input[752]), .B(p_input[736]), .Z(n10103) );
  XOR U9977 ( .A(n10104), .B(n10105), .Z(n378) );
  AND U9978 ( .A(n10106), .B(n10107), .Z(n10105) );
  XNOR U9979 ( .A(p_input[767]), .B(n10104), .Z(n10107) );
  XOR U9980 ( .A(n10104), .B(p_input[751]), .Z(n10106) );
  XOR U9981 ( .A(n10108), .B(n10109), .Z(n10104) );
  AND U9982 ( .A(n10110), .B(n10111), .Z(n10109) );
  XNOR U9983 ( .A(p_input[766]), .B(n10108), .Z(n10111) );
  XOR U9984 ( .A(n10108), .B(p_input[750]), .Z(n10110) );
  XOR U9985 ( .A(n10112), .B(n10113), .Z(n10108) );
  AND U9986 ( .A(n10114), .B(n10115), .Z(n10113) );
  XNOR U9987 ( .A(p_input[765]), .B(n10112), .Z(n10115) );
  XOR U9988 ( .A(n10112), .B(p_input[749]), .Z(n10114) );
  XOR U9989 ( .A(n10116), .B(n10117), .Z(n10112) );
  AND U9990 ( .A(n10118), .B(n10119), .Z(n10117) );
  XNOR U9991 ( .A(p_input[764]), .B(n10116), .Z(n10119) );
  XOR U9992 ( .A(n10116), .B(p_input[748]), .Z(n10118) );
  XOR U9993 ( .A(n10120), .B(n10121), .Z(n10116) );
  AND U9994 ( .A(n10122), .B(n10123), .Z(n10121) );
  XNOR U9995 ( .A(p_input[763]), .B(n10120), .Z(n10123) );
  XOR U9996 ( .A(n10120), .B(p_input[747]), .Z(n10122) );
  XOR U9997 ( .A(n10124), .B(n10125), .Z(n10120) );
  AND U9998 ( .A(n10126), .B(n10127), .Z(n10125) );
  XNOR U9999 ( .A(p_input[762]), .B(n10124), .Z(n10127) );
  XOR U10000 ( .A(n10124), .B(p_input[746]), .Z(n10126) );
  XOR U10001 ( .A(n10128), .B(n10129), .Z(n10124) );
  AND U10002 ( .A(n10130), .B(n10131), .Z(n10129) );
  XNOR U10003 ( .A(p_input[761]), .B(n10128), .Z(n10131) );
  XOR U10004 ( .A(n10128), .B(p_input[745]), .Z(n10130) );
  XOR U10005 ( .A(n10132), .B(n10133), .Z(n10128) );
  AND U10006 ( .A(n10134), .B(n10135), .Z(n10133) );
  XNOR U10007 ( .A(p_input[760]), .B(n10132), .Z(n10135) );
  XOR U10008 ( .A(n10132), .B(p_input[744]), .Z(n10134) );
  XOR U10009 ( .A(n10136), .B(n10137), .Z(n10132) );
  AND U10010 ( .A(n10138), .B(n10139), .Z(n10137) );
  XNOR U10011 ( .A(p_input[759]), .B(n10136), .Z(n10139) );
  XOR U10012 ( .A(n10136), .B(p_input[743]), .Z(n10138) );
  XOR U10013 ( .A(n10140), .B(n10141), .Z(n10136) );
  AND U10014 ( .A(n10142), .B(n10143), .Z(n10141) );
  XNOR U10015 ( .A(p_input[758]), .B(n10140), .Z(n10143) );
  XOR U10016 ( .A(n10140), .B(p_input[742]), .Z(n10142) );
  XOR U10017 ( .A(n10144), .B(n10145), .Z(n10140) );
  AND U10018 ( .A(n10146), .B(n10147), .Z(n10145) );
  XNOR U10019 ( .A(p_input[757]), .B(n10144), .Z(n10147) );
  XOR U10020 ( .A(n10144), .B(p_input[741]), .Z(n10146) );
  XOR U10021 ( .A(n10148), .B(n10149), .Z(n10144) );
  AND U10022 ( .A(n10150), .B(n10151), .Z(n10149) );
  XNOR U10023 ( .A(p_input[756]), .B(n10148), .Z(n10151) );
  XOR U10024 ( .A(n10148), .B(p_input[740]), .Z(n10150) );
  XOR U10025 ( .A(n10152), .B(n10153), .Z(n10148) );
  AND U10026 ( .A(n10154), .B(n10155), .Z(n10153) );
  XNOR U10027 ( .A(p_input[755]), .B(n10152), .Z(n10155) );
  XOR U10028 ( .A(n10152), .B(p_input[739]), .Z(n10154) );
  XOR U10029 ( .A(n10156), .B(n10157), .Z(n10152) );
  AND U10030 ( .A(n10158), .B(n10159), .Z(n10157) );
  XNOR U10031 ( .A(p_input[754]), .B(n10156), .Z(n10159) );
  XOR U10032 ( .A(n10156), .B(p_input[738]), .Z(n10158) );
  XNOR U10033 ( .A(n10160), .B(n10161), .Z(n10156) );
  AND U10034 ( .A(n10162), .B(n10163), .Z(n10161) );
  XOR U10035 ( .A(p_input[753]), .B(n10160), .Z(n10163) );
  XNOR U10036 ( .A(p_input[737]), .B(n10160), .Z(n10162) );
  AND U10037 ( .A(p_input[752]), .B(n10164), .Z(n10160) );
  IV U10038 ( .A(p_input[736]), .Z(n10164) );
  XNOR U10039 ( .A(p_input[704]), .B(n10165), .Z(n9967) );
  AND U10040 ( .A(n376), .B(n10166), .Z(n10165) );
  XOR U10041 ( .A(p_input[720]), .B(p_input[704]), .Z(n10166) );
  XOR U10042 ( .A(n10167), .B(n10168), .Z(n376) );
  AND U10043 ( .A(n10169), .B(n10170), .Z(n10168) );
  XNOR U10044 ( .A(p_input[735]), .B(n10167), .Z(n10170) );
  XOR U10045 ( .A(n10167), .B(p_input[719]), .Z(n10169) );
  XOR U10046 ( .A(n10171), .B(n10172), .Z(n10167) );
  AND U10047 ( .A(n10173), .B(n10174), .Z(n10172) );
  XNOR U10048 ( .A(p_input[734]), .B(n10171), .Z(n10174) );
  XNOR U10049 ( .A(n10171), .B(n9981), .Z(n10173) );
  IV U10050 ( .A(p_input[718]), .Z(n9981) );
  XOR U10051 ( .A(n10175), .B(n10176), .Z(n10171) );
  AND U10052 ( .A(n10177), .B(n10178), .Z(n10176) );
  XNOR U10053 ( .A(p_input[733]), .B(n10175), .Z(n10178) );
  XNOR U10054 ( .A(n10175), .B(n9990), .Z(n10177) );
  IV U10055 ( .A(p_input[717]), .Z(n9990) );
  XOR U10056 ( .A(n10179), .B(n10180), .Z(n10175) );
  AND U10057 ( .A(n10181), .B(n10182), .Z(n10180) );
  XNOR U10058 ( .A(p_input[732]), .B(n10179), .Z(n10182) );
  XNOR U10059 ( .A(n10179), .B(n9999), .Z(n10181) );
  IV U10060 ( .A(p_input[716]), .Z(n9999) );
  XOR U10061 ( .A(n10183), .B(n10184), .Z(n10179) );
  AND U10062 ( .A(n10185), .B(n10186), .Z(n10184) );
  XNOR U10063 ( .A(p_input[731]), .B(n10183), .Z(n10186) );
  XNOR U10064 ( .A(n10183), .B(n10008), .Z(n10185) );
  IV U10065 ( .A(p_input[715]), .Z(n10008) );
  XOR U10066 ( .A(n10187), .B(n10188), .Z(n10183) );
  AND U10067 ( .A(n10189), .B(n10190), .Z(n10188) );
  XNOR U10068 ( .A(p_input[730]), .B(n10187), .Z(n10190) );
  XNOR U10069 ( .A(n10187), .B(n10017), .Z(n10189) );
  IV U10070 ( .A(p_input[714]), .Z(n10017) );
  XOR U10071 ( .A(n10191), .B(n10192), .Z(n10187) );
  AND U10072 ( .A(n10193), .B(n10194), .Z(n10192) );
  XNOR U10073 ( .A(p_input[729]), .B(n10191), .Z(n10194) );
  XNOR U10074 ( .A(n10191), .B(n10026), .Z(n10193) );
  IV U10075 ( .A(p_input[713]), .Z(n10026) );
  XOR U10076 ( .A(n10195), .B(n10196), .Z(n10191) );
  AND U10077 ( .A(n10197), .B(n10198), .Z(n10196) );
  XNOR U10078 ( .A(p_input[728]), .B(n10195), .Z(n10198) );
  XNOR U10079 ( .A(n10195), .B(n10035), .Z(n10197) );
  IV U10080 ( .A(p_input[712]), .Z(n10035) );
  XOR U10081 ( .A(n10199), .B(n10200), .Z(n10195) );
  AND U10082 ( .A(n10201), .B(n10202), .Z(n10200) );
  XNOR U10083 ( .A(p_input[727]), .B(n10199), .Z(n10202) );
  XNOR U10084 ( .A(n10199), .B(n10044), .Z(n10201) );
  IV U10085 ( .A(p_input[711]), .Z(n10044) );
  XOR U10086 ( .A(n10203), .B(n10204), .Z(n10199) );
  AND U10087 ( .A(n10205), .B(n10206), .Z(n10204) );
  XNOR U10088 ( .A(p_input[726]), .B(n10203), .Z(n10206) );
  XNOR U10089 ( .A(n10203), .B(n10053), .Z(n10205) );
  IV U10090 ( .A(p_input[710]), .Z(n10053) );
  XOR U10091 ( .A(n10207), .B(n10208), .Z(n10203) );
  AND U10092 ( .A(n10209), .B(n10210), .Z(n10208) );
  XNOR U10093 ( .A(p_input[725]), .B(n10207), .Z(n10210) );
  XNOR U10094 ( .A(n10207), .B(n10062), .Z(n10209) );
  IV U10095 ( .A(p_input[709]), .Z(n10062) );
  XOR U10096 ( .A(n10211), .B(n10212), .Z(n10207) );
  AND U10097 ( .A(n10213), .B(n10214), .Z(n10212) );
  XNOR U10098 ( .A(p_input[724]), .B(n10211), .Z(n10214) );
  XNOR U10099 ( .A(n10211), .B(n10071), .Z(n10213) );
  IV U10100 ( .A(p_input[708]), .Z(n10071) );
  XOR U10101 ( .A(n10215), .B(n10216), .Z(n10211) );
  AND U10102 ( .A(n10217), .B(n10218), .Z(n10216) );
  XNOR U10103 ( .A(p_input[723]), .B(n10215), .Z(n10218) );
  XNOR U10104 ( .A(n10215), .B(n10080), .Z(n10217) );
  IV U10105 ( .A(p_input[707]), .Z(n10080) );
  XOR U10106 ( .A(n10219), .B(n10220), .Z(n10215) );
  AND U10107 ( .A(n10221), .B(n10222), .Z(n10220) );
  XNOR U10108 ( .A(p_input[722]), .B(n10219), .Z(n10222) );
  XNOR U10109 ( .A(n10219), .B(n10089), .Z(n10221) );
  IV U10110 ( .A(p_input[706]), .Z(n10089) );
  XNOR U10111 ( .A(n10223), .B(n10224), .Z(n10219) );
  AND U10112 ( .A(n10225), .B(n10226), .Z(n10224) );
  XOR U10113 ( .A(p_input[721]), .B(n10223), .Z(n10226) );
  XNOR U10114 ( .A(p_input[705]), .B(n10223), .Z(n10225) );
  AND U10115 ( .A(p_input[720]), .B(n10227), .Z(n10223) );
  IV U10116 ( .A(p_input[704]), .Z(n10227) );
  XOR U10117 ( .A(n10228), .B(n10229), .Z(n9786) );
  AND U10118 ( .A(n296), .B(n10230), .Z(n10229) );
  XNOR U10119 ( .A(n10231), .B(n10228), .Z(n10230) );
  XOR U10120 ( .A(n10232), .B(n10233), .Z(n296) );
  AND U10121 ( .A(n10234), .B(n10235), .Z(n10233) );
  XNOR U10122 ( .A(n9796), .B(n10232), .Z(n10235) );
  AND U10123 ( .A(p_input[703]), .B(p_input[687]), .Z(n9796) );
  XOR U10124 ( .A(n10232), .B(n9797), .Z(n10234) );
  AND U10125 ( .A(p_input[671]), .B(p_input[655]), .Z(n9797) );
  XOR U10126 ( .A(n10236), .B(n10237), .Z(n10232) );
  AND U10127 ( .A(n10238), .B(n10239), .Z(n10237) );
  XOR U10128 ( .A(n10236), .B(n9809), .Z(n10239) );
  XNOR U10129 ( .A(p_input[686]), .B(n10240), .Z(n9809) );
  AND U10130 ( .A(n382), .B(n10241), .Z(n10240) );
  XOR U10131 ( .A(p_input[702]), .B(p_input[686]), .Z(n10241) );
  XNOR U10132 ( .A(n9806), .B(n10236), .Z(n10238) );
  XOR U10133 ( .A(n10242), .B(n10243), .Z(n9806) );
  AND U10134 ( .A(n379), .B(n10244), .Z(n10243) );
  XOR U10135 ( .A(p_input[670]), .B(p_input[654]), .Z(n10244) );
  XOR U10136 ( .A(n10245), .B(n10246), .Z(n10236) );
  AND U10137 ( .A(n10247), .B(n10248), .Z(n10246) );
  XOR U10138 ( .A(n10245), .B(n9821), .Z(n10248) );
  XNOR U10139 ( .A(p_input[685]), .B(n10249), .Z(n9821) );
  AND U10140 ( .A(n382), .B(n10250), .Z(n10249) );
  XOR U10141 ( .A(p_input[701]), .B(p_input[685]), .Z(n10250) );
  XNOR U10142 ( .A(n9818), .B(n10245), .Z(n10247) );
  XOR U10143 ( .A(n10251), .B(n10252), .Z(n9818) );
  AND U10144 ( .A(n379), .B(n10253), .Z(n10252) );
  XOR U10145 ( .A(p_input[669]), .B(p_input[653]), .Z(n10253) );
  XOR U10146 ( .A(n10254), .B(n10255), .Z(n10245) );
  AND U10147 ( .A(n10256), .B(n10257), .Z(n10255) );
  XOR U10148 ( .A(n10254), .B(n9833), .Z(n10257) );
  XNOR U10149 ( .A(p_input[684]), .B(n10258), .Z(n9833) );
  AND U10150 ( .A(n382), .B(n10259), .Z(n10258) );
  XOR U10151 ( .A(p_input[700]), .B(p_input[684]), .Z(n10259) );
  XNOR U10152 ( .A(n9830), .B(n10254), .Z(n10256) );
  XOR U10153 ( .A(n10260), .B(n10261), .Z(n9830) );
  AND U10154 ( .A(n379), .B(n10262), .Z(n10261) );
  XOR U10155 ( .A(p_input[668]), .B(p_input[652]), .Z(n10262) );
  XOR U10156 ( .A(n10263), .B(n10264), .Z(n10254) );
  AND U10157 ( .A(n10265), .B(n10266), .Z(n10264) );
  XOR U10158 ( .A(n10263), .B(n9845), .Z(n10266) );
  XNOR U10159 ( .A(p_input[683]), .B(n10267), .Z(n9845) );
  AND U10160 ( .A(n382), .B(n10268), .Z(n10267) );
  XOR U10161 ( .A(p_input[699]), .B(p_input[683]), .Z(n10268) );
  XNOR U10162 ( .A(n9842), .B(n10263), .Z(n10265) );
  XOR U10163 ( .A(n10269), .B(n10270), .Z(n9842) );
  AND U10164 ( .A(n379), .B(n10271), .Z(n10270) );
  XOR U10165 ( .A(p_input[667]), .B(p_input[651]), .Z(n10271) );
  XOR U10166 ( .A(n10272), .B(n10273), .Z(n10263) );
  AND U10167 ( .A(n10274), .B(n10275), .Z(n10273) );
  XOR U10168 ( .A(n10272), .B(n9857), .Z(n10275) );
  XNOR U10169 ( .A(p_input[682]), .B(n10276), .Z(n9857) );
  AND U10170 ( .A(n382), .B(n10277), .Z(n10276) );
  XOR U10171 ( .A(p_input[698]), .B(p_input[682]), .Z(n10277) );
  XNOR U10172 ( .A(n9854), .B(n10272), .Z(n10274) );
  XOR U10173 ( .A(n10278), .B(n10279), .Z(n9854) );
  AND U10174 ( .A(n379), .B(n10280), .Z(n10279) );
  XOR U10175 ( .A(p_input[666]), .B(p_input[650]), .Z(n10280) );
  XOR U10176 ( .A(n10281), .B(n10282), .Z(n10272) );
  AND U10177 ( .A(n10283), .B(n10284), .Z(n10282) );
  XOR U10178 ( .A(n10281), .B(n9869), .Z(n10284) );
  XNOR U10179 ( .A(p_input[681]), .B(n10285), .Z(n9869) );
  AND U10180 ( .A(n382), .B(n10286), .Z(n10285) );
  XOR U10181 ( .A(p_input[697]), .B(p_input[681]), .Z(n10286) );
  XNOR U10182 ( .A(n9866), .B(n10281), .Z(n10283) );
  XOR U10183 ( .A(n10287), .B(n10288), .Z(n9866) );
  AND U10184 ( .A(n379), .B(n10289), .Z(n10288) );
  XOR U10185 ( .A(p_input[665]), .B(p_input[649]), .Z(n10289) );
  XOR U10186 ( .A(n10290), .B(n10291), .Z(n10281) );
  AND U10187 ( .A(n10292), .B(n10293), .Z(n10291) );
  XOR U10188 ( .A(n10290), .B(n9881), .Z(n10293) );
  XNOR U10189 ( .A(p_input[680]), .B(n10294), .Z(n9881) );
  AND U10190 ( .A(n382), .B(n10295), .Z(n10294) );
  XOR U10191 ( .A(p_input[696]), .B(p_input[680]), .Z(n10295) );
  XNOR U10192 ( .A(n9878), .B(n10290), .Z(n10292) );
  XOR U10193 ( .A(n10296), .B(n10297), .Z(n9878) );
  AND U10194 ( .A(n379), .B(n10298), .Z(n10297) );
  XOR U10195 ( .A(p_input[664]), .B(p_input[648]), .Z(n10298) );
  XOR U10196 ( .A(n10299), .B(n10300), .Z(n10290) );
  AND U10197 ( .A(n10301), .B(n10302), .Z(n10300) );
  XOR U10198 ( .A(n10299), .B(n9893), .Z(n10302) );
  XNOR U10199 ( .A(p_input[679]), .B(n10303), .Z(n9893) );
  AND U10200 ( .A(n382), .B(n10304), .Z(n10303) );
  XOR U10201 ( .A(p_input[695]), .B(p_input[679]), .Z(n10304) );
  XNOR U10202 ( .A(n9890), .B(n10299), .Z(n10301) );
  XOR U10203 ( .A(n10305), .B(n10306), .Z(n9890) );
  AND U10204 ( .A(n379), .B(n10307), .Z(n10306) );
  XOR U10205 ( .A(p_input[663]), .B(p_input[647]), .Z(n10307) );
  XOR U10206 ( .A(n10308), .B(n10309), .Z(n10299) );
  AND U10207 ( .A(n10310), .B(n10311), .Z(n10309) );
  XOR U10208 ( .A(n10308), .B(n9905), .Z(n10311) );
  XNOR U10209 ( .A(p_input[678]), .B(n10312), .Z(n9905) );
  AND U10210 ( .A(n382), .B(n10313), .Z(n10312) );
  XOR U10211 ( .A(p_input[694]), .B(p_input[678]), .Z(n10313) );
  XNOR U10212 ( .A(n9902), .B(n10308), .Z(n10310) );
  XOR U10213 ( .A(n10314), .B(n10315), .Z(n9902) );
  AND U10214 ( .A(n379), .B(n10316), .Z(n10315) );
  XOR U10215 ( .A(p_input[662]), .B(p_input[646]), .Z(n10316) );
  XOR U10216 ( .A(n10317), .B(n10318), .Z(n10308) );
  AND U10217 ( .A(n10319), .B(n10320), .Z(n10318) );
  XOR U10218 ( .A(n10317), .B(n9917), .Z(n10320) );
  XNOR U10219 ( .A(p_input[677]), .B(n10321), .Z(n9917) );
  AND U10220 ( .A(n382), .B(n10322), .Z(n10321) );
  XOR U10221 ( .A(p_input[693]), .B(p_input[677]), .Z(n10322) );
  XNOR U10222 ( .A(n9914), .B(n10317), .Z(n10319) );
  XOR U10223 ( .A(n10323), .B(n10324), .Z(n9914) );
  AND U10224 ( .A(n379), .B(n10325), .Z(n10324) );
  XOR U10225 ( .A(p_input[661]), .B(p_input[645]), .Z(n10325) );
  XOR U10226 ( .A(n10326), .B(n10327), .Z(n10317) );
  AND U10227 ( .A(n10328), .B(n10329), .Z(n10327) );
  XOR U10228 ( .A(n10326), .B(n9929), .Z(n10329) );
  XNOR U10229 ( .A(p_input[676]), .B(n10330), .Z(n9929) );
  AND U10230 ( .A(n382), .B(n10331), .Z(n10330) );
  XOR U10231 ( .A(p_input[692]), .B(p_input[676]), .Z(n10331) );
  XNOR U10232 ( .A(n9926), .B(n10326), .Z(n10328) );
  XOR U10233 ( .A(n10332), .B(n10333), .Z(n9926) );
  AND U10234 ( .A(n379), .B(n10334), .Z(n10333) );
  XOR U10235 ( .A(p_input[660]), .B(p_input[644]), .Z(n10334) );
  XOR U10236 ( .A(n10335), .B(n10336), .Z(n10326) );
  AND U10237 ( .A(n10337), .B(n10338), .Z(n10336) );
  XOR U10238 ( .A(n10335), .B(n9941), .Z(n10338) );
  XNOR U10239 ( .A(p_input[675]), .B(n10339), .Z(n9941) );
  AND U10240 ( .A(n382), .B(n10340), .Z(n10339) );
  XOR U10241 ( .A(p_input[691]), .B(p_input[675]), .Z(n10340) );
  XNOR U10242 ( .A(n9938), .B(n10335), .Z(n10337) );
  XOR U10243 ( .A(n10341), .B(n10342), .Z(n9938) );
  AND U10244 ( .A(n379), .B(n10343), .Z(n10342) );
  XOR U10245 ( .A(p_input[659]), .B(p_input[643]), .Z(n10343) );
  XOR U10246 ( .A(n10344), .B(n10345), .Z(n10335) );
  AND U10247 ( .A(n10346), .B(n10347), .Z(n10345) );
  XOR U10248 ( .A(n9953), .B(n10344), .Z(n10347) );
  XNOR U10249 ( .A(p_input[674]), .B(n10348), .Z(n9953) );
  AND U10250 ( .A(n382), .B(n10349), .Z(n10348) );
  XOR U10251 ( .A(p_input[690]), .B(p_input[674]), .Z(n10349) );
  XNOR U10252 ( .A(n10344), .B(n9950), .Z(n10346) );
  XOR U10253 ( .A(n10350), .B(n10351), .Z(n9950) );
  AND U10254 ( .A(n379), .B(n10352), .Z(n10351) );
  XOR U10255 ( .A(p_input[658]), .B(p_input[642]), .Z(n10352) );
  XOR U10256 ( .A(n10353), .B(n10354), .Z(n10344) );
  AND U10257 ( .A(n10355), .B(n10356), .Z(n10354) );
  XNOR U10258 ( .A(n10357), .B(n9966), .Z(n10356) );
  XNOR U10259 ( .A(p_input[673]), .B(n10358), .Z(n9966) );
  AND U10260 ( .A(n382), .B(n10359), .Z(n10358) );
  XNOR U10261 ( .A(p_input[689]), .B(n10360), .Z(n10359) );
  IV U10262 ( .A(p_input[673]), .Z(n10360) );
  XNOR U10263 ( .A(n9963), .B(n10353), .Z(n10355) );
  XNOR U10264 ( .A(p_input[641]), .B(n10361), .Z(n9963) );
  AND U10265 ( .A(n379), .B(n10362), .Z(n10361) );
  XOR U10266 ( .A(p_input[657]), .B(p_input[641]), .Z(n10362) );
  IV U10267 ( .A(n10357), .Z(n10353) );
  AND U10268 ( .A(n10228), .B(n10231), .Z(n10357) );
  XOR U10269 ( .A(p_input[672]), .B(n10363), .Z(n10231) );
  AND U10270 ( .A(n382), .B(n10364), .Z(n10363) );
  XOR U10271 ( .A(p_input[688]), .B(p_input[672]), .Z(n10364) );
  XOR U10272 ( .A(n10365), .B(n10366), .Z(n382) );
  AND U10273 ( .A(n10367), .B(n10368), .Z(n10366) );
  XNOR U10274 ( .A(p_input[703]), .B(n10365), .Z(n10368) );
  XOR U10275 ( .A(n10365), .B(p_input[687]), .Z(n10367) );
  XOR U10276 ( .A(n10369), .B(n10370), .Z(n10365) );
  AND U10277 ( .A(n10371), .B(n10372), .Z(n10370) );
  XNOR U10278 ( .A(p_input[702]), .B(n10369), .Z(n10372) );
  XOR U10279 ( .A(n10369), .B(p_input[686]), .Z(n10371) );
  XOR U10280 ( .A(n10373), .B(n10374), .Z(n10369) );
  AND U10281 ( .A(n10375), .B(n10376), .Z(n10374) );
  XNOR U10282 ( .A(p_input[701]), .B(n10373), .Z(n10376) );
  XOR U10283 ( .A(n10373), .B(p_input[685]), .Z(n10375) );
  XOR U10284 ( .A(n10377), .B(n10378), .Z(n10373) );
  AND U10285 ( .A(n10379), .B(n10380), .Z(n10378) );
  XNOR U10286 ( .A(p_input[700]), .B(n10377), .Z(n10380) );
  XOR U10287 ( .A(n10377), .B(p_input[684]), .Z(n10379) );
  XOR U10288 ( .A(n10381), .B(n10382), .Z(n10377) );
  AND U10289 ( .A(n10383), .B(n10384), .Z(n10382) );
  XNOR U10290 ( .A(p_input[699]), .B(n10381), .Z(n10384) );
  XOR U10291 ( .A(n10381), .B(p_input[683]), .Z(n10383) );
  XOR U10292 ( .A(n10385), .B(n10386), .Z(n10381) );
  AND U10293 ( .A(n10387), .B(n10388), .Z(n10386) );
  XNOR U10294 ( .A(p_input[698]), .B(n10385), .Z(n10388) );
  XOR U10295 ( .A(n10385), .B(p_input[682]), .Z(n10387) );
  XOR U10296 ( .A(n10389), .B(n10390), .Z(n10385) );
  AND U10297 ( .A(n10391), .B(n10392), .Z(n10390) );
  XNOR U10298 ( .A(p_input[697]), .B(n10389), .Z(n10392) );
  XOR U10299 ( .A(n10389), .B(p_input[681]), .Z(n10391) );
  XOR U10300 ( .A(n10393), .B(n10394), .Z(n10389) );
  AND U10301 ( .A(n10395), .B(n10396), .Z(n10394) );
  XNOR U10302 ( .A(p_input[696]), .B(n10393), .Z(n10396) );
  XOR U10303 ( .A(n10393), .B(p_input[680]), .Z(n10395) );
  XOR U10304 ( .A(n10397), .B(n10398), .Z(n10393) );
  AND U10305 ( .A(n10399), .B(n10400), .Z(n10398) );
  XNOR U10306 ( .A(p_input[695]), .B(n10397), .Z(n10400) );
  XOR U10307 ( .A(n10397), .B(p_input[679]), .Z(n10399) );
  XOR U10308 ( .A(n10401), .B(n10402), .Z(n10397) );
  AND U10309 ( .A(n10403), .B(n10404), .Z(n10402) );
  XNOR U10310 ( .A(p_input[694]), .B(n10401), .Z(n10404) );
  XOR U10311 ( .A(n10401), .B(p_input[678]), .Z(n10403) );
  XOR U10312 ( .A(n10405), .B(n10406), .Z(n10401) );
  AND U10313 ( .A(n10407), .B(n10408), .Z(n10406) );
  XNOR U10314 ( .A(p_input[693]), .B(n10405), .Z(n10408) );
  XOR U10315 ( .A(n10405), .B(p_input[677]), .Z(n10407) );
  XOR U10316 ( .A(n10409), .B(n10410), .Z(n10405) );
  AND U10317 ( .A(n10411), .B(n10412), .Z(n10410) );
  XNOR U10318 ( .A(p_input[692]), .B(n10409), .Z(n10412) );
  XOR U10319 ( .A(n10409), .B(p_input[676]), .Z(n10411) );
  XOR U10320 ( .A(n10413), .B(n10414), .Z(n10409) );
  AND U10321 ( .A(n10415), .B(n10416), .Z(n10414) );
  XNOR U10322 ( .A(p_input[691]), .B(n10413), .Z(n10416) );
  XOR U10323 ( .A(n10413), .B(p_input[675]), .Z(n10415) );
  XOR U10324 ( .A(n10417), .B(n10418), .Z(n10413) );
  AND U10325 ( .A(n10419), .B(n10420), .Z(n10418) );
  XNOR U10326 ( .A(p_input[690]), .B(n10417), .Z(n10420) );
  XOR U10327 ( .A(n10417), .B(p_input[674]), .Z(n10419) );
  XNOR U10328 ( .A(n10421), .B(n10422), .Z(n10417) );
  AND U10329 ( .A(n10423), .B(n10424), .Z(n10422) );
  XOR U10330 ( .A(p_input[689]), .B(n10421), .Z(n10424) );
  XNOR U10331 ( .A(p_input[673]), .B(n10421), .Z(n10423) );
  AND U10332 ( .A(p_input[688]), .B(n10425), .Z(n10421) );
  IV U10333 ( .A(p_input[672]), .Z(n10425) );
  XNOR U10334 ( .A(p_input[640]), .B(n10426), .Z(n10228) );
  AND U10335 ( .A(n379), .B(n10427), .Z(n10426) );
  XOR U10336 ( .A(p_input[656]), .B(p_input[640]), .Z(n10427) );
  XOR U10337 ( .A(n10428), .B(n10429), .Z(n379) );
  AND U10338 ( .A(n10430), .B(n10431), .Z(n10429) );
  XNOR U10339 ( .A(p_input[671]), .B(n10428), .Z(n10431) );
  XOR U10340 ( .A(n10428), .B(p_input[655]), .Z(n10430) );
  XOR U10341 ( .A(n10432), .B(n10433), .Z(n10428) );
  AND U10342 ( .A(n10434), .B(n10435), .Z(n10433) );
  XNOR U10343 ( .A(p_input[670]), .B(n10432), .Z(n10435) );
  XNOR U10344 ( .A(n10432), .B(n10242), .Z(n10434) );
  IV U10345 ( .A(p_input[654]), .Z(n10242) );
  XOR U10346 ( .A(n10436), .B(n10437), .Z(n10432) );
  AND U10347 ( .A(n10438), .B(n10439), .Z(n10437) );
  XNOR U10348 ( .A(p_input[669]), .B(n10436), .Z(n10439) );
  XNOR U10349 ( .A(n10436), .B(n10251), .Z(n10438) );
  IV U10350 ( .A(p_input[653]), .Z(n10251) );
  XOR U10351 ( .A(n10440), .B(n10441), .Z(n10436) );
  AND U10352 ( .A(n10442), .B(n10443), .Z(n10441) );
  XNOR U10353 ( .A(p_input[668]), .B(n10440), .Z(n10443) );
  XNOR U10354 ( .A(n10440), .B(n10260), .Z(n10442) );
  IV U10355 ( .A(p_input[652]), .Z(n10260) );
  XOR U10356 ( .A(n10444), .B(n10445), .Z(n10440) );
  AND U10357 ( .A(n10446), .B(n10447), .Z(n10445) );
  XNOR U10358 ( .A(p_input[667]), .B(n10444), .Z(n10447) );
  XNOR U10359 ( .A(n10444), .B(n10269), .Z(n10446) );
  IV U10360 ( .A(p_input[651]), .Z(n10269) );
  XOR U10361 ( .A(n10448), .B(n10449), .Z(n10444) );
  AND U10362 ( .A(n10450), .B(n10451), .Z(n10449) );
  XNOR U10363 ( .A(p_input[666]), .B(n10448), .Z(n10451) );
  XNOR U10364 ( .A(n10448), .B(n10278), .Z(n10450) );
  IV U10365 ( .A(p_input[650]), .Z(n10278) );
  XOR U10366 ( .A(n10452), .B(n10453), .Z(n10448) );
  AND U10367 ( .A(n10454), .B(n10455), .Z(n10453) );
  XNOR U10368 ( .A(p_input[665]), .B(n10452), .Z(n10455) );
  XNOR U10369 ( .A(n10452), .B(n10287), .Z(n10454) );
  IV U10370 ( .A(p_input[649]), .Z(n10287) );
  XOR U10371 ( .A(n10456), .B(n10457), .Z(n10452) );
  AND U10372 ( .A(n10458), .B(n10459), .Z(n10457) );
  XNOR U10373 ( .A(p_input[664]), .B(n10456), .Z(n10459) );
  XNOR U10374 ( .A(n10456), .B(n10296), .Z(n10458) );
  IV U10375 ( .A(p_input[648]), .Z(n10296) );
  XOR U10376 ( .A(n10460), .B(n10461), .Z(n10456) );
  AND U10377 ( .A(n10462), .B(n10463), .Z(n10461) );
  XNOR U10378 ( .A(p_input[663]), .B(n10460), .Z(n10463) );
  XNOR U10379 ( .A(n10460), .B(n10305), .Z(n10462) );
  IV U10380 ( .A(p_input[647]), .Z(n10305) );
  XOR U10381 ( .A(n10464), .B(n10465), .Z(n10460) );
  AND U10382 ( .A(n10466), .B(n10467), .Z(n10465) );
  XNOR U10383 ( .A(p_input[662]), .B(n10464), .Z(n10467) );
  XNOR U10384 ( .A(n10464), .B(n10314), .Z(n10466) );
  IV U10385 ( .A(p_input[646]), .Z(n10314) );
  XOR U10386 ( .A(n10468), .B(n10469), .Z(n10464) );
  AND U10387 ( .A(n10470), .B(n10471), .Z(n10469) );
  XNOR U10388 ( .A(p_input[661]), .B(n10468), .Z(n10471) );
  XNOR U10389 ( .A(n10468), .B(n10323), .Z(n10470) );
  IV U10390 ( .A(p_input[645]), .Z(n10323) );
  XOR U10391 ( .A(n10472), .B(n10473), .Z(n10468) );
  AND U10392 ( .A(n10474), .B(n10475), .Z(n10473) );
  XNOR U10393 ( .A(p_input[660]), .B(n10472), .Z(n10475) );
  XNOR U10394 ( .A(n10472), .B(n10332), .Z(n10474) );
  IV U10395 ( .A(p_input[644]), .Z(n10332) );
  XOR U10396 ( .A(n10476), .B(n10477), .Z(n10472) );
  AND U10397 ( .A(n10478), .B(n10479), .Z(n10477) );
  XNOR U10398 ( .A(p_input[659]), .B(n10476), .Z(n10479) );
  XNOR U10399 ( .A(n10476), .B(n10341), .Z(n10478) );
  IV U10400 ( .A(p_input[643]), .Z(n10341) );
  XOR U10401 ( .A(n10480), .B(n10481), .Z(n10476) );
  AND U10402 ( .A(n10482), .B(n10483), .Z(n10481) );
  XNOR U10403 ( .A(p_input[658]), .B(n10480), .Z(n10483) );
  XNOR U10404 ( .A(n10480), .B(n10350), .Z(n10482) );
  IV U10405 ( .A(p_input[642]), .Z(n10350) );
  XNOR U10406 ( .A(n10484), .B(n10485), .Z(n10480) );
  AND U10407 ( .A(n10486), .B(n10487), .Z(n10485) );
  XOR U10408 ( .A(p_input[657]), .B(n10484), .Z(n10487) );
  XNOR U10409 ( .A(p_input[641]), .B(n10484), .Z(n10486) );
  AND U10410 ( .A(p_input[656]), .B(n10488), .Z(n10484) );
  IV U10411 ( .A(p_input[640]), .Z(n10488) );
  XOR U10412 ( .A(n10489), .B(n10490), .Z(n9604) );
  AND U10413 ( .A(n439), .B(n10491), .Z(n10490) );
  XNOR U10414 ( .A(n10492), .B(n10489), .Z(n10491) );
  XOR U10415 ( .A(n10493), .B(n10494), .Z(n439) );
  AND U10416 ( .A(n10495), .B(n10496), .Z(n10494) );
  XNOR U10417 ( .A(n9616), .B(n10493), .Z(n10496) );
  AND U10418 ( .A(n10497), .B(n10498), .Z(n9616) );
  XOR U10419 ( .A(n10493), .B(n9615), .Z(n10495) );
  AND U10420 ( .A(n10499), .B(n10500), .Z(n9615) );
  XOR U10421 ( .A(n10501), .B(n10502), .Z(n10493) );
  AND U10422 ( .A(n10503), .B(n10504), .Z(n10502) );
  XOR U10423 ( .A(n10501), .B(n9628), .Z(n10504) );
  XOR U10424 ( .A(n10505), .B(n10506), .Z(n9628) );
  AND U10425 ( .A(n302), .B(n10507), .Z(n10506) );
  XOR U10426 ( .A(n10508), .B(n10505), .Z(n10507) );
  XNOR U10427 ( .A(n9625), .B(n10501), .Z(n10503) );
  XOR U10428 ( .A(n10509), .B(n10510), .Z(n9625) );
  AND U10429 ( .A(n299), .B(n10511), .Z(n10510) );
  XOR U10430 ( .A(n10512), .B(n10509), .Z(n10511) );
  XOR U10431 ( .A(n10513), .B(n10514), .Z(n10501) );
  AND U10432 ( .A(n10515), .B(n10516), .Z(n10514) );
  XOR U10433 ( .A(n10513), .B(n9640), .Z(n10516) );
  XOR U10434 ( .A(n10517), .B(n10518), .Z(n9640) );
  AND U10435 ( .A(n302), .B(n10519), .Z(n10518) );
  XOR U10436 ( .A(n10520), .B(n10517), .Z(n10519) );
  XNOR U10437 ( .A(n9637), .B(n10513), .Z(n10515) );
  XOR U10438 ( .A(n10521), .B(n10522), .Z(n9637) );
  AND U10439 ( .A(n299), .B(n10523), .Z(n10522) );
  XOR U10440 ( .A(n10524), .B(n10521), .Z(n10523) );
  XOR U10441 ( .A(n10525), .B(n10526), .Z(n10513) );
  AND U10442 ( .A(n10527), .B(n10528), .Z(n10526) );
  XOR U10443 ( .A(n10525), .B(n9652), .Z(n10528) );
  XOR U10444 ( .A(n10529), .B(n10530), .Z(n9652) );
  AND U10445 ( .A(n302), .B(n10531), .Z(n10530) );
  XOR U10446 ( .A(n10532), .B(n10529), .Z(n10531) );
  XNOR U10447 ( .A(n9649), .B(n10525), .Z(n10527) );
  XOR U10448 ( .A(n10533), .B(n10534), .Z(n9649) );
  AND U10449 ( .A(n299), .B(n10535), .Z(n10534) );
  XOR U10450 ( .A(n10536), .B(n10533), .Z(n10535) );
  XOR U10451 ( .A(n10537), .B(n10538), .Z(n10525) );
  AND U10452 ( .A(n10539), .B(n10540), .Z(n10538) );
  XOR U10453 ( .A(n10537), .B(n9664), .Z(n10540) );
  XOR U10454 ( .A(n10541), .B(n10542), .Z(n9664) );
  AND U10455 ( .A(n302), .B(n10543), .Z(n10542) );
  XOR U10456 ( .A(n10544), .B(n10541), .Z(n10543) );
  XNOR U10457 ( .A(n9661), .B(n10537), .Z(n10539) );
  XOR U10458 ( .A(n10545), .B(n10546), .Z(n9661) );
  AND U10459 ( .A(n299), .B(n10547), .Z(n10546) );
  XOR U10460 ( .A(n10548), .B(n10545), .Z(n10547) );
  XOR U10461 ( .A(n10549), .B(n10550), .Z(n10537) );
  AND U10462 ( .A(n10551), .B(n10552), .Z(n10550) );
  XOR U10463 ( .A(n10549), .B(n9676), .Z(n10552) );
  XOR U10464 ( .A(n10553), .B(n10554), .Z(n9676) );
  AND U10465 ( .A(n302), .B(n10555), .Z(n10554) );
  XOR U10466 ( .A(n10556), .B(n10553), .Z(n10555) );
  XNOR U10467 ( .A(n9673), .B(n10549), .Z(n10551) );
  XOR U10468 ( .A(n10557), .B(n10558), .Z(n9673) );
  AND U10469 ( .A(n299), .B(n10559), .Z(n10558) );
  XOR U10470 ( .A(n10560), .B(n10557), .Z(n10559) );
  XOR U10471 ( .A(n10561), .B(n10562), .Z(n10549) );
  AND U10472 ( .A(n10563), .B(n10564), .Z(n10562) );
  XOR U10473 ( .A(n10561), .B(n9688), .Z(n10564) );
  XOR U10474 ( .A(n10565), .B(n10566), .Z(n9688) );
  AND U10475 ( .A(n302), .B(n10567), .Z(n10566) );
  XOR U10476 ( .A(n10568), .B(n10565), .Z(n10567) );
  XNOR U10477 ( .A(n9685), .B(n10561), .Z(n10563) );
  XOR U10478 ( .A(n10569), .B(n10570), .Z(n9685) );
  AND U10479 ( .A(n299), .B(n10571), .Z(n10570) );
  XOR U10480 ( .A(n10572), .B(n10569), .Z(n10571) );
  XOR U10481 ( .A(n10573), .B(n10574), .Z(n10561) );
  AND U10482 ( .A(n10575), .B(n10576), .Z(n10574) );
  XOR U10483 ( .A(n10573), .B(n9700), .Z(n10576) );
  XOR U10484 ( .A(n10577), .B(n10578), .Z(n9700) );
  AND U10485 ( .A(n302), .B(n10579), .Z(n10578) );
  XOR U10486 ( .A(n10580), .B(n10577), .Z(n10579) );
  XNOR U10487 ( .A(n9697), .B(n10573), .Z(n10575) );
  XOR U10488 ( .A(n10581), .B(n10582), .Z(n9697) );
  AND U10489 ( .A(n299), .B(n10583), .Z(n10582) );
  XOR U10490 ( .A(n10584), .B(n10581), .Z(n10583) );
  XOR U10491 ( .A(n10585), .B(n10586), .Z(n10573) );
  AND U10492 ( .A(n10587), .B(n10588), .Z(n10586) );
  XOR U10493 ( .A(n10585), .B(n9712), .Z(n10588) );
  XOR U10494 ( .A(n10589), .B(n10590), .Z(n9712) );
  AND U10495 ( .A(n302), .B(n10591), .Z(n10590) );
  XOR U10496 ( .A(n10592), .B(n10589), .Z(n10591) );
  XNOR U10497 ( .A(n9709), .B(n10585), .Z(n10587) );
  XOR U10498 ( .A(n10593), .B(n10594), .Z(n9709) );
  AND U10499 ( .A(n299), .B(n10595), .Z(n10594) );
  XOR U10500 ( .A(n10596), .B(n10593), .Z(n10595) );
  XOR U10501 ( .A(n10597), .B(n10598), .Z(n10585) );
  AND U10502 ( .A(n10599), .B(n10600), .Z(n10598) );
  XOR U10503 ( .A(n10597), .B(n9724), .Z(n10600) );
  XOR U10504 ( .A(n10601), .B(n10602), .Z(n9724) );
  AND U10505 ( .A(n302), .B(n10603), .Z(n10602) );
  XOR U10506 ( .A(n10604), .B(n10601), .Z(n10603) );
  XNOR U10507 ( .A(n9721), .B(n10597), .Z(n10599) );
  XOR U10508 ( .A(n10605), .B(n10606), .Z(n9721) );
  AND U10509 ( .A(n299), .B(n10607), .Z(n10606) );
  XOR U10510 ( .A(n10608), .B(n10605), .Z(n10607) );
  XOR U10511 ( .A(n10609), .B(n10610), .Z(n10597) );
  AND U10512 ( .A(n10611), .B(n10612), .Z(n10610) );
  XOR U10513 ( .A(n10609), .B(n9736), .Z(n10612) );
  XOR U10514 ( .A(n10613), .B(n10614), .Z(n9736) );
  AND U10515 ( .A(n302), .B(n10615), .Z(n10614) );
  XOR U10516 ( .A(n10616), .B(n10613), .Z(n10615) );
  XNOR U10517 ( .A(n9733), .B(n10609), .Z(n10611) );
  XOR U10518 ( .A(n10617), .B(n10618), .Z(n9733) );
  AND U10519 ( .A(n299), .B(n10619), .Z(n10618) );
  XOR U10520 ( .A(n10620), .B(n10617), .Z(n10619) );
  XOR U10521 ( .A(n10621), .B(n10622), .Z(n10609) );
  AND U10522 ( .A(n10623), .B(n10624), .Z(n10622) );
  XOR U10523 ( .A(n10621), .B(n9748), .Z(n10624) );
  XOR U10524 ( .A(n10625), .B(n10626), .Z(n9748) );
  AND U10525 ( .A(n302), .B(n10627), .Z(n10626) );
  XOR U10526 ( .A(n10628), .B(n10625), .Z(n10627) );
  XNOR U10527 ( .A(n9745), .B(n10621), .Z(n10623) );
  XOR U10528 ( .A(n10629), .B(n10630), .Z(n9745) );
  AND U10529 ( .A(n299), .B(n10631), .Z(n10630) );
  XOR U10530 ( .A(n10632), .B(n10629), .Z(n10631) );
  XOR U10531 ( .A(n10633), .B(n10634), .Z(n10621) );
  AND U10532 ( .A(n10635), .B(n10636), .Z(n10634) );
  XOR U10533 ( .A(n10633), .B(n9760), .Z(n10636) );
  XOR U10534 ( .A(n10637), .B(n10638), .Z(n9760) );
  AND U10535 ( .A(n302), .B(n10639), .Z(n10638) );
  XOR U10536 ( .A(n10640), .B(n10637), .Z(n10639) );
  XNOR U10537 ( .A(n9757), .B(n10633), .Z(n10635) );
  XOR U10538 ( .A(n10641), .B(n10642), .Z(n9757) );
  AND U10539 ( .A(n299), .B(n10643), .Z(n10642) );
  XOR U10540 ( .A(n10644), .B(n10641), .Z(n10643) );
  XOR U10541 ( .A(n10645), .B(n10646), .Z(n10633) );
  AND U10542 ( .A(n10647), .B(n10648), .Z(n10646) );
  XOR U10543 ( .A(n9772), .B(n10645), .Z(n10648) );
  XOR U10544 ( .A(n10649), .B(n10650), .Z(n9772) );
  AND U10545 ( .A(n302), .B(n10651), .Z(n10650) );
  XOR U10546 ( .A(n10649), .B(n10652), .Z(n10651) );
  XNOR U10547 ( .A(n10645), .B(n9769), .Z(n10647) );
  XOR U10548 ( .A(n10653), .B(n10654), .Z(n9769) );
  AND U10549 ( .A(n299), .B(n10655), .Z(n10654) );
  XOR U10550 ( .A(n10653), .B(n10656), .Z(n10655) );
  XOR U10551 ( .A(n10657), .B(n10658), .Z(n10645) );
  AND U10552 ( .A(n10659), .B(n10660), .Z(n10658) );
  XNOR U10553 ( .A(n10661), .B(n9785), .Z(n10660) );
  XOR U10554 ( .A(n10662), .B(n10663), .Z(n9785) );
  AND U10555 ( .A(n302), .B(n10664), .Z(n10663) );
  XOR U10556 ( .A(n10665), .B(n10662), .Z(n10664) );
  XNOR U10557 ( .A(n9782), .B(n10657), .Z(n10659) );
  XOR U10558 ( .A(n10666), .B(n10667), .Z(n9782) );
  AND U10559 ( .A(n299), .B(n10668), .Z(n10667) );
  XOR U10560 ( .A(n10669), .B(n10666), .Z(n10668) );
  IV U10561 ( .A(n10661), .Z(n10657) );
  AND U10562 ( .A(n10489), .B(n10492), .Z(n10661) );
  XNOR U10563 ( .A(n10670), .B(n10671), .Z(n10492) );
  AND U10564 ( .A(n302), .B(n10672), .Z(n10671) );
  XNOR U10565 ( .A(n10673), .B(n10670), .Z(n10672) );
  XOR U10566 ( .A(n10674), .B(n10675), .Z(n302) );
  AND U10567 ( .A(n10676), .B(n10677), .Z(n10675) );
  XNOR U10568 ( .A(n10497), .B(n10674), .Z(n10677) );
  AND U10569 ( .A(p_input[639]), .B(p_input[623]), .Z(n10497) );
  XOR U10570 ( .A(n10674), .B(n10498), .Z(n10676) );
  AND U10571 ( .A(p_input[607]), .B(p_input[591]), .Z(n10498) );
  XOR U10572 ( .A(n10678), .B(n10679), .Z(n10674) );
  AND U10573 ( .A(n10680), .B(n10681), .Z(n10679) );
  XOR U10574 ( .A(n10678), .B(n10508), .Z(n10681) );
  XNOR U10575 ( .A(p_input[622]), .B(n10682), .Z(n10508) );
  AND U10576 ( .A(n390), .B(n10683), .Z(n10682) );
  XOR U10577 ( .A(p_input[638]), .B(p_input[622]), .Z(n10683) );
  XNOR U10578 ( .A(n10505), .B(n10678), .Z(n10680) );
  XOR U10579 ( .A(n10684), .B(n10685), .Z(n10505) );
  AND U10580 ( .A(n388), .B(n10686), .Z(n10685) );
  XOR U10581 ( .A(p_input[606]), .B(p_input[590]), .Z(n10686) );
  XOR U10582 ( .A(n10687), .B(n10688), .Z(n10678) );
  AND U10583 ( .A(n10689), .B(n10690), .Z(n10688) );
  XOR U10584 ( .A(n10687), .B(n10520), .Z(n10690) );
  XNOR U10585 ( .A(p_input[621]), .B(n10691), .Z(n10520) );
  AND U10586 ( .A(n390), .B(n10692), .Z(n10691) );
  XOR U10587 ( .A(p_input[637]), .B(p_input[621]), .Z(n10692) );
  XNOR U10588 ( .A(n10517), .B(n10687), .Z(n10689) );
  XOR U10589 ( .A(n10693), .B(n10694), .Z(n10517) );
  AND U10590 ( .A(n388), .B(n10695), .Z(n10694) );
  XOR U10591 ( .A(p_input[605]), .B(p_input[589]), .Z(n10695) );
  XOR U10592 ( .A(n10696), .B(n10697), .Z(n10687) );
  AND U10593 ( .A(n10698), .B(n10699), .Z(n10697) );
  XOR U10594 ( .A(n10696), .B(n10532), .Z(n10699) );
  XNOR U10595 ( .A(p_input[620]), .B(n10700), .Z(n10532) );
  AND U10596 ( .A(n390), .B(n10701), .Z(n10700) );
  XOR U10597 ( .A(p_input[636]), .B(p_input[620]), .Z(n10701) );
  XNOR U10598 ( .A(n10529), .B(n10696), .Z(n10698) );
  XOR U10599 ( .A(n10702), .B(n10703), .Z(n10529) );
  AND U10600 ( .A(n388), .B(n10704), .Z(n10703) );
  XOR U10601 ( .A(p_input[604]), .B(p_input[588]), .Z(n10704) );
  XOR U10602 ( .A(n10705), .B(n10706), .Z(n10696) );
  AND U10603 ( .A(n10707), .B(n10708), .Z(n10706) );
  XOR U10604 ( .A(n10705), .B(n10544), .Z(n10708) );
  XNOR U10605 ( .A(p_input[619]), .B(n10709), .Z(n10544) );
  AND U10606 ( .A(n390), .B(n10710), .Z(n10709) );
  XOR U10607 ( .A(p_input[635]), .B(p_input[619]), .Z(n10710) );
  XNOR U10608 ( .A(n10541), .B(n10705), .Z(n10707) );
  XOR U10609 ( .A(n10711), .B(n10712), .Z(n10541) );
  AND U10610 ( .A(n388), .B(n10713), .Z(n10712) );
  XOR U10611 ( .A(p_input[603]), .B(p_input[587]), .Z(n10713) );
  XOR U10612 ( .A(n10714), .B(n10715), .Z(n10705) );
  AND U10613 ( .A(n10716), .B(n10717), .Z(n10715) );
  XOR U10614 ( .A(n10714), .B(n10556), .Z(n10717) );
  XNOR U10615 ( .A(p_input[618]), .B(n10718), .Z(n10556) );
  AND U10616 ( .A(n390), .B(n10719), .Z(n10718) );
  XOR U10617 ( .A(p_input[634]), .B(p_input[618]), .Z(n10719) );
  XNOR U10618 ( .A(n10553), .B(n10714), .Z(n10716) );
  XOR U10619 ( .A(n10720), .B(n10721), .Z(n10553) );
  AND U10620 ( .A(n388), .B(n10722), .Z(n10721) );
  XOR U10621 ( .A(p_input[602]), .B(p_input[586]), .Z(n10722) );
  XOR U10622 ( .A(n10723), .B(n10724), .Z(n10714) );
  AND U10623 ( .A(n10725), .B(n10726), .Z(n10724) );
  XOR U10624 ( .A(n10723), .B(n10568), .Z(n10726) );
  XNOR U10625 ( .A(p_input[617]), .B(n10727), .Z(n10568) );
  AND U10626 ( .A(n390), .B(n10728), .Z(n10727) );
  XOR U10627 ( .A(p_input[633]), .B(p_input[617]), .Z(n10728) );
  XNOR U10628 ( .A(n10565), .B(n10723), .Z(n10725) );
  XOR U10629 ( .A(n10729), .B(n10730), .Z(n10565) );
  AND U10630 ( .A(n388), .B(n10731), .Z(n10730) );
  XOR U10631 ( .A(p_input[601]), .B(p_input[585]), .Z(n10731) );
  XOR U10632 ( .A(n10732), .B(n10733), .Z(n10723) );
  AND U10633 ( .A(n10734), .B(n10735), .Z(n10733) );
  XOR U10634 ( .A(n10732), .B(n10580), .Z(n10735) );
  XNOR U10635 ( .A(p_input[616]), .B(n10736), .Z(n10580) );
  AND U10636 ( .A(n390), .B(n10737), .Z(n10736) );
  XOR U10637 ( .A(p_input[632]), .B(p_input[616]), .Z(n10737) );
  XNOR U10638 ( .A(n10577), .B(n10732), .Z(n10734) );
  XOR U10639 ( .A(n10738), .B(n10739), .Z(n10577) );
  AND U10640 ( .A(n388), .B(n10740), .Z(n10739) );
  XOR U10641 ( .A(p_input[600]), .B(p_input[584]), .Z(n10740) );
  XOR U10642 ( .A(n10741), .B(n10742), .Z(n10732) );
  AND U10643 ( .A(n10743), .B(n10744), .Z(n10742) );
  XOR U10644 ( .A(n10741), .B(n10592), .Z(n10744) );
  XNOR U10645 ( .A(p_input[615]), .B(n10745), .Z(n10592) );
  AND U10646 ( .A(n390), .B(n10746), .Z(n10745) );
  XOR U10647 ( .A(p_input[631]), .B(p_input[615]), .Z(n10746) );
  XNOR U10648 ( .A(n10589), .B(n10741), .Z(n10743) );
  XOR U10649 ( .A(n10747), .B(n10748), .Z(n10589) );
  AND U10650 ( .A(n388), .B(n10749), .Z(n10748) );
  XOR U10651 ( .A(p_input[599]), .B(p_input[583]), .Z(n10749) );
  XOR U10652 ( .A(n10750), .B(n10751), .Z(n10741) );
  AND U10653 ( .A(n10752), .B(n10753), .Z(n10751) );
  XOR U10654 ( .A(n10750), .B(n10604), .Z(n10753) );
  XNOR U10655 ( .A(p_input[614]), .B(n10754), .Z(n10604) );
  AND U10656 ( .A(n390), .B(n10755), .Z(n10754) );
  XOR U10657 ( .A(p_input[630]), .B(p_input[614]), .Z(n10755) );
  XNOR U10658 ( .A(n10601), .B(n10750), .Z(n10752) );
  XOR U10659 ( .A(n10756), .B(n10757), .Z(n10601) );
  AND U10660 ( .A(n388), .B(n10758), .Z(n10757) );
  XOR U10661 ( .A(p_input[598]), .B(p_input[582]), .Z(n10758) );
  XOR U10662 ( .A(n10759), .B(n10760), .Z(n10750) );
  AND U10663 ( .A(n10761), .B(n10762), .Z(n10760) );
  XOR U10664 ( .A(n10759), .B(n10616), .Z(n10762) );
  XNOR U10665 ( .A(p_input[613]), .B(n10763), .Z(n10616) );
  AND U10666 ( .A(n390), .B(n10764), .Z(n10763) );
  XOR U10667 ( .A(p_input[629]), .B(p_input[613]), .Z(n10764) );
  XNOR U10668 ( .A(n10613), .B(n10759), .Z(n10761) );
  XOR U10669 ( .A(n10765), .B(n10766), .Z(n10613) );
  AND U10670 ( .A(n388), .B(n10767), .Z(n10766) );
  XOR U10671 ( .A(p_input[597]), .B(p_input[581]), .Z(n10767) );
  XOR U10672 ( .A(n10768), .B(n10769), .Z(n10759) );
  AND U10673 ( .A(n10770), .B(n10771), .Z(n10769) );
  XOR U10674 ( .A(n10768), .B(n10628), .Z(n10771) );
  XNOR U10675 ( .A(p_input[612]), .B(n10772), .Z(n10628) );
  AND U10676 ( .A(n390), .B(n10773), .Z(n10772) );
  XOR U10677 ( .A(p_input[628]), .B(p_input[612]), .Z(n10773) );
  XNOR U10678 ( .A(n10625), .B(n10768), .Z(n10770) );
  XOR U10679 ( .A(n10774), .B(n10775), .Z(n10625) );
  AND U10680 ( .A(n388), .B(n10776), .Z(n10775) );
  XOR U10681 ( .A(p_input[596]), .B(p_input[580]), .Z(n10776) );
  XOR U10682 ( .A(n10777), .B(n10778), .Z(n10768) );
  AND U10683 ( .A(n10779), .B(n10780), .Z(n10778) );
  XOR U10684 ( .A(n10777), .B(n10640), .Z(n10780) );
  XNOR U10685 ( .A(p_input[611]), .B(n10781), .Z(n10640) );
  AND U10686 ( .A(n390), .B(n10782), .Z(n10781) );
  XOR U10687 ( .A(p_input[627]), .B(p_input[611]), .Z(n10782) );
  XNOR U10688 ( .A(n10637), .B(n10777), .Z(n10779) );
  XOR U10689 ( .A(n10783), .B(n10784), .Z(n10637) );
  AND U10690 ( .A(n388), .B(n10785), .Z(n10784) );
  XOR U10691 ( .A(p_input[595]), .B(p_input[579]), .Z(n10785) );
  XOR U10692 ( .A(n10786), .B(n10787), .Z(n10777) );
  AND U10693 ( .A(n10788), .B(n10789), .Z(n10787) );
  XOR U10694 ( .A(n10652), .B(n10786), .Z(n10789) );
  XNOR U10695 ( .A(p_input[610]), .B(n10790), .Z(n10652) );
  AND U10696 ( .A(n390), .B(n10791), .Z(n10790) );
  XOR U10697 ( .A(p_input[626]), .B(p_input[610]), .Z(n10791) );
  XNOR U10698 ( .A(n10786), .B(n10649), .Z(n10788) );
  XOR U10699 ( .A(n10792), .B(n10793), .Z(n10649) );
  AND U10700 ( .A(n388), .B(n10794), .Z(n10793) );
  XOR U10701 ( .A(p_input[594]), .B(p_input[578]), .Z(n10794) );
  XOR U10702 ( .A(n10795), .B(n10796), .Z(n10786) );
  AND U10703 ( .A(n10797), .B(n10798), .Z(n10796) );
  XNOR U10704 ( .A(n10799), .B(n10665), .Z(n10798) );
  XNOR U10705 ( .A(p_input[609]), .B(n10800), .Z(n10665) );
  AND U10706 ( .A(n390), .B(n10801), .Z(n10800) );
  XNOR U10707 ( .A(p_input[625]), .B(n10802), .Z(n10801) );
  IV U10708 ( .A(p_input[609]), .Z(n10802) );
  XNOR U10709 ( .A(n10662), .B(n10795), .Z(n10797) );
  XNOR U10710 ( .A(p_input[577]), .B(n10803), .Z(n10662) );
  AND U10711 ( .A(n388), .B(n10804), .Z(n10803) );
  XOR U10712 ( .A(p_input[593]), .B(p_input[577]), .Z(n10804) );
  IV U10713 ( .A(n10799), .Z(n10795) );
  AND U10714 ( .A(n10670), .B(n10673), .Z(n10799) );
  XOR U10715 ( .A(p_input[608]), .B(n10805), .Z(n10673) );
  AND U10716 ( .A(n390), .B(n10806), .Z(n10805) );
  XOR U10717 ( .A(p_input[624]), .B(p_input[608]), .Z(n10806) );
  XOR U10718 ( .A(n10807), .B(n10808), .Z(n390) );
  AND U10719 ( .A(n10809), .B(n10810), .Z(n10808) );
  XNOR U10720 ( .A(p_input[639]), .B(n10807), .Z(n10810) );
  XOR U10721 ( .A(n10807), .B(p_input[623]), .Z(n10809) );
  XOR U10722 ( .A(n10811), .B(n10812), .Z(n10807) );
  AND U10723 ( .A(n10813), .B(n10814), .Z(n10812) );
  XNOR U10724 ( .A(p_input[638]), .B(n10811), .Z(n10814) );
  XOR U10725 ( .A(n10811), .B(p_input[622]), .Z(n10813) );
  XOR U10726 ( .A(n10815), .B(n10816), .Z(n10811) );
  AND U10727 ( .A(n10817), .B(n10818), .Z(n10816) );
  XNOR U10728 ( .A(p_input[637]), .B(n10815), .Z(n10818) );
  XOR U10729 ( .A(n10815), .B(p_input[621]), .Z(n10817) );
  XOR U10730 ( .A(n10819), .B(n10820), .Z(n10815) );
  AND U10731 ( .A(n10821), .B(n10822), .Z(n10820) );
  XNOR U10732 ( .A(p_input[636]), .B(n10819), .Z(n10822) );
  XOR U10733 ( .A(n10819), .B(p_input[620]), .Z(n10821) );
  XOR U10734 ( .A(n10823), .B(n10824), .Z(n10819) );
  AND U10735 ( .A(n10825), .B(n10826), .Z(n10824) );
  XNOR U10736 ( .A(p_input[635]), .B(n10823), .Z(n10826) );
  XOR U10737 ( .A(n10823), .B(p_input[619]), .Z(n10825) );
  XOR U10738 ( .A(n10827), .B(n10828), .Z(n10823) );
  AND U10739 ( .A(n10829), .B(n10830), .Z(n10828) );
  XNOR U10740 ( .A(p_input[634]), .B(n10827), .Z(n10830) );
  XOR U10741 ( .A(n10827), .B(p_input[618]), .Z(n10829) );
  XOR U10742 ( .A(n10831), .B(n10832), .Z(n10827) );
  AND U10743 ( .A(n10833), .B(n10834), .Z(n10832) );
  XNOR U10744 ( .A(p_input[633]), .B(n10831), .Z(n10834) );
  XOR U10745 ( .A(n10831), .B(p_input[617]), .Z(n10833) );
  XOR U10746 ( .A(n10835), .B(n10836), .Z(n10831) );
  AND U10747 ( .A(n10837), .B(n10838), .Z(n10836) );
  XNOR U10748 ( .A(p_input[632]), .B(n10835), .Z(n10838) );
  XOR U10749 ( .A(n10835), .B(p_input[616]), .Z(n10837) );
  XOR U10750 ( .A(n10839), .B(n10840), .Z(n10835) );
  AND U10751 ( .A(n10841), .B(n10842), .Z(n10840) );
  XNOR U10752 ( .A(p_input[631]), .B(n10839), .Z(n10842) );
  XOR U10753 ( .A(n10839), .B(p_input[615]), .Z(n10841) );
  XOR U10754 ( .A(n10843), .B(n10844), .Z(n10839) );
  AND U10755 ( .A(n10845), .B(n10846), .Z(n10844) );
  XNOR U10756 ( .A(p_input[630]), .B(n10843), .Z(n10846) );
  XOR U10757 ( .A(n10843), .B(p_input[614]), .Z(n10845) );
  XOR U10758 ( .A(n10847), .B(n10848), .Z(n10843) );
  AND U10759 ( .A(n10849), .B(n10850), .Z(n10848) );
  XNOR U10760 ( .A(p_input[629]), .B(n10847), .Z(n10850) );
  XOR U10761 ( .A(n10847), .B(p_input[613]), .Z(n10849) );
  XOR U10762 ( .A(n10851), .B(n10852), .Z(n10847) );
  AND U10763 ( .A(n10853), .B(n10854), .Z(n10852) );
  XNOR U10764 ( .A(p_input[628]), .B(n10851), .Z(n10854) );
  XOR U10765 ( .A(n10851), .B(p_input[612]), .Z(n10853) );
  XOR U10766 ( .A(n10855), .B(n10856), .Z(n10851) );
  AND U10767 ( .A(n10857), .B(n10858), .Z(n10856) );
  XNOR U10768 ( .A(p_input[627]), .B(n10855), .Z(n10858) );
  XOR U10769 ( .A(n10855), .B(p_input[611]), .Z(n10857) );
  XOR U10770 ( .A(n10859), .B(n10860), .Z(n10855) );
  AND U10771 ( .A(n10861), .B(n10862), .Z(n10860) );
  XNOR U10772 ( .A(p_input[626]), .B(n10859), .Z(n10862) );
  XOR U10773 ( .A(n10859), .B(p_input[610]), .Z(n10861) );
  XNOR U10774 ( .A(n10863), .B(n10864), .Z(n10859) );
  AND U10775 ( .A(n10865), .B(n10866), .Z(n10864) );
  XOR U10776 ( .A(p_input[625]), .B(n10863), .Z(n10866) );
  XNOR U10777 ( .A(p_input[609]), .B(n10863), .Z(n10865) );
  AND U10778 ( .A(p_input[624]), .B(n10867), .Z(n10863) );
  IV U10779 ( .A(p_input[608]), .Z(n10867) );
  XNOR U10780 ( .A(p_input[576]), .B(n10868), .Z(n10670) );
  AND U10781 ( .A(n388), .B(n10869), .Z(n10868) );
  XOR U10782 ( .A(p_input[592]), .B(p_input[576]), .Z(n10869) );
  XOR U10783 ( .A(n10870), .B(n10871), .Z(n388) );
  AND U10784 ( .A(n10872), .B(n10873), .Z(n10871) );
  XNOR U10785 ( .A(p_input[607]), .B(n10870), .Z(n10873) );
  XOR U10786 ( .A(n10870), .B(p_input[591]), .Z(n10872) );
  XOR U10787 ( .A(n10874), .B(n10875), .Z(n10870) );
  AND U10788 ( .A(n10876), .B(n10877), .Z(n10875) );
  XNOR U10789 ( .A(p_input[606]), .B(n10874), .Z(n10877) );
  XNOR U10790 ( .A(n10874), .B(n10684), .Z(n10876) );
  IV U10791 ( .A(p_input[590]), .Z(n10684) );
  XOR U10792 ( .A(n10878), .B(n10879), .Z(n10874) );
  AND U10793 ( .A(n10880), .B(n10881), .Z(n10879) );
  XNOR U10794 ( .A(p_input[605]), .B(n10878), .Z(n10881) );
  XNOR U10795 ( .A(n10878), .B(n10693), .Z(n10880) );
  IV U10796 ( .A(p_input[589]), .Z(n10693) );
  XOR U10797 ( .A(n10882), .B(n10883), .Z(n10878) );
  AND U10798 ( .A(n10884), .B(n10885), .Z(n10883) );
  XNOR U10799 ( .A(p_input[604]), .B(n10882), .Z(n10885) );
  XNOR U10800 ( .A(n10882), .B(n10702), .Z(n10884) );
  IV U10801 ( .A(p_input[588]), .Z(n10702) );
  XOR U10802 ( .A(n10886), .B(n10887), .Z(n10882) );
  AND U10803 ( .A(n10888), .B(n10889), .Z(n10887) );
  XNOR U10804 ( .A(p_input[603]), .B(n10886), .Z(n10889) );
  XNOR U10805 ( .A(n10886), .B(n10711), .Z(n10888) );
  IV U10806 ( .A(p_input[587]), .Z(n10711) );
  XOR U10807 ( .A(n10890), .B(n10891), .Z(n10886) );
  AND U10808 ( .A(n10892), .B(n10893), .Z(n10891) );
  XNOR U10809 ( .A(p_input[602]), .B(n10890), .Z(n10893) );
  XNOR U10810 ( .A(n10890), .B(n10720), .Z(n10892) );
  IV U10811 ( .A(p_input[586]), .Z(n10720) );
  XOR U10812 ( .A(n10894), .B(n10895), .Z(n10890) );
  AND U10813 ( .A(n10896), .B(n10897), .Z(n10895) );
  XNOR U10814 ( .A(p_input[601]), .B(n10894), .Z(n10897) );
  XNOR U10815 ( .A(n10894), .B(n10729), .Z(n10896) );
  IV U10816 ( .A(p_input[585]), .Z(n10729) );
  XOR U10817 ( .A(n10898), .B(n10899), .Z(n10894) );
  AND U10818 ( .A(n10900), .B(n10901), .Z(n10899) );
  XNOR U10819 ( .A(p_input[600]), .B(n10898), .Z(n10901) );
  XNOR U10820 ( .A(n10898), .B(n10738), .Z(n10900) );
  IV U10821 ( .A(p_input[584]), .Z(n10738) );
  XOR U10822 ( .A(n10902), .B(n10903), .Z(n10898) );
  AND U10823 ( .A(n10904), .B(n10905), .Z(n10903) );
  XNOR U10824 ( .A(p_input[599]), .B(n10902), .Z(n10905) );
  XNOR U10825 ( .A(n10902), .B(n10747), .Z(n10904) );
  IV U10826 ( .A(p_input[583]), .Z(n10747) );
  XOR U10827 ( .A(n10906), .B(n10907), .Z(n10902) );
  AND U10828 ( .A(n10908), .B(n10909), .Z(n10907) );
  XNOR U10829 ( .A(p_input[598]), .B(n10906), .Z(n10909) );
  XNOR U10830 ( .A(n10906), .B(n10756), .Z(n10908) );
  IV U10831 ( .A(p_input[582]), .Z(n10756) );
  XOR U10832 ( .A(n10910), .B(n10911), .Z(n10906) );
  AND U10833 ( .A(n10912), .B(n10913), .Z(n10911) );
  XNOR U10834 ( .A(p_input[597]), .B(n10910), .Z(n10913) );
  XNOR U10835 ( .A(n10910), .B(n10765), .Z(n10912) );
  IV U10836 ( .A(p_input[581]), .Z(n10765) );
  XOR U10837 ( .A(n10914), .B(n10915), .Z(n10910) );
  AND U10838 ( .A(n10916), .B(n10917), .Z(n10915) );
  XNOR U10839 ( .A(p_input[596]), .B(n10914), .Z(n10917) );
  XNOR U10840 ( .A(n10914), .B(n10774), .Z(n10916) );
  IV U10841 ( .A(p_input[580]), .Z(n10774) );
  XOR U10842 ( .A(n10918), .B(n10919), .Z(n10914) );
  AND U10843 ( .A(n10920), .B(n10921), .Z(n10919) );
  XNOR U10844 ( .A(p_input[595]), .B(n10918), .Z(n10921) );
  XNOR U10845 ( .A(n10918), .B(n10783), .Z(n10920) );
  IV U10846 ( .A(p_input[579]), .Z(n10783) );
  XOR U10847 ( .A(n10922), .B(n10923), .Z(n10918) );
  AND U10848 ( .A(n10924), .B(n10925), .Z(n10923) );
  XNOR U10849 ( .A(p_input[594]), .B(n10922), .Z(n10925) );
  XNOR U10850 ( .A(n10922), .B(n10792), .Z(n10924) );
  IV U10851 ( .A(p_input[578]), .Z(n10792) );
  XNOR U10852 ( .A(n10926), .B(n10927), .Z(n10922) );
  AND U10853 ( .A(n10928), .B(n10929), .Z(n10927) );
  XOR U10854 ( .A(p_input[593]), .B(n10926), .Z(n10929) );
  XNOR U10855 ( .A(p_input[577]), .B(n10926), .Z(n10928) );
  AND U10856 ( .A(p_input[592]), .B(n10930), .Z(n10926) );
  IV U10857 ( .A(p_input[576]), .Z(n10930) );
  XOR U10858 ( .A(n10931), .B(n10932), .Z(n10489) );
  AND U10859 ( .A(n299), .B(n10933), .Z(n10932) );
  XNOR U10860 ( .A(n10934), .B(n10931), .Z(n10933) );
  XOR U10861 ( .A(n10935), .B(n10936), .Z(n299) );
  AND U10862 ( .A(n10937), .B(n10938), .Z(n10936) );
  XNOR U10863 ( .A(n10500), .B(n10935), .Z(n10938) );
  AND U10864 ( .A(p_input[575]), .B(p_input[559]), .Z(n10500) );
  XOR U10865 ( .A(n10935), .B(n10499), .Z(n10937) );
  AND U10866 ( .A(p_input[527]), .B(p_input[543]), .Z(n10499) );
  XOR U10867 ( .A(n10939), .B(n10940), .Z(n10935) );
  AND U10868 ( .A(n10941), .B(n10942), .Z(n10940) );
  XOR U10869 ( .A(n10939), .B(n10512), .Z(n10942) );
  XNOR U10870 ( .A(p_input[558]), .B(n10943), .Z(n10512) );
  AND U10871 ( .A(n394), .B(n10944), .Z(n10943) );
  XOR U10872 ( .A(p_input[574]), .B(p_input[558]), .Z(n10944) );
  XNOR U10873 ( .A(n10509), .B(n10939), .Z(n10941) );
  XOR U10874 ( .A(n10945), .B(n10946), .Z(n10509) );
  AND U10875 ( .A(n391), .B(n10947), .Z(n10946) );
  XOR U10876 ( .A(p_input[542]), .B(p_input[526]), .Z(n10947) );
  XOR U10877 ( .A(n10948), .B(n10949), .Z(n10939) );
  AND U10878 ( .A(n10950), .B(n10951), .Z(n10949) );
  XOR U10879 ( .A(n10948), .B(n10524), .Z(n10951) );
  XNOR U10880 ( .A(p_input[557]), .B(n10952), .Z(n10524) );
  AND U10881 ( .A(n394), .B(n10953), .Z(n10952) );
  XOR U10882 ( .A(p_input[573]), .B(p_input[557]), .Z(n10953) );
  XNOR U10883 ( .A(n10521), .B(n10948), .Z(n10950) );
  XOR U10884 ( .A(n10954), .B(n10955), .Z(n10521) );
  AND U10885 ( .A(n391), .B(n10956), .Z(n10955) );
  XOR U10886 ( .A(p_input[541]), .B(p_input[525]), .Z(n10956) );
  XOR U10887 ( .A(n10957), .B(n10958), .Z(n10948) );
  AND U10888 ( .A(n10959), .B(n10960), .Z(n10958) );
  XOR U10889 ( .A(n10957), .B(n10536), .Z(n10960) );
  XNOR U10890 ( .A(p_input[556]), .B(n10961), .Z(n10536) );
  AND U10891 ( .A(n394), .B(n10962), .Z(n10961) );
  XOR U10892 ( .A(p_input[572]), .B(p_input[556]), .Z(n10962) );
  XNOR U10893 ( .A(n10533), .B(n10957), .Z(n10959) );
  XOR U10894 ( .A(n10963), .B(n10964), .Z(n10533) );
  AND U10895 ( .A(n391), .B(n10965), .Z(n10964) );
  XOR U10896 ( .A(p_input[540]), .B(p_input[524]), .Z(n10965) );
  XOR U10897 ( .A(n10966), .B(n10967), .Z(n10957) );
  AND U10898 ( .A(n10968), .B(n10969), .Z(n10967) );
  XOR U10899 ( .A(n10966), .B(n10548), .Z(n10969) );
  XNOR U10900 ( .A(p_input[555]), .B(n10970), .Z(n10548) );
  AND U10901 ( .A(n394), .B(n10971), .Z(n10970) );
  XOR U10902 ( .A(p_input[571]), .B(p_input[555]), .Z(n10971) );
  XNOR U10903 ( .A(n10545), .B(n10966), .Z(n10968) );
  XOR U10904 ( .A(n10972), .B(n10973), .Z(n10545) );
  AND U10905 ( .A(n391), .B(n10974), .Z(n10973) );
  XOR U10906 ( .A(p_input[539]), .B(p_input[523]), .Z(n10974) );
  XOR U10907 ( .A(n10975), .B(n10976), .Z(n10966) );
  AND U10908 ( .A(n10977), .B(n10978), .Z(n10976) );
  XOR U10909 ( .A(n10975), .B(n10560), .Z(n10978) );
  XNOR U10910 ( .A(p_input[554]), .B(n10979), .Z(n10560) );
  AND U10911 ( .A(n394), .B(n10980), .Z(n10979) );
  XOR U10912 ( .A(p_input[570]), .B(p_input[554]), .Z(n10980) );
  XNOR U10913 ( .A(n10557), .B(n10975), .Z(n10977) );
  XOR U10914 ( .A(n10981), .B(n10982), .Z(n10557) );
  AND U10915 ( .A(n391), .B(n10983), .Z(n10982) );
  XOR U10916 ( .A(p_input[538]), .B(p_input[522]), .Z(n10983) );
  XOR U10917 ( .A(n10984), .B(n10985), .Z(n10975) );
  AND U10918 ( .A(n10986), .B(n10987), .Z(n10985) );
  XOR U10919 ( .A(n10984), .B(n10572), .Z(n10987) );
  XNOR U10920 ( .A(p_input[553]), .B(n10988), .Z(n10572) );
  AND U10921 ( .A(n394), .B(n10989), .Z(n10988) );
  XOR U10922 ( .A(p_input[569]), .B(p_input[553]), .Z(n10989) );
  XNOR U10923 ( .A(n10569), .B(n10984), .Z(n10986) );
  XOR U10924 ( .A(n10990), .B(n10991), .Z(n10569) );
  AND U10925 ( .A(n391), .B(n10992), .Z(n10991) );
  XOR U10926 ( .A(p_input[537]), .B(p_input[521]), .Z(n10992) );
  XOR U10927 ( .A(n10993), .B(n10994), .Z(n10984) );
  AND U10928 ( .A(n10995), .B(n10996), .Z(n10994) );
  XOR U10929 ( .A(n10993), .B(n10584), .Z(n10996) );
  XNOR U10930 ( .A(p_input[552]), .B(n10997), .Z(n10584) );
  AND U10931 ( .A(n394), .B(n10998), .Z(n10997) );
  XOR U10932 ( .A(p_input[568]), .B(p_input[552]), .Z(n10998) );
  XNOR U10933 ( .A(n10581), .B(n10993), .Z(n10995) );
  XOR U10934 ( .A(n10999), .B(n11000), .Z(n10581) );
  AND U10935 ( .A(n391), .B(n11001), .Z(n11000) );
  XOR U10936 ( .A(p_input[536]), .B(p_input[520]), .Z(n11001) );
  XOR U10937 ( .A(n11002), .B(n11003), .Z(n10993) );
  AND U10938 ( .A(n11004), .B(n11005), .Z(n11003) );
  XOR U10939 ( .A(n11002), .B(n10596), .Z(n11005) );
  XNOR U10940 ( .A(p_input[551]), .B(n11006), .Z(n10596) );
  AND U10941 ( .A(n394), .B(n11007), .Z(n11006) );
  XOR U10942 ( .A(p_input[567]), .B(p_input[551]), .Z(n11007) );
  XNOR U10943 ( .A(n10593), .B(n11002), .Z(n11004) );
  XOR U10944 ( .A(n11008), .B(n11009), .Z(n10593) );
  AND U10945 ( .A(n391), .B(n11010), .Z(n11009) );
  XOR U10946 ( .A(p_input[535]), .B(p_input[519]), .Z(n11010) );
  XOR U10947 ( .A(n11011), .B(n11012), .Z(n11002) );
  AND U10948 ( .A(n11013), .B(n11014), .Z(n11012) );
  XOR U10949 ( .A(n11011), .B(n10608), .Z(n11014) );
  XNOR U10950 ( .A(p_input[550]), .B(n11015), .Z(n10608) );
  AND U10951 ( .A(n394), .B(n11016), .Z(n11015) );
  XOR U10952 ( .A(p_input[566]), .B(p_input[550]), .Z(n11016) );
  XNOR U10953 ( .A(n10605), .B(n11011), .Z(n11013) );
  XOR U10954 ( .A(n11017), .B(n11018), .Z(n10605) );
  AND U10955 ( .A(n391), .B(n11019), .Z(n11018) );
  XOR U10956 ( .A(p_input[534]), .B(p_input[518]), .Z(n11019) );
  XOR U10957 ( .A(n11020), .B(n11021), .Z(n11011) );
  AND U10958 ( .A(n11022), .B(n11023), .Z(n11021) );
  XOR U10959 ( .A(n11020), .B(n10620), .Z(n11023) );
  XNOR U10960 ( .A(p_input[549]), .B(n11024), .Z(n10620) );
  AND U10961 ( .A(n394), .B(n11025), .Z(n11024) );
  XOR U10962 ( .A(p_input[565]), .B(p_input[549]), .Z(n11025) );
  XNOR U10963 ( .A(n10617), .B(n11020), .Z(n11022) );
  XOR U10964 ( .A(n11026), .B(n11027), .Z(n10617) );
  AND U10965 ( .A(n391), .B(n11028), .Z(n11027) );
  XOR U10966 ( .A(p_input[533]), .B(p_input[517]), .Z(n11028) );
  XOR U10967 ( .A(n11029), .B(n11030), .Z(n11020) );
  AND U10968 ( .A(n11031), .B(n11032), .Z(n11030) );
  XOR U10969 ( .A(n11029), .B(n10632), .Z(n11032) );
  XNOR U10970 ( .A(p_input[548]), .B(n11033), .Z(n10632) );
  AND U10971 ( .A(n394), .B(n11034), .Z(n11033) );
  XOR U10972 ( .A(p_input[564]), .B(p_input[548]), .Z(n11034) );
  XNOR U10973 ( .A(n10629), .B(n11029), .Z(n11031) );
  XOR U10974 ( .A(n11035), .B(n11036), .Z(n10629) );
  AND U10975 ( .A(n391), .B(n11037), .Z(n11036) );
  XOR U10976 ( .A(p_input[532]), .B(p_input[516]), .Z(n11037) );
  XOR U10977 ( .A(n11038), .B(n11039), .Z(n11029) );
  AND U10978 ( .A(n11040), .B(n11041), .Z(n11039) );
  XOR U10979 ( .A(n11038), .B(n10644), .Z(n11041) );
  XNOR U10980 ( .A(p_input[547]), .B(n11042), .Z(n10644) );
  AND U10981 ( .A(n394), .B(n11043), .Z(n11042) );
  XOR U10982 ( .A(p_input[563]), .B(p_input[547]), .Z(n11043) );
  XNOR U10983 ( .A(n10641), .B(n11038), .Z(n11040) );
  XOR U10984 ( .A(n11044), .B(n11045), .Z(n10641) );
  AND U10985 ( .A(n391), .B(n11046), .Z(n11045) );
  XOR U10986 ( .A(p_input[531]), .B(p_input[515]), .Z(n11046) );
  XOR U10987 ( .A(n11047), .B(n11048), .Z(n11038) );
  AND U10988 ( .A(n11049), .B(n11050), .Z(n11048) );
  XOR U10989 ( .A(n10656), .B(n11047), .Z(n11050) );
  XNOR U10990 ( .A(p_input[546]), .B(n11051), .Z(n10656) );
  AND U10991 ( .A(n394), .B(n11052), .Z(n11051) );
  XOR U10992 ( .A(p_input[562]), .B(p_input[546]), .Z(n11052) );
  XNOR U10993 ( .A(n11047), .B(n10653), .Z(n11049) );
  XOR U10994 ( .A(n11053), .B(n11054), .Z(n10653) );
  AND U10995 ( .A(n391), .B(n11055), .Z(n11054) );
  XOR U10996 ( .A(p_input[530]), .B(p_input[514]), .Z(n11055) );
  XOR U10997 ( .A(n11056), .B(n11057), .Z(n11047) );
  AND U10998 ( .A(n11058), .B(n11059), .Z(n11057) );
  XNOR U10999 ( .A(n11060), .B(n10669), .Z(n11059) );
  XNOR U11000 ( .A(p_input[545]), .B(n11061), .Z(n10669) );
  AND U11001 ( .A(n394), .B(n11062), .Z(n11061) );
  XNOR U11002 ( .A(p_input[561]), .B(n11063), .Z(n11062) );
  IV U11003 ( .A(p_input[545]), .Z(n11063) );
  XNOR U11004 ( .A(n10666), .B(n11056), .Z(n11058) );
  XNOR U11005 ( .A(p_input[513]), .B(n11064), .Z(n10666) );
  AND U11006 ( .A(n391), .B(n11065), .Z(n11064) );
  XOR U11007 ( .A(p_input[529]), .B(p_input[513]), .Z(n11065) );
  IV U11008 ( .A(n11060), .Z(n11056) );
  AND U11009 ( .A(n10931), .B(n10934), .Z(n11060) );
  XOR U11010 ( .A(p_input[544]), .B(n11066), .Z(n10934) );
  AND U11011 ( .A(n394), .B(n11067), .Z(n11066) );
  XOR U11012 ( .A(p_input[560]), .B(p_input[544]), .Z(n11067) );
  XOR U11013 ( .A(n11068), .B(n11069), .Z(n394) );
  AND U11014 ( .A(n11070), .B(n11071), .Z(n11069) );
  XNOR U11015 ( .A(p_input[575]), .B(n11068), .Z(n11071) );
  XOR U11016 ( .A(n11068), .B(p_input[559]), .Z(n11070) );
  XOR U11017 ( .A(n11072), .B(n11073), .Z(n11068) );
  AND U11018 ( .A(n11074), .B(n11075), .Z(n11073) );
  XNOR U11019 ( .A(p_input[574]), .B(n11072), .Z(n11075) );
  XOR U11020 ( .A(n11072), .B(p_input[558]), .Z(n11074) );
  XOR U11021 ( .A(n11076), .B(n11077), .Z(n11072) );
  AND U11022 ( .A(n11078), .B(n11079), .Z(n11077) );
  XNOR U11023 ( .A(p_input[573]), .B(n11076), .Z(n11079) );
  XOR U11024 ( .A(n11076), .B(p_input[557]), .Z(n11078) );
  XOR U11025 ( .A(n11080), .B(n11081), .Z(n11076) );
  AND U11026 ( .A(n11082), .B(n11083), .Z(n11081) );
  XNOR U11027 ( .A(p_input[572]), .B(n11080), .Z(n11083) );
  XOR U11028 ( .A(n11080), .B(p_input[556]), .Z(n11082) );
  XOR U11029 ( .A(n11084), .B(n11085), .Z(n11080) );
  AND U11030 ( .A(n11086), .B(n11087), .Z(n11085) );
  XNOR U11031 ( .A(p_input[571]), .B(n11084), .Z(n11087) );
  XOR U11032 ( .A(n11084), .B(p_input[555]), .Z(n11086) );
  XOR U11033 ( .A(n11088), .B(n11089), .Z(n11084) );
  AND U11034 ( .A(n11090), .B(n11091), .Z(n11089) );
  XNOR U11035 ( .A(p_input[570]), .B(n11088), .Z(n11091) );
  XOR U11036 ( .A(n11088), .B(p_input[554]), .Z(n11090) );
  XOR U11037 ( .A(n11092), .B(n11093), .Z(n11088) );
  AND U11038 ( .A(n11094), .B(n11095), .Z(n11093) );
  XNOR U11039 ( .A(p_input[569]), .B(n11092), .Z(n11095) );
  XOR U11040 ( .A(n11092), .B(p_input[553]), .Z(n11094) );
  XOR U11041 ( .A(n11096), .B(n11097), .Z(n11092) );
  AND U11042 ( .A(n11098), .B(n11099), .Z(n11097) );
  XNOR U11043 ( .A(p_input[568]), .B(n11096), .Z(n11099) );
  XOR U11044 ( .A(n11096), .B(p_input[552]), .Z(n11098) );
  XOR U11045 ( .A(n11100), .B(n11101), .Z(n11096) );
  AND U11046 ( .A(n11102), .B(n11103), .Z(n11101) );
  XNOR U11047 ( .A(p_input[567]), .B(n11100), .Z(n11103) );
  XOR U11048 ( .A(n11100), .B(p_input[551]), .Z(n11102) );
  XOR U11049 ( .A(n11104), .B(n11105), .Z(n11100) );
  AND U11050 ( .A(n11106), .B(n11107), .Z(n11105) );
  XNOR U11051 ( .A(p_input[566]), .B(n11104), .Z(n11107) );
  XOR U11052 ( .A(n11104), .B(p_input[550]), .Z(n11106) );
  XOR U11053 ( .A(n11108), .B(n11109), .Z(n11104) );
  AND U11054 ( .A(n11110), .B(n11111), .Z(n11109) );
  XNOR U11055 ( .A(p_input[565]), .B(n11108), .Z(n11111) );
  XOR U11056 ( .A(n11108), .B(p_input[549]), .Z(n11110) );
  XOR U11057 ( .A(n11112), .B(n11113), .Z(n11108) );
  AND U11058 ( .A(n11114), .B(n11115), .Z(n11113) );
  XNOR U11059 ( .A(p_input[564]), .B(n11112), .Z(n11115) );
  XOR U11060 ( .A(n11112), .B(p_input[548]), .Z(n11114) );
  XOR U11061 ( .A(n11116), .B(n11117), .Z(n11112) );
  AND U11062 ( .A(n11118), .B(n11119), .Z(n11117) );
  XNOR U11063 ( .A(p_input[563]), .B(n11116), .Z(n11119) );
  XOR U11064 ( .A(n11116), .B(p_input[547]), .Z(n11118) );
  XOR U11065 ( .A(n11120), .B(n11121), .Z(n11116) );
  AND U11066 ( .A(n11122), .B(n11123), .Z(n11121) );
  XNOR U11067 ( .A(p_input[562]), .B(n11120), .Z(n11123) );
  XOR U11068 ( .A(n11120), .B(p_input[546]), .Z(n11122) );
  XNOR U11069 ( .A(n11124), .B(n11125), .Z(n11120) );
  AND U11070 ( .A(n11126), .B(n11127), .Z(n11125) );
  XOR U11071 ( .A(p_input[561]), .B(n11124), .Z(n11127) );
  XNOR U11072 ( .A(p_input[545]), .B(n11124), .Z(n11126) );
  AND U11073 ( .A(p_input[560]), .B(n11128), .Z(n11124) );
  IV U11074 ( .A(p_input[544]), .Z(n11128) );
  XNOR U11075 ( .A(p_input[512]), .B(n11129), .Z(n10931) );
  AND U11076 ( .A(n391), .B(n11130), .Z(n11129) );
  XOR U11077 ( .A(p_input[528]), .B(p_input[512]), .Z(n11130) );
  XOR U11078 ( .A(n11131), .B(n11132), .Z(n391) );
  AND U11079 ( .A(n11133), .B(n11134), .Z(n11132) );
  XNOR U11080 ( .A(p_input[543]), .B(n11131), .Z(n11134) );
  XOR U11081 ( .A(n11131), .B(p_input[527]), .Z(n11133) );
  XOR U11082 ( .A(n11135), .B(n11136), .Z(n11131) );
  AND U11083 ( .A(n11137), .B(n11138), .Z(n11136) );
  XNOR U11084 ( .A(p_input[542]), .B(n11135), .Z(n11138) );
  XNOR U11085 ( .A(n11135), .B(n10945), .Z(n11137) );
  IV U11086 ( .A(p_input[526]), .Z(n10945) );
  XOR U11087 ( .A(n11139), .B(n11140), .Z(n11135) );
  AND U11088 ( .A(n11141), .B(n11142), .Z(n11140) );
  XNOR U11089 ( .A(p_input[541]), .B(n11139), .Z(n11142) );
  XNOR U11090 ( .A(n11139), .B(n10954), .Z(n11141) );
  IV U11091 ( .A(p_input[525]), .Z(n10954) );
  XOR U11092 ( .A(n11143), .B(n11144), .Z(n11139) );
  AND U11093 ( .A(n11145), .B(n11146), .Z(n11144) );
  XNOR U11094 ( .A(p_input[540]), .B(n11143), .Z(n11146) );
  XNOR U11095 ( .A(n11143), .B(n10963), .Z(n11145) );
  IV U11096 ( .A(p_input[524]), .Z(n10963) );
  XOR U11097 ( .A(n11147), .B(n11148), .Z(n11143) );
  AND U11098 ( .A(n11149), .B(n11150), .Z(n11148) );
  XNOR U11099 ( .A(p_input[539]), .B(n11147), .Z(n11150) );
  XNOR U11100 ( .A(n11147), .B(n10972), .Z(n11149) );
  IV U11101 ( .A(p_input[523]), .Z(n10972) );
  XOR U11102 ( .A(n11151), .B(n11152), .Z(n11147) );
  AND U11103 ( .A(n11153), .B(n11154), .Z(n11152) );
  XNOR U11104 ( .A(p_input[538]), .B(n11151), .Z(n11154) );
  XNOR U11105 ( .A(n11151), .B(n10981), .Z(n11153) );
  IV U11106 ( .A(p_input[522]), .Z(n10981) );
  XOR U11107 ( .A(n11155), .B(n11156), .Z(n11151) );
  AND U11108 ( .A(n11157), .B(n11158), .Z(n11156) );
  XNOR U11109 ( .A(p_input[537]), .B(n11155), .Z(n11158) );
  XNOR U11110 ( .A(n11155), .B(n10990), .Z(n11157) );
  IV U11111 ( .A(p_input[521]), .Z(n10990) );
  XOR U11112 ( .A(n11159), .B(n11160), .Z(n11155) );
  AND U11113 ( .A(n11161), .B(n11162), .Z(n11160) );
  XNOR U11114 ( .A(p_input[536]), .B(n11159), .Z(n11162) );
  XNOR U11115 ( .A(n11159), .B(n10999), .Z(n11161) );
  IV U11116 ( .A(p_input[520]), .Z(n10999) );
  XOR U11117 ( .A(n11163), .B(n11164), .Z(n11159) );
  AND U11118 ( .A(n11165), .B(n11166), .Z(n11164) );
  XNOR U11119 ( .A(p_input[535]), .B(n11163), .Z(n11166) );
  XNOR U11120 ( .A(n11163), .B(n11008), .Z(n11165) );
  IV U11121 ( .A(p_input[519]), .Z(n11008) );
  XOR U11122 ( .A(n11167), .B(n11168), .Z(n11163) );
  AND U11123 ( .A(n11169), .B(n11170), .Z(n11168) );
  XNOR U11124 ( .A(p_input[534]), .B(n11167), .Z(n11170) );
  XNOR U11125 ( .A(n11167), .B(n11017), .Z(n11169) );
  IV U11126 ( .A(p_input[518]), .Z(n11017) );
  XOR U11127 ( .A(n11171), .B(n11172), .Z(n11167) );
  AND U11128 ( .A(n11173), .B(n11174), .Z(n11172) );
  XNOR U11129 ( .A(p_input[533]), .B(n11171), .Z(n11174) );
  XNOR U11130 ( .A(n11171), .B(n11026), .Z(n11173) );
  IV U11131 ( .A(p_input[517]), .Z(n11026) );
  XOR U11132 ( .A(n11175), .B(n11176), .Z(n11171) );
  AND U11133 ( .A(n11177), .B(n11178), .Z(n11176) );
  XNOR U11134 ( .A(p_input[532]), .B(n11175), .Z(n11178) );
  XNOR U11135 ( .A(n11175), .B(n11035), .Z(n11177) );
  IV U11136 ( .A(p_input[516]), .Z(n11035) );
  XOR U11137 ( .A(n11179), .B(n11180), .Z(n11175) );
  AND U11138 ( .A(n11181), .B(n11182), .Z(n11180) );
  XNOR U11139 ( .A(p_input[531]), .B(n11179), .Z(n11182) );
  XNOR U11140 ( .A(n11179), .B(n11044), .Z(n11181) );
  IV U11141 ( .A(p_input[515]), .Z(n11044) );
  XOR U11142 ( .A(n11183), .B(n11184), .Z(n11179) );
  AND U11143 ( .A(n11185), .B(n11186), .Z(n11184) );
  XNOR U11144 ( .A(p_input[530]), .B(n11183), .Z(n11186) );
  XNOR U11145 ( .A(n11183), .B(n11053), .Z(n11185) );
  IV U11146 ( .A(p_input[514]), .Z(n11053) );
  XNOR U11147 ( .A(n11187), .B(n11188), .Z(n11183) );
  AND U11148 ( .A(n11189), .B(n11190), .Z(n11188) );
  XOR U11149 ( .A(p_input[529]), .B(n11187), .Z(n11190) );
  XNOR U11150 ( .A(p_input[513]), .B(n11187), .Z(n11189) );
  AND U11151 ( .A(p_input[528]), .B(n11191), .Z(n11187) );
  IV U11152 ( .A(p_input[512]), .Z(n11191) );
  XOR U11153 ( .A(n11192), .B(n11193), .Z(n7646) );
  AND U11154 ( .A(n539), .B(n11194), .Z(n11193) );
  XNOR U11155 ( .A(n11195), .B(n11192), .Z(n11194) );
  XOR U11156 ( .A(n11196), .B(n11197), .Z(n539) );
  AND U11157 ( .A(n11198), .B(n11199), .Z(n11197) );
  XOR U11158 ( .A(n11196), .B(n7661), .Z(n11199) );
  XNOR U11159 ( .A(n11200), .B(n11201), .Z(n7661) );
  AND U11160 ( .A(n11202), .B(n514), .Z(n11201) );
  AND U11161 ( .A(n11200), .B(n11203), .Z(n11202) );
  XNOR U11162 ( .A(n7658), .B(n11196), .Z(n11198) );
  XOR U11163 ( .A(n11204), .B(n11205), .Z(n7658) );
  AND U11164 ( .A(n11206), .B(n511), .Z(n11205) );
  NOR U11165 ( .A(n11204), .B(n11207), .Z(n11206) );
  XOR U11166 ( .A(n11208), .B(n11209), .Z(n11196) );
  AND U11167 ( .A(n11210), .B(n11211), .Z(n11209) );
  XOR U11168 ( .A(n11208), .B(n7673), .Z(n11211) );
  XOR U11169 ( .A(n11212), .B(n11213), .Z(n7673) );
  AND U11170 ( .A(n514), .B(n11214), .Z(n11213) );
  XOR U11171 ( .A(n11215), .B(n11212), .Z(n11214) );
  XNOR U11172 ( .A(n7670), .B(n11208), .Z(n11210) );
  XOR U11173 ( .A(n11216), .B(n11217), .Z(n7670) );
  AND U11174 ( .A(n511), .B(n11218), .Z(n11217) );
  XOR U11175 ( .A(n11219), .B(n11216), .Z(n11218) );
  XOR U11176 ( .A(n11220), .B(n11221), .Z(n11208) );
  AND U11177 ( .A(n11222), .B(n11223), .Z(n11221) );
  XOR U11178 ( .A(n11220), .B(n7685), .Z(n11223) );
  XOR U11179 ( .A(n11224), .B(n11225), .Z(n7685) );
  AND U11180 ( .A(n514), .B(n11226), .Z(n11225) );
  XOR U11181 ( .A(n11227), .B(n11224), .Z(n11226) );
  XNOR U11182 ( .A(n7682), .B(n11220), .Z(n11222) );
  XOR U11183 ( .A(n11228), .B(n11229), .Z(n7682) );
  AND U11184 ( .A(n511), .B(n11230), .Z(n11229) );
  XOR U11185 ( .A(n11231), .B(n11228), .Z(n11230) );
  XOR U11186 ( .A(n11232), .B(n11233), .Z(n11220) );
  AND U11187 ( .A(n11234), .B(n11235), .Z(n11233) );
  XOR U11188 ( .A(n11232), .B(n7697), .Z(n11235) );
  XOR U11189 ( .A(n11236), .B(n11237), .Z(n7697) );
  AND U11190 ( .A(n514), .B(n11238), .Z(n11237) );
  XOR U11191 ( .A(n11239), .B(n11236), .Z(n11238) );
  XNOR U11192 ( .A(n7694), .B(n11232), .Z(n11234) );
  XOR U11193 ( .A(n11240), .B(n11241), .Z(n7694) );
  AND U11194 ( .A(n511), .B(n11242), .Z(n11241) );
  XOR U11195 ( .A(n11243), .B(n11240), .Z(n11242) );
  XOR U11196 ( .A(n11244), .B(n11245), .Z(n11232) );
  AND U11197 ( .A(n11246), .B(n11247), .Z(n11245) );
  XOR U11198 ( .A(n11244), .B(n7709), .Z(n11247) );
  XOR U11199 ( .A(n11248), .B(n11249), .Z(n7709) );
  AND U11200 ( .A(n514), .B(n11250), .Z(n11249) );
  XOR U11201 ( .A(n11251), .B(n11248), .Z(n11250) );
  XNOR U11202 ( .A(n7706), .B(n11244), .Z(n11246) );
  XOR U11203 ( .A(n11252), .B(n11253), .Z(n7706) );
  AND U11204 ( .A(n511), .B(n11254), .Z(n11253) );
  XOR U11205 ( .A(n11255), .B(n11252), .Z(n11254) );
  XOR U11206 ( .A(n11256), .B(n11257), .Z(n11244) );
  AND U11207 ( .A(n11258), .B(n11259), .Z(n11257) );
  XOR U11208 ( .A(n11256), .B(n7721), .Z(n11259) );
  XOR U11209 ( .A(n11260), .B(n11261), .Z(n7721) );
  AND U11210 ( .A(n514), .B(n11262), .Z(n11261) );
  XOR U11211 ( .A(n11263), .B(n11260), .Z(n11262) );
  XNOR U11212 ( .A(n7718), .B(n11256), .Z(n11258) );
  XOR U11213 ( .A(n11264), .B(n11265), .Z(n7718) );
  AND U11214 ( .A(n511), .B(n11266), .Z(n11265) );
  XOR U11215 ( .A(n11267), .B(n11264), .Z(n11266) );
  XOR U11216 ( .A(n11268), .B(n11269), .Z(n11256) );
  AND U11217 ( .A(n11270), .B(n11271), .Z(n11269) );
  XOR U11218 ( .A(n11268), .B(n7733), .Z(n11271) );
  XOR U11219 ( .A(n11272), .B(n11273), .Z(n7733) );
  AND U11220 ( .A(n514), .B(n11274), .Z(n11273) );
  XOR U11221 ( .A(n11275), .B(n11272), .Z(n11274) );
  XNOR U11222 ( .A(n7730), .B(n11268), .Z(n11270) );
  XOR U11223 ( .A(n11276), .B(n11277), .Z(n7730) );
  AND U11224 ( .A(n511), .B(n11278), .Z(n11277) );
  XOR U11225 ( .A(n11279), .B(n11276), .Z(n11278) );
  XOR U11226 ( .A(n11280), .B(n11281), .Z(n11268) );
  AND U11227 ( .A(n11282), .B(n11283), .Z(n11281) );
  XOR U11228 ( .A(n11280), .B(n7745), .Z(n11283) );
  XOR U11229 ( .A(n11284), .B(n11285), .Z(n7745) );
  AND U11230 ( .A(n514), .B(n11286), .Z(n11285) );
  XOR U11231 ( .A(n11287), .B(n11284), .Z(n11286) );
  XNOR U11232 ( .A(n7742), .B(n11280), .Z(n11282) );
  XOR U11233 ( .A(n11288), .B(n11289), .Z(n7742) );
  AND U11234 ( .A(n511), .B(n11290), .Z(n11289) );
  XOR U11235 ( .A(n11291), .B(n11288), .Z(n11290) );
  XOR U11236 ( .A(n11292), .B(n11293), .Z(n11280) );
  AND U11237 ( .A(n11294), .B(n11295), .Z(n11293) );
  XOR U11238 ( .A(n11292), .B(n7757), .Z(n11295) );
  XOR U11239 ( .A(n11296), .B(n11297), .Z(n7757) );
  AND U11240 ( .A(n514), .B(n11298), .Z(n11297) );
  XOR U11241 ( .A(n11299), .B(n11296), .Z(n11298) );
  XNOR U11242 ( .A(n7754), .B(n11292), .Z(n11294) );
  XOR U11243 ( .A(n11300), .B(n11301), .Z(n7754) );
  AND U11244 ( .A(n511), .B(n11302), .Z(n11301) );
  XOR U11245 ( .A(n11303), .B(n11300), .Z(n11302) );
  XOR U11246 ( .A(n11304), .B(n11305), .Z(n11292) );
  AND U11247 ( .A(n11306), .B(n11307), .Z(n11305) );
  XOR U11248 ( .A(n11304), .B(n7769), .Z(n11307) );
  XOR U11249 ( .A(n11308), .B(n11309), .Z(n7769) );
  AND U11250 ( .A(n514), .B(n11310), .Z(n11309) );
  XOR U11251 ( .A(n11311), .B(n11308), .Z(n11310) );
  XNOR U11252 ( .A(n7766), .B(n11304), .Z(n11306) );
  XOR U11253 ( .A(n11312), .B(n11313), .Z(n7766) );
  AND U11254 ( .A(n511), .B(n11314), .Z(n11313) );
  XOR U11255 ( .A(n11315), .B(n11312), .Z(n11314) );
  XOR U11256 ( .A(n11316), .B(n11317), .Z(n11304) );
  AND U11257 ( .A(n11318), .B(n11319), .Z(n11317) );
  XOR U11258 ( .A(n11316), .B(n7781), .Z(n11319) );
  XOR U11259 ( .A(n11320), .B(n11321), .Z(n7781) );
  AND U11260 ( .A(n514), .B(n11322), .Z(n11321) );
  XOR U11261 ( .A(n11323), .B(n11320), .Z(n11322) );
  XNOR U11262 ( .A(n7778), .B(n11316), .Z(n11318) );
  XOR U11263 ( .A(n11324), .B(n11325), .Z(n7778) );
  AND U11264 ( .A(n511), .B(n11326), .Z(n11325) );
  XOR U11265 ( .A(n11327), .B(n11324), .Z(n11326) );
  XOR U11266 ( .A(n11328), .B(n11329), .Z(n11316) );
  AND U11267 ( .A(n11330), .B(n11331), .Z(n11329) );
  XOR U11268 ( .A(n11328), .B(n7793), .Z(n11331) );
  XOR U11269 ( .A(n11332), .B(n11333), .Z(n7793) );
  AND U11270 ( .A(n514), .B(n11334), .Z(n11333) );
  XOR U11271 ( .A(n11335), .B(n11332), .Z(n11334) );
  XNOR U11272 ( .A(n7790), .B(n11328), .Z(n11330) );
  XOR U11273 ( .A(n11336), .B(n11337), .Z(n7790) );
  AND U11274 ( .A(n511), .B(n11338), .Z(n11337) );
  XOR U11275 ( .A(n11339), .B(n11336), .Z(n11338) );
  XOR U11276 ( .A(n11340), .B(n11341), .Z(n11328) );
  AND U11277 ( .A(n11342), .B(n11343), .Z(n11341) );
  XOR U11278 ( .A(n11340), .B(n7805), .Z(n11343) );
  XOR U11279 ( .A(n11344), .B(n11345), .Z(n7805) );
  AND U11280 ( .A(n514), .B(n11346), .Z(n11345) );
  XOR U11281 ( .A(n11347), .B(n11344), .Z(n11346) );
  XNOR U11282 ( .A(n7802), .B(n11340), .Z(n11342) );
  XOR U11283 ( .A(n11348), .B(n11349), .Z(n7802) );
  AND U11284 ( .A(n511), .B(n11350), .Z(n11349) );
  XOR U11285 ( .A(n11351), .B(n11348), .Z(n11350) );
  XOR U11286 ( .A(n11352), .B(n11353), .Z(n11340) );
  AND U11287 ( .A(n11354), .B(n11355), .Z(n11353) );
  XOR U11288 ( .A(n7817), .B(n11352), .Z(n11355) );
  XOR U11289 ( .A(n11356), .B(n11357), .Z(n7817) );
  AND U11290 ( .A(n514), .B(n11358), .Z(n11357) );
  XOR U11291 ( .A(n11356), .B(n11359), .Z(n11358) );
  XNOR U11292 ( .A(n11352), .B(n7814), .Z(n11354) );
  XOR U11293 ( .A(n11360), .B(n11361), .Z(n7814) );
  AND U11294 ( .A(n511), .B(n11362), .Z(n11361) );
  XOR U11295 ( .A(n11360), .B(n11363), .Z(n11362) );
  XOR U11296 ( .A(n11364), .B(n11365), .Z(n11352) );
  AND U11297 ( .A(n11366), .B(n11367), .Z(n11365) );
  XNOR U11298 ( .A(n11368), .B(n7830), .Z(n11367) );
  XOR U11299 ( .A(n11369), .B(n11370), .Z(n7830) );
  AND U11300 ( .A(n514), .B(n11371), .Z(n11370) );
  XOR U11301 ( .A(n11372), .B(n11369), .Z(n11371) );
  XNOR U11302 ( .A(n7827), .B(n11364), .Z(n11366) );
  XOR U11303 ( .A(n11373), .B(n11374), .Z(n7827) );
  AND U11304 ( .A(n511), .B(n11375), .Z(n11374) );
  XOR U11305 ( .A(n11376), .B(n11373), .Z(n11375) );
  IV U11306 ( .A(n11368), .Z(n11364) );
  AND U11307 ( .A(n11192), .B(n11195), .Z(n11368) );
  XNOR U11308 ( .A(n11377), .B(n11378), .Z(n11195) );
  AND U11309 ( .A(n514), .B(n11379), .Z(n11378) );
  XNOR U11310 ( .A(n11380), .B(n11377), .Z(n11379) );
  XOR U11311 ( .A(n11381), .B(n11382), .Z(n514) );
  AND U11312 ( .A(n11383), .B(n11384), .Z(n11382) );
  XOR U11313 ( .A(n11203), .B(n11381), .Z(n11384) );
  IV U11314 ( .A(n11385), .Z(n11203) );
  AND U11315 ( .A(n11386), .B(n11387), .Z(n11385) );
  XOR U11316 ( .A(n11381), .B(n11200), .Z(n11383) );
  AND U11317 ( .A(n11388), .B(n11389), .Z(n11200) );
  XOR U11318 ( .A(n11390), .B(n11391), .Z(n11381) );
  AND U11319 ( .A(n11392), .B(n11393), .Z(n11391) );
  XOR U11320 ( .A(n11390), .B(n11215), .Z(n11393) );
  XOR U11321 ( .A(n11394), .B(n11395), .Z(n11215) );
  AND U11322 ( .A(n450), .B(n11396), .Z(n11395) );
  XOR U11323 ( .A(n11397), .B(n11394), .Z(n11396) );
  XNOR U11324 ( .A(n11212), .B(n11390), .Z(n11392) );
  XOR U11325 ( .A(n11398), .B(n11399), .Z(n11212) );
  AND U11326 ( .A(n448), .B(n11400), .Z(n11399) );
  XOR U11327 ( .A(n11401), .B(n11398), .Z(n11400) );
  XOR U11328 ( .A(n11402), .B(n11403), .Z(n11390) );
  AND U11329 ( .A(n11404), .B(n11405), .Z(n11403) );
  XOR U11330 ( .A(n11402), .B(n11227), .Z(n11405) );
  XOR U11331 ( .A(n11406), .B(n11407), .Z(n11227) );
  AND U11332 ( .A(n450), .B(n11408), .Z(n11407) );
  XOR U11333 ( .A(n11409), .B(n11406), .Z(n11408) );
  XNOR U11334 ( .A(n11224), .B(n11402), .Z(n11404) );
  XOR U11335 ( .A(n11410), .B(n11411), .Z(n11224) );
  AND U11336 ( .A(n448), .B(n11412), .Z(n11411) );
  XOR U11337 ( .A(n11413), .B(n11410), .Z(n11412) );
  XOR U11338 ( .A(n11414), .B(n11415), .Z(n11402) );
  AND U11339 ( .A(n11416), .B(n11417), .Z(n11415) );
  XOR U11340 ( .A(n11414), .B(n11239), .Z(n11417) );
  XOR U11341 ( .A(n11418), .B(n11419), .Z(n11239) );
  AND U11342 ( .A(n450), .B(n11420), .Z(n11419) );
  XOR U11343 ( .A(n11421), .B(n11418), .Z(n11420) );
  XNOR U11344 ( .A(n11236), .B(n11414), .Z(n11416) );
  XOR U11345 ( .A(n11422), .B(n11423), .Z(n11236) );
  AND U11346 ( .A(n448), .B(n11424), .Z(n11423) );
  XOR U11347 ( .A(n11425), .B(n11422), .Z(n11424) );
  XOR U11348 ( .A(n11426), .B(n11427), .Z(n11414) );
  AND U11349 ( .A(n11428), .B(n11429), .Z(n11427) );
  XOR U11350 ( .A(n11426), .B(n11251), .Z(n11429) );
  XOR U11351 ( .A(n11430), .B(n11431), .Z(n11251) );
  AND U11352 ( .A(n450), .B(n11432), .Z(n11431) );
  XOR U11353 ( .A(n11433), .B(n11430), .Z(n11432) );
  XNOR U11354 ( .A(n11248), .B(n11426), .Z(n11428) );
  XOR U11355 ( .A(n11434), .B(n11435), .Z(n11248) );
  AND U11356 ( .A(n448), .B(n11436), .Z(n11435) );
  XOR U11357 ( .A(n11437), .B(n11434), .Z(n11436) );
  XOR U11358 ( .A(n11438), .B(n11439), .Z(n11426) );
  AND U11359 ( .A(n11440), .B(n11441), .Z(n11439) );
  XOR U11360 ( .A(n11438), .B(n11263), .Z(n11441) );
  XOR U11361 ( .A(n11442), .B(n11443), .Z(n11263) );
  AND U11362 ( .A(n450), .B(n11444), .Z(n11443) );
  XOR U11363 ( .A(n11445), .B(n11442), .Z(n11444) );
  XNOR U11364 ( .A(n11260), .B(n11438), .Z(n11440) );
  XOR U11365 ( .A(n11446), .B(n11447), .Z(n11260) );
  AND U11366 ( .A(n448), .B(n11448), .Z(n11447) );
  XOR U11367 ( .A(n11449), .B(n11446), .Z(n11448) );
  XOR U11368 ( .A(n11450), .B(n11451), .Z(n11438) );
  AND U11369 ( .A(n11452), .B(n11453), .Z(n11451) );
  XOR U11370 ( .A(n11450), .B(n11275), .Z(n11453) );
  XOR U11371 ( .A(n11454), .B(n11455), .Z(n11275) );
  AND U11372 ( .A(n450), .B(n11456), .Z(n11455) );
  XOR U11373 ( .A(n11457), .B(n11454), .Z(n11456) );
  XNOR U11374 ( .A(n11272), .B(n11450), .Z(n11452) );
  XOR U11375 ( .A(n11458), .B(n11459), .Z(n11272) );
  AND U11376 ( .A(n448), .B(n11460), .Z(n11459) );
  XOR U11377 ( .A(n11461), .B(n11458), .Z(n11460) );
  XOR U11378 ( .A(n11462), .B(n11463), .Z(n11450) );
  AND U11379 ( .A(n11464), .B(n11465), .Z(n11463) );
  XOR U11380 ( .A(n11462), .B(n11287), .Z(n11465) );
  XOR U11381 ( .A(n11466), .B(n11467), .Z(n11287) );
  AND U11382 ( .A(n450), .B(n11468), .Z(n11467) );
  XOR U11383 ( .A(n11469), .B(n11466), .Z(n11468) );
  XNOR U11384 ( .A(n11284), .B(n11462), .Z(n11464) );
  XOR U11385 ( .A(n11470), .B(n11471), .Z(n11284) );
  AND U11386 ( .A(n448), .B(n11472), .Z(n11471) );
  XOR U11387 ( .A(n11473), .B(n11470), .Z(n11472) );
  XOR U11388 ( .A(n11474), .B(n11475), .Z(n11462) );
  AND U11389 ( .A(n11476), .B(n11477), .Z(n11475) );
  XOR U11390 ( .A(n11474), .B(n11299), .Z(n11477) );
  XOR U11391 ( .A(n11478), .B(n11479), .Z(n11299) );
  AND U11392 ( .A(n450), .B(n11480), .Z(n11479) );
  XOR U11393 ( .A(n11481), .B(n11478), .Z(n11480) );
  XNOR U11394 ( .A(n11296), .B(n11474), .Z(n11476) );
  XOR U11395 ( .A(n11482), .B(n11483), .Z(n11296) );
  AND U11396 ( .A(n448), .B(n11484), .Z(n11483) );
  XOR U11397 ( .A(n11485), .B(n11482), .Z(n11484) );
  XOR U11398 ( .A(n11486), .B(n11487), .Z(n11474) );
  AND U11399 ( .A(n11488), .B(n11489), .Z(n11487) );
  XOR U11400 ( .A(n11486), .B(n11311), .Z(n11489) );
  XOR U11401 ( .A(n11490), .B(n11491), .Z(n11311) );
  AND U11402 ( .A(n450), .B(n11492), .Z(n11491) );
  XOR U11403 ( .A(n11493), .B(n11490), .Z(n11492) );
  XNOR U11404 ( .A(n11308), .B(n11486), .Z(n11488) );
  XOR U11405 ( .A(n11494), .B(n11495), .Z(n11308) );
  AND U11406 ( .A(n448), .B(n11496), .Z(n11495) );
  XOR U11407 ( .A(n11497), .B(n11494), .Z(n11496) );
  XOR U11408 ( .A(n11498), .B(n11499), .Z(n11486) );
  AND U11409 ( .A(n11500), .B(n11501), .Z(n11499) );
  XOR U11410 ( .A(n11498), .B(n11323), .Z(n11501) );
  XOR U11411 ( .A(n11502), .B(n11503), .Z(n11323) );
  AND U11412 ( .A(n450), .B(n11504), .Z(n11503) );
  XOR U11413 ( .A(n11505), .B(n11502), .Z(n11504) );
  XNOR U11414 ( .A(n11320), .B(n11498), .Z(n11500) );
  XOR U11415 ( .A(n11506), .B(n11507), .Z(n11320) );
  AND U11416 ( .A(n448), .B(n11508), .Z(n11507) );
  XOR U11417 ( .A(n11509), .B(n11506), .Z(n11508) );
  XOR U11418 ( .A(n11510), .B(n11511), .Z(n11498) );
  AND U11419 ( .A(n11512), .B(n11513), .Z(n11511) );
  XOR U11420 ( .A(n11510), .B(n11335), .Z(n11513) );
  XOR U11421 ( .A(n11514), .B(n11515), .Z(n11335) );
  AND U11422 ( .A(n450), .B(n11516), .Z(n11515) );
  XOR U11423 ( .A(n11517), .B(n11514), .Z(n11516) );
  XNOR U11424 ( .A(n11332), .B(n11510), .Z(n11512) );
  XOR U11425 ( .A(n11518), .B(n11519), .Z(n11332) );
  AND U11426 ( .A(n448), .B(n11520), .Z(n11519) );
  XOR U11427 ( .A(n11521), .B(n11518), .Z(n11520) );
  XOR U11428 ( .A(n11522), .B(n11523), .Z(n11510) );
  AND U11429 ( .A(n11524), .B(n11525), .Z(n11523) );
  XOR U11430 ( .A(n11522), .B(n11347), .Z(n11525) );
  XOR U11431 ( .A(n11526), .B(n11527), .Z(n11347) );
  AND U11432 ( .A(n450), .B(n11528), .Z(n11527) );
  XOR U11433 ( .A(n11529), .B(n11526), .Z(n11528) );
  XNOR U11434 ( .A(n11344), .B(n11522), .Z(n11524) );
  XOR U11435 ( .A(n11530), .B(n11531), .Z(n11344) );
  AND U11436 ( .A(n448), .B(n11532), .Z(n11531) );
  XOR U11437 ( .A(n11533), .B(n11530), .Z(n11532) );
  XOR U11438 ( .A(n11534), .B(n11535), .Z(n11522) );
  AND U11439 ( .A(n11536), .B(n11537), .Z(n11535) );
  XOR U11440 ( .A(n11359), .B(n11534), .Z(n11537) );
  XOR U11441 ( .A(n11538), .B(n11539), .Z(n11359) );
  AND U11442 ( .A(n450), .B(n11540), .Z(n11539) );
  XOR U11443 ( .A(n11538), .B(n11541), .Z(n11540) );
  XNOR U11444 ( .A(n11534), .B(n11356), .Z(n11536) );
  XOR U11445 ( .A(n11542), .B(n11543), .Z(n11356) );
  AND U11446 ( .A(n448), .B(n11544), .Z(n11543) );
  XOR U11447 ( .A(n11542), .B(n11545), .Z(n11544) );
  XOR U11448 ( .A(n11546), .B(n11547), .Z(n11534) );
  AND U11449 ( .A(n11548), .B(n11549), .Z(n11547) );
  XNOR U11450 ( .A(n11550), .B(n11372), .Z(n11549) );
  XOR U11451 ( .A(n11551), .B(n11552), .Z(n11372) );
  AND U11452 ( .A(n450), .B(n11553), .Z(n11552) );
  XOR U11453 ( .A(n11554), .B(n11551), .Z(n11553) );
  XNOR U11454 ( .A(n11369), .B(n11546), .Z(n11548) );
  XOR U11455 ( .A(n11555), .B(n11556), .Z(n11369) );
  AND U11456 ( .A(n448), .B(n11557), .Z(n11556) );
  XOR U11457 ( .A(n11558), .B(n11555), .Z(n11557) );
  IV U11458 ( .A(n11550), .Z(n11546) );
  AND U11459 ( .A(n11377), .B(n11380), .Z(n11550) );
  XNOR U11460 ( .A(n11559), .B(n11560), .Z(n11380) );
  AND U11461 ( .A(n450), .B(n11561), .Z(n11560) );
  XNOR U11462 ( .A(n11562), .B(n11559), .Z(n11561) );
  XOR U11463 ( .A(n11563), .B(n11564), .Z(n450) );
  AND U11464 ( .A(n11565), .B(n11566), .Z(n11564) );
  XNOR U11465 ( .A(n11386), .B(n11563), .Z(n11566) );
  AND U11466 ( .A(n11567), .B(n11568), .Z(n11386) );
  XOR U11467 ( .A(n11563), .B(n11387), .Z(n11565) );
  AND U11468 ( .A(n11569), .B(n11570), .Z(n11387) );
  XOR U11469 ( .A(n11571), .B(n11572), .Z(n11563) );
  AND U11470 ( .A(n11573), .B(n11574), .Z(n11572) );
  XOR U11471 ( .A(n11571), .B(n11397), .Z(n11574) );
  XOR U11472 ( .A(n11575), .B(n11576), .Z(n11397) );
  AND U11473 ( .A(n314), .B(n11577), .Z(n11576) );
  XOR U11474 ( .A(n11578), .B(n11575), .Z(n11577) );
  XNOR U11475 ( .A(n11394), .B(n11571), .Z(n11573) );
  XOR U11476 ( .A(n11579), .B(n11580), .Z(n11394) );
  AND U11477 ( .A(n312), .B(n11581), .Z(n11580) );
  XOR U11478 ( .A(n11582), .B(n11579), .Z(n11581) );
  XOR U11479 ( .A(n11583), .B(n11584), .Z(n11571) );
  AND U11480 ( .A(n11585), .B(n11586), .Z(n11584) );
  XOR U11481 ( .A(n11583), .B(n11409), .Z(n11586) );
  XOR U11482 ( .A(n11587), .B(n11588), .Z(n11409) );
  AND U11483 ( .A(n314), .B(n11589), .Z(n11588) );
  XOR U11484 ( .A(n11590), .B(n11587), .Z(n11589) );
  XNOR U11485 ( .A(n11406), .B(n11583), .Z(n11585) );
  XOR U11486 ( .A(n11591), .B(n11592), .Z(n11406) );
  AND U11487 ( .A(n312), .B(n11593), .Z(n11592) );
  XOR U11488 ( .A(n11594), .B(n11591), .Z(n11593) );
  XOR U11489 ( .A(n11595), .B(n11596), .Z(n11583) );
  AND U11490 ( .A(n11597), .B(n11598), .Z(n11596) );
  XOR U11491 ( .A(n11595), .B(n11421), .Z(n11598) );
  XOR U11492 ( .A(n11599), .B(n11600), .Z(n11421) );
  AND U11493 ( .A(n314), .B(n11601), .Z(n11600) );
  XOR U11494 ( .A(n11602), .B(n11599), .Z(n11601) );
  XNOR U11495 ( .A(n11418), .B(n11595), .Z(n11597) );
  XOR U11496 ( .A(n11603), .B(n11604), .Z(n11418) );
  AND U11497 ( .A(n312), .B(n11605), .Z(n11604) );
  XOR U11498 ( .A(n11606), .B(n11603), .Z(n11605) );
  XOR U11499 ( .A(n11607), .B(n11608), .Z(n11595) );
  AND U11500 ( .A(n11609), .B(n11610), .Z(n11608) );
  XOR U11501 ( .A(n11607), .B(n11433), .Z(n11610) );
  XOR U11502 ( .A(n11611), .B(n11612), .Z(n11433) );
  AND U11503 ( .A(n314), .B(n11613), .Z(n11612) );
  XOR U11504 ( .A(n11614), .B(n11611), .Z(n11613) );
  XNOR U11505 ( .A(n11430), .B(n11607), .Z(n11609) );
  XOR U11506 ( .A(n11615), .B(n11616), .Z(n11430) );
  AND U11507 ( .A(n312), .B(n11617), .Z(n11616) );
  XOR U11508 ( .A(n11618), .B(n11615), .Z(n11617) );
  XOR U11509 ( .A(n11619), .B(n11620), .Z(n11607) );
  AND U11510 ( .A(n11621), .B(n11622), .Z(n11620) );
  XOR U11511 ( .A(n11619), .B(n11445), .Z(n11622) );
  XOR U11512 ( .A(n11623), .B(n11624), .Z(n11445) );
  AND U11513 ( .A(n314), .B(n11625), .Z(n11624) );
  XOR U11514 ( .A(n11626), .B(n11623), .Z(n11625) );
  XNOR U11515 ( .A(n11442), .B(n11619), .Z(n11621) );
  XOR U11516 ( .A(n11627), .B(n11628), .Z(n11442) );
  AND U11517 ( .A(n312), .B(n11629), .Z(n11628) );
  XOR U11518 ( .A(n11630), .B(n11627), .Z(n11629) );
  XOR U11519 ( .A(n11631), .B(n11632), .Z(n11619) );
  AND U11520 ( .A(n11633), .B(n11634), .Z(n11632) );
  XOR U11521 ( .A(n11631), .B(n11457), .Z(n11634) );
  XOR U11522 ( .A(n11635), .B(n11636), .Z(n11457) );
  AND U11523 ( .A(n314), .B(n11637), .Z(n11636) );
  XOR U11524 ( .A(n11638), .B(n11635), .Z(n11637) );
  XNOR U11525 ( .A(n11454), .B(n11631), .Z(n11633) );
  XOR U11526 ( .A(n11639), .B(n11640), .Z(n11454) );
  AND U11527 ( .A(n312), .B(n11641), .Z(n11640) );
  XOR U11528 ( .A(n11642), .B(n11639), .Z(n11641) );
  XOR U11529 ( .A(n11643), .B(n11644), .Z(n11631) );
  AND U11530 ( .A(n11645), .B(n11646), .Z(n11644) );
  XOR U11531 ( .A(n11643), .B(n11469), .Z(n11646) );
  XOR U11532 ( .A(n11647), .B(n11648), .Z(n11469) );
  AND U11533 ( .A(n314), .B(n11649), .Z(n11648) );
  XOR U11534 ( .A(n11650), .B(n11647), .Z(n11649) );
  XNOR U11535 ( .A(n11466), .B(n11643), .Z(n11645) );
  XOR U11536 ( .A(n11651), .B(n11652), .Z(n11466) );
  AND U11537 ( .A(n312), .B(n11653), .Z(n11652) );
  XOR U11538 ( .A(n11654), .B(n11651), .Z(n11653) );
  XOR U11539 ( .A(n11655), .B(n11656), .Z(n11643) );
  AND U11540 ( .A(n11657), .B(n11658), .Z(n11656) );
  XOR U11541 ( .A(n11655), .B(n11481), .Z(n11658) );
  XOR U11542 ( .A(n11659), .B(n11660), .Z(n11481) );
  AND U11543 ( .A(n314), .B(n11661), .Z(n11660) );
  XOR U11544 ( .A(n11662), .B(n11659), .Z(n11661) );
  XNOR U11545 ( .A(n11478), .B(n11655), .Z(n11657) );
  XOR U11546 ( .A(n11663), .B(n11664), .Z(n11478) );
  AND U11547 ( .A(n312), .B(n11665), .Z(n11664) );
  XOR U11548 ( .A(n11666), .B(n11663), .Z(n11665) );
  XOR U11549 ( .A(n11667), .B(n11668), .Z(n11655) );
  AND U11550 ( .A(n11669), .B(n11670), .Z(n11668) );
  XOR U11551 ( .A(n11667), .B(n11493), .Z(n11670) );
  XOR U11552 ( .A(n11671), .B(n11672), .Z(n11493) );
  AND U11553 ( .A(n314), .B(n11673), .Z(n11672) );
  XOR U11554 ( .A(n11674), .B(n11671), .Z(n11673) );
  XNOR U11555 ( .A(n11490), .B(n11667), .Z(n11669) );
  XOR U11556 ( .A(n11675), .B(n11676), .Z(n11490) );
  AND U11557 ( .A(n312), .B(n11677), .Z(n11676) );
  XOR U11558 ( .A(n11678), .B(n11675), .Z(n11677) );
  XOR U11559 ( .A(n11679), .B(n11680), .Z(n11667) );
  AND U11560 ( .A(n11681), .B(n11682), .Z(n11680) );
  XOR U11561 ( .A(n11679), .B(n11505), .Z(n11682) );
  XOR U11562 ( .A(n11683), .B(n11684), .Z(n11505) );
  AND U11563 ( .A(n314), .B(n11685), .Z(n11684) );
  XOR U11564 ( .A(n11686), .B(n11683), .Z(n11685) );
  XNOR U11565 ( .A(n11502), .B(n11679), .Z(n11681) );
  XOR U11566 ( .A(n11687), .B(n11688), .Z(n11502) );
  AND U11567 ( .A(n312), .B(n11689), .Z(n11688) );
  XOR U11568 ( .A(n11690), .B(n11687), .Z(n11689) );
  XOR U11569 ( .A(n11691), .B(n11692), .Z(n11679) );
  AND U11570 ( .A(n11693), .B(n11694), .Z(n11692) );
  XOR U11571 ( .A(n11691), .B(n11517), .Z(n11694) );
  XOR U11572 ( .A(n11695), .B(n11696), .Z(n11517) );
  AND U11573 ( .A(n314), .B(n11697), .Z(n11696) );
  XOR U11574 ( .A(n11698), .B(n11695), .Z(n11697) );
  XNOR U11575 ( .A(n11514), .B(n11691), .Z(n11693) );
  XOR U11576 ( .A(n11699), .B(n11700), .Z(n11514) );
  AND U11577 ( .A(n312), .B(n11701), .Z(n11700) );
  XOR U11578 ( .A(n11702), .B(n11699), .Z(n11701) );
  XOR U11579 ( .A(n11703), .B(n11704), .Z(n11691) );
  AND U11580 ( .A(n11705), .B(n11706), .Z(n11704) );
  XOR U11581 ( .A(n11703), .B(n11529), .Z(n11706) );
  XOR U11582 ( .A(n11707), .B(n11708), .Z(n11529) );
  AND U11583 ( .A(n314), .B(n11709), .Z(n11708) );
  XOR U11584 ( .A(n11710), .B(n11707), .Z(n11709) );
  XNOR U11585 ( .A(n11526), .B(n11703), .Z(n11705) );
  XOR U11586 ( .A(n11711), .B(n11712), .Z(n11526) );
  AND U11587 ( .A(n312), .B(n11713), .Z(n11712) );
  XOR U11588 ( .A(n11714), .B(n11711), .Z(n11713) );
  XOR U11589 ( .A(n11715), .B(n11716), .Z(n11703) );
  AND U11590 ( .A(n11717), .B(n11718), .Z(n11716) );
  XOR U11591 ( .A(n11541), .B(n11715), .Z(n11718) );
  XOR U11592 ( .A(n11719), .B(n11720), .Z(n11541) );
  AND U11593 ( .A(n314), .B(n11721), .Z(n11720) );
  XOR U11594 ( .A(n11719), .B(n11722), .Z(n11721) );
  XNOR U11595 ( .A(n11715), .B(n11538), .Z(n11717) );
  XOR U11596 ( .A(n11723), .B(n11724), .Z(n11538) );
  AND U11597 ( .A(n312), .B(n11725), .Z(n11724) );
  XOR U11598 ( .A(n11723), .B(n11726), .Z(n11725) );
  XOR U11599 ( .A(n11727), .B(n11728), .Z(n11715) );
  AND U11600 ( .A(n11729), .B(n11730), .Z(n11728) );
  XNOR U11601 ( .A(n11731), .B(n11554), .Z(n11730) );
  XOR U11602 ( .A(n11732), .B(n11733), .Z(n11554) );
  AND U11603 ( .A(n314), .B(n11734), .Z(n11733) );
  XOR U11604 ( .A(n11735), .B(n11732), .Z(n11734) );
  XNOR U11605 ( .A(n11551), .B(n11727), .Z(n11729) );
  XOR U11606 ( .A(n11736), .B(n11737), .Z(n11551) );
  AND U11607 ( .A(n312), .B(n11738), .Z(n11737) );
  XOR U11608 ( .A(n11739), .B(n11736), .Z(n11738) );
  IV U11609 ( .A(n11731), .Z(n11727) );
  AND U11610 ( .A(n11559), .B(n11562), .Z(n11731) );
  XNOR U11611 ( .A(n11740), .B(n11741), .Z(n11562) );
  AND U11612 ( .A(n314), .B(n11742), .Z(n11741) );
  XNOR U11613 ( .A(n11743), .B(n11740), .Z(n11742) );
  XOR U11614 ( .A(n11744), .B(n11745), .Z(n314) );
  AND U11615 ( .A(n11746), .B(n11747), .Z(n11745) );
  XNOR U11616 ( .A(n11567), .B(n11744), .Z(n11747) );
  AND U11617 ( .A(p_input[511]), .B(p_input[495]), .Z(n11567) );
  XOR U11618 ( .A(n11744), .B(n11568), .Z(n11746) );
  AND U11619 ( .A(p_input[479]), .B(p_input[463]), .Z(n11568) );
  XOR U11620 ( .A(n11748), .B(n11749), .Z(n11744) );
  AND U11621 ( .A(n11750), .B(n11751), .Z(n11749) );
  XOR U11622 ( .A(n11748), .B(n11578), .Z(n11751) );
  XNOR U11623 ( .A(p_input[494]), .B(n11752), .Z(n11578) );
  AND U11624 ( .A(n470), .B(n11753), .Z(n11752) );
  XOR U11625 ( .A(p_input[510]), .B(p_input[494]), .Z(n11753) );
  XNOR U11626 ( .A(n11575), .B(n11748), .Z(n11750) );
  XOR U11627 ( .A(n11754), .B(n11755), .Z(n11575) );
  AND U11628 ( .A(n468), .B(n11756), .Z(n11755) );
  XOR U11629 ( .A(p_input[478]), .B(p_input[462]), .Z(n11756) );
  XOR U11630 ( .A(n11757), .B(n11758), .Z(n11748) );
  AND U11631 ( .A(n11759), .B(n11760), .Z(n11758) );
  XOR U11632 ( .A(n11757), .B(n11590), .Z(n11760) );
  XNOR U11633 ( .A(p_input[493]), .B(n11761), .Z(n11590) );
  AND U11634 ( .A(n470), .B(n11762), .Z(n11761) );
  XOR U11635 ( .A(p_input[509]), .B(p_input[493]), .Z(n11762) );
  XNOR U11636 ( .A(n11587), .B(n11757), .Z(n11759) );
  XOR U11637 ( .A(n11763), .B(n11764), .Z(n11587) );
  AND U11638 ( .A(n468), .B(n11765), .Z(n11764) );
  XOR U11639 ( .A(p_input[477]), .B(p_input[461]), .Z(n11765) );
  XOR U11640 ( .A(n11766), .B(n11767), .Z(n11757) );
  AND U11641 ( .A(n11768), .B(n11769), .Z(n11767) );
  XOR U11642 ( .A(n11766), .B(n11602), .Z(n11769) );
  XNOR U11643 ( .A(p_input[492]), .B(n11770), .Z(n11602) );
  AND U11644 ( .A(n470), .B(n11771), .Z(n11770) );
  XOR U11645 ( .A(p_input[508]), .B(p_input[492]), .Z(n11771) );
  XNOR U11646 ( .A(n11599), .B(n11766), .Z(n11768) );
  XOR U11647 ( .A(n11772), .B(n11773), .Z(n11599) );
  AND U11648 ( .A(n468), .B(n11774), .Z(n11773) );
  XOR U11649 ( .A(p_input[476]), .B(p_input[460]), .Z(n11774) );
  XOR U11650 ( .A(n11775), .B(n11776), .Z(n11766) );
  AND U11651 ( .A(n11777), .B(n11778), .Z(n11776) );
  XOR U11652 ( .A(n11775), .B(n11614), .Z(n11778) );
  XNOR U11653 ( .A(p_input[491]), .B(n11779), .Z(n11614) );
  AND U11654 ( .A(n470), .B(n11780), .Z(n11779) );
  XOR U11655 ( .A(p_input[507]), .B(p_input[491]), .Z(n11780) );
  XNOR U11656 ( .A(n11611), .B(n11775), .Z(n11777) );
  XOR U11657 ( .A(n11781), .B(n11782), .Z(n11611) );
  AND U11658 ( .A(n468), .B(n11783), .Z(n11782) );
  XOR U11659 ( .A(p_input[475]), .B(p_input[459]), .Z(n11783) );
  XOR U11660 ( .A(n11784), .B(n11785), .Z(n11775) );
  AND U11661 ( .A(n11786), .B(n11787), .Z(n11785) );
  XOR U11662 ( .A(n11784), .B(n11626), .Z(n11787) );
  XNOR U11663 ( .A(p_input[490]), .B(n11788), .Z(n11626) );
  AND U11664 ( .A(n470), .B(n11789), .Z(n11788) );
  XOR U11665 ( .A(p_input[506]), .B(p_input[490]), .Z(n11789) );
  XNOR U11666 ( .A(n11623), .B(n11784), .Z(n11786) );
  XOR U11667 ( .A(n11790), .B(n11791), .Z(n11623) );
  AND U11668 ( .A(n468), .B(n11792), .Z(n11791) );
  XOR U11669 ( .A(p_input[474]), .B(p_input[458]), .Z(n11792) );
  XOR U11670 ( .A(n11793), .B(n11794), .Z(n11784) );
  AND U11671 ( .A(n11795), .B(n11796), .Z(n11794) );
  XOR U11672 ( .A(n11793), .B(n11638), .Z(n11796) );
  XNOR U11673 ( .A(p_input[489]), .B(n11797), .Z(n11638) );
  AND U11674 ( .A(n470), .B(n11798), .Z(n11797) );
  XOR U11675 ( .A(p_input[505]), .B(p_input[489]), .Z(n11798) );
  XNOR U11676 ( .A(n11635), .B(n11793), .Z(n11795) );
  XOR U11677 ( .A(n11799), .B(n11800), .Z(n11635) );
  AND U11678 ( .A(n468), .B(n11801), .Z(n11800) );
  XOR U11679 ( .A(p_input[473]), .B(p_input[457]), .Z(n11801) );
  XOR U11680 ( .A(n11802), .B(n11803), .Z(n11793) );
  AND U11681 ( .A(n11804), .B(n11805), .Z(n11803) );
  XOR U11682 ( .A(n11802), .B(n11650), .Z(n11805) );
  XNOR U11683 ( .A(p_input[488]), .B(n11806), .Z(n11650) );
  AND U11684 ( .A(n470), .B(n11807), .Z(n11806) );
  XOR U11685 ( .A(p_input[504]), .B(p_input[488]), .Z(n11807) );
  XNOR U11686 ( .A(n11647), .B(n11802), .Z(n11804) );
  XOR U11687 ( .A(n11808), .B(n11809), .Z(n11647) );
  AND U11688 ( .A(n468), .B(n11810), .Z(n11809) );
  XOR U11689 ( .A(p_input[472]), .B(p_input[456]), .Z(n11810) );
  XOR U11690 ( .A(n11811), .B(n11812), .Z(n11802) );
  AND U11691 ( .A(n11813), .B(n11814), .Z(n11812) );
  XOR U11692 ( .A(n11811), .B(n11662), .Z(n11814) );
  XNOR U11693 ( .A(p_input[487]), .B(n11815), .Z(n11662) );
  AND U11694 ( .A(n470), .B(n11816), .Z(n11815) );
  XOR U11695 ( .A(p_input[503]), .B(p_input[487]), .Z(n11816) );
  XNOR U11696 ( .A(n11659), .B(n11811), .Z(n11813) );
  XOR U11697 ( .A(n11817), .B(n11818), .Z(n11659) );
  AND U11698 ( .A(n468), .B(n11819), .Z(n11818) );
  XOR U11699 ( .A(p_input[471]), .B(p_input[455]), .Z(n11819) );
  XOR U11700 ( .A(n11820), .B(n11821), .Z(n11811) );
  AND U11701 ( .A(n11822), .B(n11823), .Z(n11821) );
  XOR U11702 ( .A(n11820), .B(n11674), .Z(n11823) );
  XNOR U11703 ( .A(p_input[486]), .B(n11824), .Z(n11674) );
  AND U11704 ( .A(n470), .B(n11825), .Z(n11824) );
  XOR U11705 ( .A(p_input[502]), .B(p_input[486]), .Z(n11825) );
  XNOR U11706 ( .A(n11671), .B(n11820), .Z(n11822) );
  XOR U11707 ( .A(n11826), .B(n11827), .Z(n11671) );
  AND U11708 ( .A(n468), .B(n11828), .Z(n11827) );
  XOR U11709 ( .A(p_input[470]), .B(p_input[454]), .Z(n11828) );
  XOR U11710 ( .A(n11829), .B(n11830), .Z(n11820) );
  AND U11711 ( .A(n11831), .B(n11832), .Z(n11830) );
  XOR U11712 ( .A(n11829), .B(n11686), .Z(n11832) );
  XNOR U11713 ( .A(p_input[485]), .B(n11833), .Z(n11686) );
  AND U11714 ( .A(n470), .B(n11834), .Z(n11833) );
  XOR U11715 ( .A(p_input[501]), .B(p_input[485]), .Z(n11834) );
  XNOR U11716 ( .A(n11683), .B(n11829), .Z(n11831) );
  XOR U11717 ( .A(n11835), .B(n11836), .Z(n11683) );
  AND U11718 ( .A(n468), .B(n11837), .Z(n11836) );
  XOR U11719 ( .A(p_input[469]), .B(p_input[453]), .Z(n11837) );
  XOR U11720 ( .A(n11838), .B(n11839), .Z(n11829) );
  AND U11721 ( .A(n11840), .B(n11841), .Z(n11839) );
  XOR U11722 ( .A(n11838), .B(n11698), .Z(n11841) );
  XNOR U11723 ( .A(p_input[484]), .B(n11842), .Z(n11698) );
  AND U11724 ( .A(n470), .B(n11843), .Z(n11842) );
  XOR U11725 ( .A(p_input[500]), .B(p_input[484]), .Z(n11843) );
  XNOR U11726 ( .A(n11695), .B(n11838), .Z(n11840) );
  XOR U11727 ( .A(n11844), .B(n11845), .Z(n11695) );
  AND U11728 ( .A(n468), .B(n11846), .Z(n11845) );
  XOR U11729 ( .A(p_input[468]), .B(p_input[452]), .Z(n11846) );
  XOR U11730 ( .A(n11847), .B(n11848), .Z(n11838) );
  AND U11731 ( .A(n11849), .B(n11850), .Z(n11848) );
  XOR U11732 ( .A(n11847), .B(n11710), .Z(n11850) );
  XNOR U11733 ( .A(p_input[483]), .B(n11851), .Z(n11710) );
  AND U11734 ( .A(n470), .B(n11852), .Z(n11851) );
  XOR U11735 ( .A(p_input[499]), .B(p_input[483]), .Z(n11852) );
  XNOR U11736 ( .A(n11707), .B(n11847), .Z(n11849) );
  XOR U11737 ( .A(n11853), .B(n11854), .Z(n11707) );
  AND U11738 ( .A(n468), .B(n11855), .Z(n11854) );
  XOR U11739 ( .A(p_input[467]), .B(p_input[451]), .Z(n11855) );
  XOR U11740 ( .A(n11856), .B(n11857), .Z(n11847) );
  AND U11741 ( .A(n11858), .B(n11859), .Z(n11857) );
  XOR U11742 ( .A(n11722), .B(n11856), .Z(n11859) );
  XNOR U11743 ( .A(p_input[482]), .B(n11860), .Z(n11722) );
  AND U11744 ( .A(n470), .B(n11861), .Z(n11860) );
  XOR U11745 ( .A(p_input[498]), .B(p_input[482]), .Z(n11861) );
  XNOR U11746 ( .A(n11856), .B(n11719), .Z(n11858) );
  XOR U11747 ( .A(n11862), .B(n11863), .Z(n11719) );
  AND U11748 ( .A(n468), .B(n11864), .Z(n11863) );
  XOR U11749 ( .A(p_input[466]), .B(p_input[450]), .Z(n11864) );
  XOR U11750 ( .A(n11865), .B(n11866), .Z(n11856) );
  AND U11751 ( .A(n11867), .B(n11868), .Z(n11866) );
  XNOR U11752 ( .A(n11869), .B(n11735), .Z(n11868) );
  XNOR U11753 ( .A(p_input[481]), .B(n11870), .Z(n11735) );
  AND U11754 ( .A(n470), .B(n11871), .Z(n11870) );
  XNOR U11755 ( .A(p_input[497]), .B(n11872), .Z(n11871) );
  IV U11756 ( .A(p_input[481]), .Z(n11872) );
  XNOR U11757 ( .A(n11732), .B(n11865), .Z(n11867) );
  XNOR U11758 ( .A(p_input[449]), .B(n11873), .Z(n11732) );
  AND U11759 ( .A(n468), .B(n11874), .Z(n11873) );
  XOR U11760 ( .A(p_input[465]), .B(p_input[449]), .Z(n11874) );
  IV U11761 ( .A(n11869), .Z(n11865) );
  AND U11762 ( .A(n11740), .B(n11743), .Z(n11869) );
  XOR U11763 ( .A(p_input[480]), .B(n11875), .Z(n11743) );
  AND U11764 ( .A(n470), .B(n11876), .Z(n11875) );
  XOR U11765 ( .A(p_input[496]), .B(p_input[480]), .Z(n11876) );
  XOR U11766 ( .A(n11877), .B(n11878), .Z(n470) );
  AND U11767 ( .A(n11879), .B(n11880), .Z(n11878) );
  XNOR U11768 ( .A(p_input[511]), .B(n11877), .Z(n11880) );
  XOR U11769 ( .A(n11877), .B(p_input[495]), .Z(n11879) );
  XOR U11770 ( .A(n11881), .B(n11882), .Z(n11877) );
  AND U11771 ( .A(n11883), .B(n11884), .Z(n11882) );
  XNOR U11772 ( .A(p_input[510]), .B(n11881), .Z(n11884) );
  XOR U11773 ( .A(n11881), .B(p_input[494]), .Z(n11883) );
  XOR U11774 ( .A(n11885), .B(n11886), .Z(n11881) );
  AND U11775 ( .A(n11887), .B(n11888), .Z(n11886) );
  XNOR U11776 ( .A(p_input[509]), .B(n11885), .Z(n11888) );
  XOR U11777 ( .A(n11885), .B(p_input[493]), .Z(n11887) );
  XOR U11778 ( .A(n11889), .B(n11890), .Z(n11885) );
  AND U11779 ( .A(n11891), .B(n11892), .Z(n11890) );
  XNOR U11780 ( .A(p_input[508]), .B(n11889), .Z(n11892) );
  XOR U11781 ( .A(n11889), .B(p_input[492]), .Z(n11891) );
  XOR U11782 ( .A(n11893), .B(n11894), .Z(n11889) );
  AND U11783 ( .A(n11895), .B(n11896), .Z(n11894) );
  XNOR U11784 ( .A(p_input[507]), .B(n11893), .Z(n11896) );
  XOR U11785 ( .A(n11893), .B(p_input[491]), .Z(n11895) );
  XOR U11786 ( .A(n11897), .B(n11898), .Z(n11893) );
  AND U11787 ( .A(n11899), .B(n11900), .Z(n11898) );
  XNOR U11788 ( .A(p_input[506]), .B(n11897), .Z(n11900) );
  XOR U11789 ( .A(n11897), .B(p_input[490]), .Z(n11899) );
  XOR U11790 ( .A(n11901), .B(n11902), .Z(n11897) );
  AND U11791 ( .A(n11903), .B(n11904), .Z(n11902) );
  XNOR U11792 ( .A(p_input[505]), .B(n11901), .Z(n11904) );
  XOR U11793 ( .A(n11901), .B(p_input[489]), .Z(n11903) );
  XOR U11794 ( .A(n11905), .B(n11906), .Z(n11901) );
  AND U11795 ( .A(n11907), .B(n11908), .Z(n11906) );
  XNOR U11796 ( .A(p_input[504]), .B(n11905), .Z(n11908) );
  XOR U11797 ( .A(n11905), .B(p_input[488]), .Z(n11907) );
  XOR U11798 ( .A(n11909), .B(n11910), .Z(n11905) );
  AND U11799 ( .A(n11911), .B(n11912), .Z(n11910) );
  XNOR U11800 ( .A(p_input[503]), .B(n11909), .Z(n11912) );
  XOR U11801 ( .A(n11909), .B(p_input[487]), .Z(n11911) );
  XOR U11802 ( .A(n11913), .B(n11914), .Z(n11909) );
  AND U11803 ( .A(n11915), .B(n11916), .Z(n11914) );
  XNOR U11804 ( .A(p_input[502]), .B(n11913), .Z(n11916) );
  XOR U11805 ( .A(n11913), .B(p_input[486]), .Z(n11915) );
  XOR U11806 ( .A(n11917), .B(n11918), .Z(n11913) );
  AND U11807 ( .A(n11919), .B(n11920), .Z(n11918) );
  XNOR U11808 ( .A(p_input[501]), .B(n11917), .Z(n11920) );
  XOR U11809 ( .A(n11917), .B(p_input[485]), .Z(n11919) );
  XOR U11810 ( .A(n11921), .B(n11922), .Z(n11917) );
  AND U11811 ( .A(n11923), .B(n11924), .Z(n11922) );
  XNOR U11812 ( .A(p_input[500]), .B(n11921), .Z(n11924) );
  XOR U11813 ( .A(n11921), .B(p_input[484]), .Z(n11923) );
  XOR U11814 ( .A(n11925), .B(n11926), .Z(n11921) );
  AND U11815 ( .A(n11927), .B(n11928), .Z(n11926) );
  XNOR U11816 ( .A(p_input[499]), .B(n11925), .Z(n11928) );
  XOR U11817 ( .A(n11925), .B(p_input[483]), .Z(n11927) );
  XOR U11818 ( .A(n11929), .B(n11930), .Z(n11925) );
  AND U11819 ( .A(n11931), .B(n11932), .Z(n11930) );
  XNOR U11820 ( .A(p_input[498]), .B(n11929), .Z(n11932) );
  XOR U11821 ( .A(n11929), .B(p_input[482]), .Z(n11931) );
  XNOR U11822 ( .A(n11933), .B(n11934), .Z(n11929) );
  AND U11823 ( .A(n11935), .B(n11936), .Z(n11934) );
  XOR U11824 ( .A(p_input[497]), .B(n11933), .Z(n11936) );
  XNOR U11825 ( .A(p_input[481]), .B(n11933), .Z(n11935) );
  AND U11826 ( .A(p_input[496]), .B(n11937), .Z(n11933) );
  IV U11827 ( .A(p_input[480]), .Z(n11937) );
  XNOR U11828 ( .A(p_input[448]), .B(n11938), .Z(n11740) );
  AND U11829 ( .A(n468), .B(n11939), .Z(n11938) );
  XOR U11830 ( .A(p_input[464]), .B(p_input[448]), .Z(n11939) );
  XOR U11831 ( .A(n11940), .B(n11941), .Z(n468) );
  AND U11832 ( .A(n11942), .B(n11943), .Z(n11941) );
  XNOR U11833 ( .A(p_input[479]), .B(n11940), .Z(n11943) );
  XOR U11834 ( .A(n11940), .B(p_input[463]), .Z(n11942) );
  XOR U11835 ( .A(n11944), .B(n11945), .Z(n11940) );
  AND U11836 ( .A(n11946), .B(n11947), .Z(n11945) );
  XNOR U11837 ( .A(p_input[478]), .B(n11944), .Z(n11947) );
  XNOR U11838 ( .A(n11944), .B(n11754), .Z(n11946) );
  IV U11839 ( .A(p_input[462]), .Z(n11754) );
  XOR U11840 ( .A(n11948), .B(n11949), .Z(n11944) );
  AND U11841 ( .A(n11950), .B(n11951), .Z(n11949) );
  XNOR U11842 ( .A(p_input[477]), .B(n11948), .Z(n11951) );
  XNOR U11843 ( .A(n11948), .B(n11763), .Z(n11950) );
  IV U11844 ( .A(p_input[461]), .Z(n11763) );
  XOR U11845 ( .A(n11952), .B(n11953), .Z(n11948) );
  AND U11846 ( .A(n11954), .B(n11955), .Z(n11953) );
  XNOR U11847 ( .A(p_input[476]), .B(n11952), .Z(n11955) );
  XNOR U11848 ( .A(n11952), .B(n11772), .Z(n11954) );
  IV U11849 ( .A(p_input[460]), .Z(n11772) );
  XOR U11850 ( .A(n11956), .B(n11957), .Z(n11952) );
  AND U11851 ( .A(n11958), .B(n11959), .Z(n11957) );
  XNOR U11852 ( .A(p_input[475]), .B(n11956), .Z(n11959) );
  XNOR U11853 ( .A(n11956), .B(n11781), .Z(n11958) );
  IV U11854 ( .A(p_input[459]), .Z(n11781) );
  XOR U11855 ( .A(n11960), .B(n11961), .Z(n11956) );
  AND U11856 ( .A(n11962), .B(n11963), .Z(n11961) );
  XNOR U11857 ( .A(p_input[474]), .B(n11960), .Z(n11963) );
  XNOR U11858 ( .A(n11960), .B(n11790), .Z(n11962) );
  IV U11859 ( .A(p_input[458]), .Z(n11790) );
  XOR U11860 ( .A(n11964), .B(n11965), .Z(n11960) );
  AND U11861 ( .A(n11966), .B(n11967), .Z(n11965) );
  XNOR U11862 ( .A(p_input[473]), .B(n11964), .Z(n11967) );
  XNOR U11863 ( .A(n11964), .B(n11799), .Z(n11966) );
  IV U11864 ( .A(p_input[457]), .Z(n11799) );
  XOR U11865 ( .A(n11968), .B(n11969), .Z(n11964) );
  AND U11866 ( .A(n11970), .B(n11971), .Z(n11969) );
  XNOR U11867 ( .A(p_input[472]), .B(n11968), .Z(n11971) );
  XNOR U11868 ( .A(n11968), .B(n11808), .Z(n11970) );
  IV U11869 ( .A(p_input[456]), .Z(n11808) );
  XOR U11870 ( .A(n11972), .B(n11973), .Z(n11968) );
  AND U11871 ( .A(n11974), .B(n11975), .Z(n11973) );
  XNOR U11872 ( .A(p_input[471]), .B(n11972), .Z(n11975) );
  XNOR U11873 ( .A(n11972), .B(n11817), .Z(n11974) );
  IV U11874 ( .A(p_input[455]), .Z(n11817) );
  XOR U11875 ( .A(n11976), .B(n11977), .Z(n11972) );
  AND U11876 ( .A(n11978), .B(n11979), .Z(n11977) );
  XNOR U11877 ( .A(p_input[470]), .B(n11976), .Z(n11979) );
  XNOR U11878 ( .A(n11976), .B(n11826), .Z(n11978) );
  IV U11879 ( .A(p_input[454]), .Z(n11826) );
  XOR U11880 ( .A(n11980), .B(n11981), .Z(n11976) );
  AND U11881 ( .A(n11982), .B(n11983), .Z(n11981) );
  XNOR U11882 ( .A(p_input[469]), .B(n11980), .Z(n11983) );
  XNOR U11883 ( .A(n11980), .B(n11835), .Z(n11982) );
  IV U11884 ( .A(p_input[453]), .Z(n11835) );
  XOR U11885 ( .A(n11984), .B(n11985), .Z(n11980) );
  AND U11886 ( .A(n11986), .B(n11987), .Z(n11985) );
  XNOR U11887 ( .A(p_input[468]), .B(n11984), .Z(n11987) );
  XNOR U11888 ( .A(n11984), .B(n11844), .Z(n11986) );
  IV U11889 ( .A(p_input[452]), .Z(n11844) );
  XOR U11890 ( .A(n11988), .B(n11989), .Z(n11984) );
  AND U11891 ( .A(n11990), .B(n11991), .Z(n11989) );
  XNOR U11892 ( .A(p_input[467]), .B(n11988), .Z(n11991) );
  XNOR U11893 ( .A(n11988), .B(n11853), .Z(n11990) );
  IV U11894 ( .A(p_input[451]), .Z(n11853) );
  XOR U11895 ( .A(n11992), .B(n11993), .Z(n11988) );
  AND U11896 ( .A(n11994), .B(n11995), .Z(n11993) );
  XNOR U11897 ( .A(p_input[466]), .B(n11992), .Z(n11995) );
  XNOR U11898 ( .A(n11992), .B(n11862), .Z(n11994) );
  IV U11899 ( .A(p_input[450]), .Z(n11862) );
  XNOR U11900 ( .A(n11996), .B(n11997), .Z(n11992) );
  AND U11901 ( .A(n11998), .B(n11999), .Z(n11997) );
  XOR U11902 ( .A(p_input[465]), .B(n11996), .Z(n11999) );
  XNOR U11903 ( .A(p_input[449]), .B(n11996), .Z(n11998) );
  AND U11904 ( .A(p_input[464]), .B(n12000), .Z(n11996) );
  IV U11905 ( .A(p_input[448]), .Z(n12000) );
  XOR U11906 ( .A(n12001), .B(n12002), .Z(n11559) );
  AND U11907 ( .A(n312), .B(n12003), .Z(n12002) );
  XNOR U11908 ( .A(n12004), .B(n12001), .Z(n12003) );
  XOR U11909 ( .A(n12005), .B(n12006), .Z(n312) );
  AND U11910 ( .A(n12007), .B(n12008), .Z(n12006) );
  XNOR U11911 ( .A(n11569), .B(n12005), .Z(n12008) );
  AND U11912 ( .A(p_input[447]), .B(p_input[431]), .Z(n11569) );
  XOR U11913 ( .A(n12005), .B(n11570), .Z(n12007) );
  AND U11914 ( .A(p_input[415]), .B(p_input[399]), .Z(n11570) );
  XOR U11915 ( .A(n12009), .B(n12010), .Z(n12005) );
  AND U11916 ( .A(n12011), .B(n12012), .Z(n12010) );
  XOR U11917 ( .A(n12009), .B(n11582), .Z(n12012) );
  XNOR U11918 ( .A(p_input[430]), .B(n12013), .Z(n11582) );
  AND U11919 ( .A(n474), .B(n12014), .Z(n12013) );
  XOR U11920 ( .A(p_input[446]), .B(p_input[430]), .Z(n12014) );
  XNOR U11921 ( .A(n11579), .B(n12009), .Z(n12011) );
  XOR U11922 ( .A(n12015), .B(n12016), .Z(n11579) );
  AND U11923 ( .A(n471), .B(n12017), .Z(n12016) );
  XOR U11924 ( .A(p_input[414]), .B(p_input[398]), .Z(n12017) );
  XOR U11925 ( .A(n12018), .B(n12019), .Z(n12009) );
  AND U11926 ( .A(n12020), .B(n12021), .Z(n12019) );
  XOR U11927 ( .A(n12018), .B(n11594), .Z(n12021) );
  XNOR U11928 ( .A(p_input[429]), .B(n12022), .Z(n11594) );
  AND U11929 ( .A(n474), .B(n12023), .Z(n12022) );
  XOR U11930 ( .A(p_input[445]), .B(p_input[429]), .Z(n12023) );
  XNOR U11931 ( .A(n11591), .B(n12018), .Z(n12020) );
  XOR U11932 ( .A(n12024), .B(n12025), .Z(n11591) );
  AND U11933 ( .A(n471), .B(n12026), .Z(n12025) );
  XOR U11934 ( .A(p_input[413]), .B(p_input[397]), .Z(n12026) );
  XOR U11935 ( .A(n12027), .B(n12028), .Z(n12018) );
  AND U11936 ( .A(n12029), .B(n12030), .Z(n12028) );
  XOR U11937 ( .A(n12027), .B(n11606), .Z(n12030) );
  XNOR U11938 ( .A(p_input[428]), .B(n12031), .Z(n11606) );
  AND U11939 ( .A(n474), .B(n12032), .Z(n12031) );
  XOR U11940 ( .A(p_input[444]), .B(p_input[428]), .Z(n12032) );
  XNOR U11941 ( .A(n11603), .B(n12027), .Z(n12029) );
  XOR U11942 ( .A(n12033), .B(n12034), .Z(n11603) );
  AND U11943 ( .A(n471), .B(n12035), .Z(n12034) );
  XOR U11944 ( .A(p_input[412]), .B(p_input[396]), .Z(n12035) );
  XOR U11945 ( .A(n12036), .B(n12037), .Z(n12027) );
  AND U11946 ( .A(n12038), .B(n12039), .Z(n12037) );
  XOR U11947 ( .A(n12036), .B(n11618), .Z(n12039) );
  XNOR U11948 ( .A(p_input[427]), .B(n12040), .Z(n11618) );
  AND U11949 ( .A(n474), .B(n12041), .Z(n12040) );
  XOR U11950 ( .A(p_input[443]), .B(p_input[427]), .Z(n12041) );
  XNOR U11951 ( .A(n11615), .B(n12036), .Z(n12038) );
  XOR U11952 ( .A(n12042), .B(n12043), .Z(n11615) );
  AND U11953 ( .A(n471), .B(n12044), .Z(n12043) );
  XOR U11954 ( .A(p_input[411]), .B(p_input[395]), .Z(n12044) );
  XOR U11955 ( .A(n12045), .B(n12046), .Z(n12036) );
  AND U11956 ( .A(n12047), .B(n12048), .Z(n12046) );
  XOR U11957 ( .A(n12045), .B(n11630), .Z(n12048) );
  XNOR U11958 ( .A(p_input[426]), .B(n12049), .Z(n11630) );
  AND U11959 ( .A(n474), .B(n12050), .Z(n12049) );
  XOR U11960 ( .A(p_input[442]), .B(p_input[426]), .Z(n12050) );
  XNOR U11961 ( .A(n11627), .B(n12045), .Z(n12047) );
  XOR U11962 ( .A(n12051), .B(n12052), .Z(n11627) );
  AND U11963 ( .A(n471), .B(n12053), .Z(n12052) );
  XOR U11964 ( .A(p_input[410]), .B(p_input[394]), .Z(n12053) );
  XOR U11965 ( .A(n12054), .B(n12055), .Z(n12045) );
  AND U11966 ( .A(n12056), .B(n12057), .Z(n12055) );
  XOR U11967 ( .A(n12054), .B(n11642), .Z(n12057) );
  XNOR U11968 ( .A(p_input[425]), .B(n12058), .Z(n11642) );
  AND U11969 ( .A(n474), .B(n12059), .Z(n12058) );
  XOR U11970 ( .A(p_input[441]), .B(p_input[425]), .Z(n12059) );
  XNOR U11971 ( .A(n11639), .B(n12054), .Z(n12056) );
  XOR U11972 ( .A(n12060), .B(n12061), .Z(n11639) );
  AND U11973 ( .A(n471), .B(n12062), .Z(n12061) );
  XOR U11974 ( .A(p_input[409]), .B(p_input[393]), .Z(n12062) );
  XOR U11975 ( .A(n12063), .B(n12064), .Z(n12054) );
  AND U11976 ( .A(n12065), .B(n12066), .Z(n12064) );
  XOR U11977 ( .A(n12063), .B(n11654), .Z(n12066) );
  XNOR U11978 ( .A(p_input[424]), .B(n12067), .Z(n11654) );
  AND U11979 ( .A(n474), .B(n12068), .Z(n12067) );
  XOR U11980 ( .A(p_input[440]), .B(p_input[424]), .Z(n12068) );
  XNOR U11981 ( .A(n11651), .B(n12063), .Z(n12065) );
  XOR U11982 ( .A(n12069), .B(n12070), .Z(n11651) );
  AND U11983 ( .A(n471), .B(n12071), .Z(n12070) );
  XOR U11984 ( .A(p_input[408]), .B(p_input[392]), .Z(n12071) );
  XOR U11985 ( .A(n12072), .B(n12073), .Z(n12063) );
  AND U11986 ( .A(n12074), .B(n12075), .Z(n12073) );
  XOR U11987 ( .A(n12072), .B(n11666), .Z(n12075) );
  XNOR U11988 ( .A(p_input[423]), .B(n12076), .Z(n11666) );
  AND U11989 ( .A(n474), .B(n12077), .Z(n12076) );
  XOR U11990 ( .A(p_input[439]), .B(p_input[423]), .Z(n12077) );
  XNOR U11991 ( .A(n11663), .B(n12072), .Z(n12074) );
  XOR U11992 ( .A(n12078), .B(n12079), .Z(n11663) );
  AND U11993 ( .A(n471), .B(n12080), .Z(n12079) );
  XOR U11994 ( .A(p_input[407]), .B(p_input[391]), .Z(n12080) );
  XOR U11995 ( .A(n12081), .B(n12082), .Z(n12072) );
  AND U11996 ( .A(n12083), .B(n12084), .Z(n12082) );
  XOR U11997 ( .A(n12081), .B(n11678), .Z(n12084) );
  XNOR U11998 ( .A(p_input[422]), .B(n12085), .Z(n11678) );
  AND U11999 ( .A(n474), .B(n12086), .Z(n12085) );
  XOR U12000 ( .A(p_input[438]), .B(p_input[422]), .Z(n12086) );
  XNOR U12001 ( .A(n11675), .B(n12081), .Z(n12083) );
  XOR U12002 ( .A(n12087), .B(n12088), .Z(n11675) );
  AND U12003 ( .A(n471), .B(n12089), .Z(n12088) );
  XOR U12004 ( .A(p_input[406]), .B(p_input[390]), .Z(n12089) );
  XOR U12005 ( .A(n12090), .B(n12091), .Z(n12081) );
  AND U12006 ( .A(n12092), .B(n12093), .Z(n12091) );
  XOR U12007 ( .A(n12090), .B(n11690), .Z(n12093) );
  XNOR U12008 ( .A(p_input[421]), .B(n12094), .Z(n11690) );
  AND U12009 ( .A(n474), .B(n12095), .Z(n12094) );
  XOR U12010 ( .A(p_input[437]), .B(p_input[421]), .Z(n12095) );
  XNOR U12011 ( .A(n11687), .B(n12090), .Z(n12092) );
  XOR U12012 ( .A(n12096), .B(n12097), .Z(n11687) );
  AND U12013 ( .A(n471), .B(n12098), .Z(n12097) );
  XOR U12014 ( .A(p_input[405]), .B(p_input[389]), .Z(n12098) );
  XOR U12015 ( .A(n12099), .B(n12100), .Z(n12090) );
  AND U12016 ( .A(n12101), .B(n12102), .Z(n12100) );
  XOR U12017 ( .A(n12099), .B(n11702), .Z(n12102) );
  XNOR U12018 ( .A(p_input[420]), .B(n12103), .Z(n11702) );
  AND U12019 ( .A(n474), .B(n12104), .Z(n12103) );
  XOR U12020 ( .A(p_input[436]), .B(p_input[420]), .Z(n12104) );
  XNOR U12021 ( .A(n11699), .B(n12099), .Z(n12101) );
  XOR U12022 ( .A(n12105), .B(n12106), .Z(n11699) );
  AND U12023 ( .A(n471), .B(n12107), .Z(n12106) );
  XOR U12024 ( .A(p_input[404]), .B(p_input[388]), .Z(n12107) );
  XOR U12025 ( .A(n12108), .B(n12109), .Z(n12099) );
  AND U12026 ( .A(n12110), .B(n12111), .Z(n12109) );
  XOR U12027 ( .A(n12108), .B(n11714), .Z(n12111) );
  XNOR U12028 ( .A(p_input[419]), .B(n12112), .Z(n11714) );
  AND U12029 ( .A(n474), .B(n12113), .Z(n12112) );
  XOR U12030 ( .A(p_input[435]), .B(p_input[419]), .Z(n12113) );
  XNOR U12031 ( .A(n11711), .B(n12108), .Z(n12110) );
  XOR U12032 ( .A(n12114), .B(n12115), .Z(n11711) );
  AND U12033 ( .A(n471), .B(n12116), .Z(n12115) );
  XOR U12034 ( .A(p_input[403]), .B(p_input[387]), .Z(n12116) );
  XOR U12035 ( .A(n12117), .B(n12118), .Z(n12108) );
  AND U12036 ( .A(n12119), .B(n12120), .Z(n12118) );
  XOR U12037 ( .A(n11726), .B(n12117), .Z(n12120) );
  XNOR U12038 ( .A(p_input[418]), .B(n12121), .Z(n11726) );
  AND U12039 ( .A(n474), .B(n12122), .Z(n12121) );
  XOR U12040 ( .A(p_input[434]), .B(p_input[418]), .Z(n12122) );
  XNOR U12041 ( .A(n12117), .B(n11723), .Z(n12119) );
  XOR U12042 ( .A(n12123), .B(n12124), .Z(n11723) );
  AND U12043 ( .A(n471), .B(n12125), .Z(n12124) );
  XOR U12044 ( .A(p_input[402]), .B(p_input[386]), .Z(n12125) );
  XOR U12045 ( .A(n12126), .B(n12127), .Z(n12117) );
  AND U12046 ( .A(n12128), .B(n12129), .Z(n12127) );
  XNOR U12047 ( .A(n12130), .B(n11739), .Z(n12129) );
  XNOR U12048 ( .A(p_input[417]), .B(n12131), .Z(n11739) );
  AND U12049 ( .A(n474), .B(n12132), .Z(n12131) );
  XNOR U12050 ( .A(p_input[433]), .B(n12133), .Z(n12132) );
  IV U12051 ( .A(p_input[417]), .Z(n12133) );
  XNOR U12052 ( .A(n11736), .B(n12126), .Z(n12128) );
  XNOR U12053 ( .A(p_input[385]), .B(n12134), .Z(n11736) );
  AND U12054 ( .A(n471), .B(n12135), .Z(n12134) );
  XOR U12055 ( .A(p_input[401]), .B(p_input[385]), .Z(n12135) );
  IV U12056 ( .A(n12130), .Z(n12126) );
  AND U12057 ( .A(n12001), .B(n12004), .Z(n12130) );
  XOR U12058 ( .A(p_input[416]), .B(n12136), .Z(n12004) );
  AND U12059 ( .A(n474), .B(n12137), .Z(n12136) );
  XOR U12060 ( .A(p_input[432]), .B(p_input[416]), .Z(n12137) );
  XOR U12061 ( .A(n12138), .B(n12139), .Z(n474) );
  AND U12062 ( .A(n12140), .B(n12141), .Z(n12139) );
  XNOR U12063 ( .A(p_input[447]), .B(n12138), .Z(n12141) );
  XOR U12064 ( .A(n12138), .B(p_input[431]), .Z(n12140) );
  XOR U12065 ( .A(n12142), .B(n12143), .Z(n12138) );
  AND U12066 ( .A(n12144), .B(n12145), .Z(n12143) );
  XNOR U12067 ( .A(p_input[446]), .B(n12142), .Z(n12145) );
  XOR U12068 ( .A(n12142), .B(p_input[430]), .Z(n12144) );
  XOR U12069 ( .A(n12146), .B(n12147), .Z(n12142) );
  AND U12070 ( .A(n12148), .B(n12149), .Z(n12147) );
  XNOR U12071 ( .A(p_input[445]), .B(n12146), .Z(n12149) );
  XOR U12072 ( .A(n12146), .B(p_input[429]), .Z(n12148) );
  XOR U12073 ( .A(n12150), .B(n12151), .Z(n12146) );
  AND U12074 ( .A(n12152), .B(n12153), .Z(n12151) );
  XNOR U12075 ( .A(p_input[444]), .B(n12150), .Z(n12153) );
  XOR U12076 ( .A(n12150), .B(p_input[428]), .Z(n12152) );
  XOR U12077 ( .A(n12154), .B(n12155), .Z(n12150) );
  AND U12078 ( .A(n12156), .B(n12157), .Z(n12155) );
  XNOR U12079 ( .A(p_input[443]), .B(n12154), .Z(n12157) );
  XOR U12080 ( .A(n12154), .B(p_input[427]), .Z(n12156) );
  XOR U12081 ( .A(n12158), .B(n12159), .Z(n12154) );
  AND U12082 ( .A(n12160), .B(n12161), .Z(n12159) );
  XNOR U12083 ( .A(p_input[442]), .B(n12158), .Z(n12161) );
  XOR U12084 ( .A(n12158), .B(p_input[426]), .Z(n12160) );
  XOR U12085 ( .A(n12162), .B(n12163), .Z(n12158) );
  AND U12086 ( .A(n12164), .B(n12165), .Z(n12163) );
  XNOR U12087 ( .A(p_input[441]), .B(n12162), .Z(n12165) );
  XOR U12088 ( .A(n12162), .B(p_input[425]), .Z(n12164) );
  XOR U12089 ( .A(n12166), .B(n12167), .Z(n12162) );
  AND U12090 ( .A(n12168), .B(n12169), .Z(n12167) );
  XNOR U12091 ( .A(p_input[440]), .B(n12166), .Z(n12169) );
  XOR U12092 ( .A(n12166), .B(p_input[424]), .Z(n12168) );
  XOR U12093 ( .A(n12170), .B(n12171), .Z(n12166) );
  AND U12094 ( .A(n12172), .B(n12173), .Z(n12171) );
  XNOR U12095 ( .A(p_input[439]), .B(n12170), .Z(n12173) );
  XOR U12096 ( .A(n12170), .B(p_input[423]), .Z(n12172) );
  XOR U12097 ( .A(n12174), .B(n12175), .Z(n12170) );
  AND U12098 ( .A(n12176), .B(n12177), .Z(n12175) );
  XNOR U12099 ( .A(p_input[438]), .B(n12174), .Z(n12177) );
  XOR U12100 ( .A(n12174), .B(p_input[422]), .Z(n12176) );
  XOR U12101 ( .A(n12178), .B(n12179), .Z(n12174) );
  AND U12102 ( .A(n12180), .B(n12181), .Z(n12179) );
  XNOR U12103 ( .A(p_input[437]), .B(n12178), .Z(n12181) );
  XOR U12104 ( .A(n12178), .B(p_input[421]), .Z(n12180) );
  XOR U12105 ( .A(n12182), .B(n12183), .Z(n12178) );
  AND U12106 ( .A(n12184), .B(n12185), .Z(n12183) );
  XNOR U12107 ( .A(p_input[436]), .B(n12182), .Z(n12185) );
  XOR U12108 ( .A(n12182), .B(p_input[420]), .Z(n12184) );
  XOR U12109 ( .A(n12186), .B(n12187), .Z(n12182) );
  AND U12110 ( .A(n12188), .B(n12189), .Z(n12187) );
  XNOR U12111 ( .A(p_input[435]), .B(n12186), .Z(n12189) );
  XOR U12112 ( .A(n12186), .B(p_input[419]), .Z(n12188) );
  XOR U12113 ( .A(n12190), .B(n12191), .Z(n12186) );
  AND U12114 ( .A(n12192), .B(n12193), .Z(n12191) );
  XNOR U12115 ( .A(p_input[434]), .B(n12190), .Z(n12193) );
  XOR U12116 ( .A(n12190), .B(p_input[418]), .Z(n12192) );
  XNOR U12117 ( .A(n12194), .B(n12195), .Z(n12190) );
  AND U12118 ( .A(n12196), .B(n12197), .Z(n12195) );
  XOR U12119 ( .A(p_input[433]), .B(n12194), .Z(n12197) );
  XNOR U12120 ( .A(p_input[417]), .B(n12194), .Z(n12196) );
  AND U12121 ( .A(p_input[432]), .B(n12198), .Z(n12194) );
  IV U12122 ( .A(p_input[416]), .Z(n12198) );
  XNOR U12123 ( .A(p_input[384]), .B(n12199), .Z(n12001) );
  AND U12124 ( .A(n471), .B(n12200), .Z(n12199) );
  XOR U12125 ( .A(p_input[400]), .B(p_input[384]), .Z(n12200) );
  XOR U12126 ( .A(n12201), .B(n12202), .Z(n471) );
  AND U12127 ( .A(n12203), .B(n12204), .Z(n12202) );
  XNOR U12128 ( .A(p_input[415]), .B(n12201), .Z(n12204) );
  XOR U12129 ( .A(n12201), .B(p_input[399]), .Z(n12203) );
  XOR U12130 ( .A(n12205), .B(n12206), .Z(n12201) );
  AND U12131 ( .A(n12207), .B(n12208), .Z(n12206) );
  XNOR U12132 ( .A(p_input[414]), .B(n12205), .Z(n12208) );
  XNOR U12133 ( .A(n12205), .B(n12015), .Z(n12207) );
  IV U12134 ( .A(p_input[398]), .Z(n12015) );
  XOR U12135 ( .A(n12209), .B(n12210), .Z(n12205) );
  AND U12136 ( .A(n12211), .B(n12212), .Z(n12210) );
  XNOR U12137 ( .A(p_input[413]), .B(n12209), .Z(n12212) );
  XNOR U12138 ( .A(n12209), .B(n12024), .Z(n12211) );
  IV U12139 ( .A(p_input[397]), .Z(n12024) );
  XOR U12140 ( .A(n12213), .B(n12214), .Z(n12209) );
  AND U12141 ( .A(n12215), .B(n12216), .Z(n12214) );
  XNOR U12142 ( .A(p_input[412]), .B(n12213), .Z(n12216) );
  XNOR U12143 ( .A(n12213), .B(n12033), .Z(n12215) );
  IV U12144 ( .A(p_input[396]), .Z(n12033) );
  XOR U12145 ( .A(n12217), .B(n12218), .Z(n12213) );
  AND U12146 ( .A(n12219), .B(n12220), .Z(n12218) );
  XNOR U12147 ( .A(p_input[411]), .B(n12217), .Z(n12220) );
  XNOR U12148 ( .A(n12217), .B(n12042), .Z(n12219) );
  IV U12149 ( .A(p_input[395]), .Z(n12042) );
  XOR U12150 ( .A(n12221), .B(n12222), .Z(n12217) );
  AND U12151 ( .A(n12223), .B(n12224), .Z(n12222) );
  XNOR U12152 ( .A(p_input[410]), .B(n12221), .Z(n12224) );
  XNOR U12153 ( .A(n12221), .B(n12051), .Z(n12223) );
  IV U12154 ( .A(p_input[394]), .Z(n12051) );
  XOR U12155 ( .A(n12225), .B(n12226), .Z(n12221) );
  AND U12156 ( .A(n12227), .B(n12228), .Z(n12226) );
  XNOR U12157 ( .A(p_input[409]), .B(n12225), .Z(n12228) );
  XNOR U12158 ( .A(n12225), .B(n12060), .Z(n12227) );
  IV U12159 ( .A(p_input[393]), .Z(n12060) );
  XOR U12160 ( .A(n12229), .B(n12230), .Z(n12225) );
  AND U12161 ( .A(n12231), .B(n12232), .Z(n12230) );
  XNOR U12162 ( .A(p_input[408]), .B(n12229), .Z(n12232) );
  XNOR U12163 ( .A(n12229), .B(n12069), .Z(n12231) );
  IV U12164 ( .A(p_input[392]), .Z(n12069) );
  XOR U12165 ( .A(n12233), .B(n12234), .Z(n12229) );
  AND U12166 ( .A(n12235), .B(n12236), .Z(n12234) );
  XNOR U12167 ( .A(p_input[407]), .B(n12233), .Z(n12236) );
  XNOR U12168 ( .A(n12233), .B(n12078), .Z(n12235) );
  IV U12169 ( .A(p_input[391]), .Z(n12078) );
  XOR U12170 ( .A(n12237), .B(n12238), .Z(n12233) );
  AND U12171 ( .A(n12239), .B(n12240), .Z(n12238) );
  XNOR U12172 ( .A(p_input[406]), .B(n12237), .Z(n12240) );
  XNOR U12173 ( .A(n12237), .B(n12087), .Z(n12239) );
  IV U12174 ( .A(p_input[390]), .Z(n12087) );
  XOR U12175 ( .A(n12241), .B(n12242), .Z(n12237) );
  AND U12176 ( .A(n12243), .B(n12244), .Z(n12242) );
  XNOR U12177 ( .A(p_input[405]), .B(n12241), .Z(n12244) );
  XNOR U12178 ( .A(n12241), .B(n12096), .Z(n12243) );
  IV U12179 ( .A(p_input[389]), .Z(n12096) );
  XOR U12180 ( .A(n12245), .B(n12246), .Z(n12241) );
  AND U12181 ( .A(n12247), .B(n12248), .Z(n12246) );
  XNOR U12182 ( .A(p_input[404]), .B(n12245), .Z(n12248) );
  XNOR U12183 ( .A(n12245), .B(n12105), .Z(n12247) );
  IV U12184 ( .A(p_input[388]), .Z(n12105) );
  XOR U12185 ( .A(n12249), .B(n12250), .Z(n12245) );
  AND U12186 ( .A(n12251), .B(n12252), .Z(n12250) );
  XNOR U12187 ( .A(p_input[403]), .B(n12249), .Z(n12252) );
  XNOR U12188 ( .A(n12249), .B(n12114), .Z(n12251) );
  IV U12189 ( .A(p_input[387]), .Z(n12114) );
  XOR U12190 ( .A(n12253), .B(n12254), .Z(n12249) );
  AND U12191 ( .A(n12255), .B(n12256), .Z(n12254) );
  XNOR U12192 ( .A(p_input[402]), .B(n12253), .Z(n12256) );
  XNOR U12193 ( .A(n12253), .B(n12123), .Z(n12255) );
  IV U12194 ( .A(p_input[386]), .Z(n12123) );
  XNOR U12195 ( .A(n12257), .B(n12258), .Z(n12253) );
  AND U12196 ( .A(n12259), .B(n12260), .Z(n12258) );
  XOR U12197 ( .A(p_input[401]), .B(n12257), .Z(n12260) );
  XNOR U12198 ( .A(p_input[385]), .B(n12257), .Z(n12259) );
  AND U12199 ( .A(p_input[400]), .B(n12261), .Z(n12257) );
  IV U12200 ( .A(p_input[384]), .Z(n12261) );
  XOR U12201 ( .A(n12262), .B(n12263), .Z(n11377) );
  AND U12202 ( .A(n448), .B(n12264), .Z(n12263) );
  XNOR U12203 ( .A(n12265), .B(n12262), .Z(n12264) );
  XOR U12204 ( .A(n12266), .B(n12267), .Z(n448) );
  AND U12205 ( .A(n12268), .B(n12269), .Z(n12267) );
  XNOR U12206 ( .A(n11389), .B(n12266), .Z(n12269) );
  AND U12207 ( .A(n12270), .B(n12271), .Z(n11389) );
  XOR U12208 ( .A(n12266), .B(n11388), .Z(n12268) );
  AND U12209 ( .A(n12272), .B(n12273), .Z(n11388) );
  XOR U12210 ( .A(n12274), .B(n12275), .Z(n12266) );
  AND U12211 ( .A(n12276), .B(n12277), .Z(n12275) );
  XOR U12212 ( .A(n12274), .B(n11401), .Z(n12277) );
  XOR U12213 ( .A(n12278), .B(n12279), .Z(n11401) );
  AND U12214 ( .A(n318), .B(n12280), .Z(n12279) );
  XOR U12215 ( .A(n12281), .B(n12278), .Z(n12280) );
  XNOR U12216 ( .A(n11398), .B(n12274), .Z(n12276) );
  XOR U12217 ( .A(n12282), .B(n12283), .Z(n11398) );
  AND U12218 ( .A(n315), .B(n12284), .Z(n12283) );
  XOR U12219 ( .A(n12285), .B(n12282), .Z(n12284) );
  XOR U12220 ( .A(n12286), .B(n12287), .Z(n12274) );
  AND U12221 ( .A(n12288), .B(n12289), .Z(n12287) );
  XOR U12222 ( .A(n12286), .B(n11413), .Z(n12289) );
  XOR U12223 ( .A(n12290), .B(n12291), .Z(n11413) );
  AND U12224 ( .A(n318), .B(n12292), .Z(n12291) );
  XOR U12225 ( .A(n12293), .B(n12290), .Z(n12292) );
  XNOR U12226 ( .A(n11410), .B(n12286), .Z(n12288) );
  XOR U12227 ( .A(n12294), .B(n12295), .Z(n11410) );
  AND U12228 ( .A(n315), .B(n12296), .Z(n12295) );
  XOR U12229 ( .A(n12297), .B(n12294), .Z(n12296) );
  XOR U12230 ( .A(n12298), .B(n12299), .Z(n12286) );
  AND U12231 ( .A(n12300), .B(n12301), .Z(n12299) );
  XOR U12232 ( .A(n12298), .B(n11425), .Z(n12301) );
  XOR U12233 ( .A(n12302), .B(n12303), .Z(n11425) );
  AND U12234 ( .A(n318), .B(n12304), .Z(n12303) );
  XOR U12235 ( .A(n12305), .B(n12302), .Z(n12304) );
  XNOR U12236 ( .A(n11422), .B(n12298), .Z(n12300) );
  XOR U12237 ( .A(n12306), .B(n12307), .Z(n11422) );
  AND U12238 ( .A(n315), .B(n12308), .Z(n12307) );
  XOR U12239 ( .A(n12309), .B(n12306), .Z(n12308) );
  XOR U12240 ( .A(n12310), .B(n12311), .Z(n12298) );
  AND U12241 ( .A(n12312), .B(n12313), .Z(n12311) );
  XOR U12242 ( .A(n12310), .B(n11437), .Z(n12313) );
  XOR U12243 ( .A(n12314), .B(n12315), .Z(n11437) );
  AND U12244 ( .A(n318), .B(n12316), .Z(n12315) );
  XOR U12245 ( .A(n12317), .B(n12314), .Z(n12316) );
  XNOR U12246 ( .A(n11434), .B(n12310), .Z(n12312) );
  XOR U12247 ( .A(n12318), .B(n12319), .Z(n11434) );
  AND U12248 ( .A(n315), .B(n12320), .Z(n12319) );
  XOR U12249 ( .A(n12321), .B(n12318), .Z(n12320) );
  XOR U12250 ( .A(n12322), .B(n12323), .Z(n12310) );
  AND U12251 ( .A(n12324), .B(n12325), .Z(n12323) );
  XOR U12252 ( .A(n12322), .B(n11449), .Z(n12325) );
  XOR U12253 ( .A(n12326), .B(n12327), .Z(n11449) );
  AND U12254 ( .A(n318), .B(n12328), .Z(n12327) );
  XOR U12255 ( .A(n12329), .B(n12326), .Z(n12328) );
  XNOR U12256 ( .A(n11446), .B(n12322), .Z(n12324) );
  XOR U12257 ( .A(n12330), .B(n12331), .Z(n11446) );
  AND U12258 ( .A(n315), .B(n12332), .Z(n12331) );
  XOR U12259 ( .A(n12333), .B(n12330), .Z(n12332) );
  XOR U12260 ( .A(n12334), .B(n12335), .Z(n12322) );
  AND U12261 ( .A(n12336), .B(n12337), .Z(n12335) );
  XOR U12262 ( .A(n12334), .B(n11461), .Z(n12337) );
  XOR U12263 ( .A(n12338), .B(n12339), .Z(n11461) );
  AND U12264 ( .A(n318), .B(n12340), .Z(n12339) );
  XOR U12265 ( .A(n12341), .B(n12338), .Z(n12340) );
  XNOR U12266 ( .A(n11458), .B(n12334), .Z(n12336) );
  XOR U12267 ( .A(n12342), .B(n12343), .Z(n11458) );
  AND U12268 ( .A(n315), .B(n12344), .Z(n12343) );
  XOR U12269 ( .A(n12345), .B(n12342), .Z(n12344) );
  XOR U12270 ( .A(n12346), .B(n12347), .Z(n12334) );
  AND U12271 ( .A(n12348), .B(n12349), .Z(n12347) );
  XOR U12272 ( .A(n12346), .B(n11473), .Z(n12349) );
  XOR U12273 ( .A(n12350), .B(n12351), .Z(n11473) );
  AND U12274 ( .A(n318), .B(n12352), .Z(n12351) );
  XOR U12275 ( .A(n12353), .B(n12350), .Z(n12352) );
  XNOR U12276 ( .A(n11470), .B(n12346), .Z(n12348) );
  XOR U12277 ( .A(n12354), .B(n12355), .Z(n11470) );
  AND U12278 ( .A(n315), .B(n12356), .Z(n12355) );
  XOR U12279 ( .A(n12357), .B(n12354), .Z(n12356) );
  XOR U12280 ( .A(n12358), .B(n12359), .Z(n12346) );
  AND U12281 ( .A(n12360), .B(n12361), .Z(n12359) );
  XOR U12282 ( .A(n12358), .B(n11485), .Z(n12361) );
  XOR U12283 ( .A(n12362), .B(n12363), .Z(n11485) );
  AND U12284 ( .A(n318), .B(n12364), .Z(n12363) );
  XOR U12285 ( .A(n12365), .B(n12362), .Z(n12364) );
  XNOR U12286 ( .A(n11482), .B(n12358), .Z(n12360) );
  XOR U12287 ( .A(n12366), .B(n12367), .Z(n11482) );
  AND U12288 ( .A(n315), .B(n12368), .Z(n12367) );
  XOR U12289 ( .A(n12369), .B(n12366), .Z(n12368) );
  XOR U12290 ( .A(n12370), .B(n12371), .Z(n12358) );
  AND U12291 ( .A(n12372), .B(n12373), .Z(n12371) );
  XOR U12292 ( .A(n12370), .B(n11497), .Z(n12373) );
  XOR U12293 ( .A(n12374), .B(n12375), .Z(n11497) );
  AND U12294 ( .A(n318), .B(n12376), .Z(n12375) );
  XOR U12295 ( .A(n12377), .B(n12374), .Z(n12376) );
  XNOR U12296 ( .A(n11494), .B(n12370), .Z(n12372) );
  XOR U12297 ( .A(n12378), .B(n12379), .Z(n11494) );
  AND U12298 ( .A(n315), .B(n12380), .Z(n12379) );
  XOR U12299 ( .A(n12381), .B(n12378), .Z(n12380) );
  XOR U12300 ( .A(n12382), .B(n12383), .Z(n12370) );
  AND U12301 ( .A(n12384), .B(n12385), .Z(n12383) );
  XOR U12302 ( .A(n12382), .B(n11509), .Z(n12385) );
  XOR U12303 ( .A(n12386), .B(n12387), .Z(n11509) );
  AND U12304 ( .A(n318), .B(n12388), .Z(n12387) );
  XOR U12305 ( .A(n12389), .B(n12386), .Z(n12388) );
  XNOR U12306 ( .A(n11506), .B(n12382), .Z(n12384) );
  XOR U12307 ( .A(n12390), .B(n12391), .Z(n11506) );
  AND U12308 ( .A(n315), .B(n12392), .Z(n12391) );
  XOR U12309 ( .A(n12393), .B(n12390), .Z(n12392) );
  XOR U12310 ( .A(n12394), .B(n12395), .Z(n12382) );
  AND U12311 ( .A(n12396), .B(n12397), .Z(n12395) );
  XOR U12312 ( .A(n12394), .B(n11521), .Z(n12397) );
  XOR U12313 ( .A(n12398), .B(n12399), .Z(n11521) );
  AND U12314 ( .A(n318), .B(n12400), .Z(n12399) );
  XOR U12315 ( .A(n12401), .B(n12398), .Z(n12400) );
  XNOR U12316 ( .A(n11518), .B(n12394), .Z(n12396) );
  XOR U12317 ( .A(n12402), .B(n12403), .Z(n11518) );
  AND U12318 ( .A(n315), .B(n12404), .Z(n12403) );
  XOR U12319 ( .A(n12405), .B(n12402), .Z(n12404) );
  XOR U12320 ( .A(n12406), .B(n12407), .Z(n12394) );
  AND U12321 ( .A(n12408), .B(n12409), .Z(n12407) );
  XOR U12322 ( .A(n12406), .B(n11533), .Z(n12409) );
  XOR U12323 ( .A(n12410), .B(n12411), .Z(n11533) );
  AND U12324 ( .A(n318), .B(n12412), .Z(n12411) );
  XOR U12325 ( .A(n12413), .B(n12410), .Z(n12412) );
  XNOR U12326 ( .A(n11530), .B(n12406), .Z(n12408) );
  XOR U12327 ( .A(n12414), .B(n12415), .Z(n11530) );
  AND U12328 ( .A(n315), .B(n12416), .Z(n12415) );
  XOR U12329 ( .A(n12417), .B(n12414), .Z(n12416) );
  XOR U12330 ( .A(n12418), .B(n12419), .Z(n12406) );
  AND U12331 ( .A(n12420), .B(n12421), .Z(n12419) );
  XOR U12332 ( .A(n11545), .B(n12418), .Z(n12421) );
  XOR U12333 ( .A(n12422), .B(n12423), .Z(n11545) );
  AND U12334 ( .A(n318), .B(n12424), .Z(n12423) );
  XOR U12335 ( .A(n12422), .B(n12425), .Z(n12424) );
  XNOR U12336 ( .A(n12418), .B(n11542), .Z(n12420) );
  XOR U12337 ( .A(n12426), .B(n12427), .Z(n11542) );
  AND U12338 ( .A(n315), .B(n12428), .Z(n12427) );
  XOR U12339 ( .A(n12426), .B(n12429), .Z(n12428) );
  XOR U12340 ( .A(n12430), .B(n12431), .Z(n12418) );
  AND U12341 ( .A(n12432), .B(n12433), .Z(n12431) );
  XNOR U12342 ( .A(n12434), .B(n11558), .Z(n12433) );
  XOR U12343 ( .A(n12435), .B(n12436), .Z(n11558) );
  AND U12344 ( .A(n318), .B(n12437), .Z(n12436) );
  XOR U12345 ( .A(n12438), .B(n12435), .Z(n12437) );
  XNOR U12346 ( .A(n11555), .B(n12430), .Z(n12432) );
  XOR U12347 ( .A(n12439), .B(n12440), .Z(n11555) );
  AND U12348 ( .A(n315), .B(n12441), .Z(n12440) );
  XOR U12349 ( .A(n12442), .B(n12439), .Z(n12441) );
  IV U12350 ( .A(n12434), .Z(n12430) );
  AND U12351 ( .A(n12262), .B(n12265), .Z(n12434) );
  XNOR U12352 ( .A(n12443), .B(n12444), .Z(n12265) );
  AND U12353 ( .A(n318), .B(n12445), .Z(n12444) );
  XNOR U12354 ( .A(n12446), .B(n12443), .Z(n12445) );
  XOR U12355 ( .A(n12447), .B(n12448), .Z(n318) );
  AND U12356 ( .A(n12449), .B(n12450), .Z(n12448) );
  XNOR U12357 ( .A(n12270), .B(n12447), .Z(n12450) );
  AND U12358 ( .A(p_input[383]), .B(p_input[367]), .Z(n12270) );
  XOR U12359 ( .A(n12447), .B(n12271), .Z(n12449) );
  AND U12360 ( .A(p_input[351]), .B(p_input[335]), .Z(n12271) );
  XOR U12361 ( .A(n12451), .B(n12452), .Z(n12447) );
  AND U12362 ( .A(n12453), .B(n12454), .Z(n12452) );
  XOR U12363 ( .A(n12451), .B(n12281), .Z(n12454) );
  XNOR U12364 ( .A(p_input[366]), .B(n12455), .Z(n12281) );
  AND U12365 ( .A(n482), .B(n12456), .Z(n12455) );
  XOR U12366 ( .A(p_input[382]), .B(p_input[366]), .Z(n12456) );
  XNOR U12367 ( .A(n12278), .B(n12451), .Z(n12453) );
  XOR U12368 ( .A(n12457), .B(n12458), .Z(n12278) );
  AND U12369 ( .A(n480), .B(n12459), .Z(n12458) );
  XOR U12370 ( .A(p_input[350]), .B(p_input[334]), .Z(n12459) );
  XOR U12371 ( .A(n12460), .B(n12461), .Z(n12451) );
  AND U12372 ( .A(n12462), .B(n12463), .Z(n12461) );
  XOR U12373 ( .A(n12460), .B(n12293), .Z(n12463) );
  XNOR U12374 ( .A(p_input[365]), .B(n12464), .Z(n12293) );
  AND U12375 ( .A(n482), .B(n12465), .Z(n12464) );
  XOR U12376 ( .A(p_input[381]), .B(p_input[365]), .Z(n12465) );
  XNOR U12377 ( .A(n12290), .B(n12460), .Z(n12462) );
  XOR U12378 ( .A(n12466), .B(n12467), .Z(n12290) );
  AND U12379 ( .A(n480), .B(n12468), .Z(n12467) );
  XOR U12380 ( .A(p_input[349]), .B(p_input[333]), .Z(n12468) );
  XOR U12381 ( .A(n12469), .B(n12470), .Z(n12460) );
  AND U12382 ( .A(n12471), .B(n12472), .Z(n12470) );
  XOR U12383 ( .A(n12469), .B(n12305), .Z(n12472) );
  XNOR U12384 ( .A(p_input[364]), .B(n12473), .Z(n12305) );
  AND U12385 ( .A(n482), .B(n12474), .Z(n12473) );
  XOR U12386 ( .A(p_input[380]), .B(p_input[364]), .Z(n12474) );
  XNOR U12387 ( .A(n12302), .B(n12469), .Z(n12471) );
  XOR U12388 ( .A(n12475), .B(n12476), .Z(n12302) );
  AND U12389 ( .A(n480), .B(n12477), .Z(n12476) );
  XOR U12390 ( .A(p_input[348]), .B(p_input[332]), .Z(n12477) );
  XOR U12391 ( .A(n12478), .B(n12479), .Z(n12469) );
  AND U12392 ( .A(n12480), .B(n12481), .Z(n12479) );
  XOR U12393 ( .A(n12478), .B(n12317), .Z(n12481) );
  XNOR U12394 ( .A(p_input[363]), .B(n12482), .Z(n12317) );
  AND U12395 ( .A(n482), .B(n12483), .Z(n12482) );
  XOR U12396 ( .A(p_input[379]), .B(p_input[363]), .Z(n12483) );
  XNOR U12397 ( .A(n12314), .B(n12478), .Z(n12480) );
  XOR U12398 ( .A(n12484), .B(n12485), .Z(n12314) );
  AND U12399 ( .A(n480), .B(n12486), .Z(n12485) );
  XOR U12400 ( .A(p_input[347]), .B(p_input[331]), .Z(n12486) );
  XOR U12401 ( .A(n12487), .B(n12488), .Z(n12478) );
  AND U12402 ( .A(n12489), .B(n12490), .Z(n12488) );
  XOR U12403 ( .A(n12487), .B(n12329), .Z(n12490) );
  XNOR U12404 ( .A(p_input[362]), .B(n12491), .Z(n12329) );
  AND U12405 ( .A(n482), .B(n12492), .Z(n12491) );
  XOR U12406 ( .A(p_input[378]), .B(p_input[362]), .Z(n12492) );
  XNOR U12407 ( .A(n12326), .B(n12487), .Z(n12489) );
  XOR U12408 ( .A(n12493), .B(n12494), .Z(n12326) );
  AND U12409 ( .A(n480), .B(n12495), .Z(n12494) );
  XOR U12410 ( .A(p_input[346]), .B(p_input[330]), .Z(n12495) );
  XOR U12411 ( .A(n12496), .B(n12497), .Z(n12487) );
  AND U12412 ( .A(n12498), .B(n12499), .Z(n12497) );
  XOR U12413 ( .A(n12496), .B(n12341), .Z(n12499) );
  XNOR U12414 ( .A(p_input[361]), .B(n12500), .Z(n12341) );
  AND U12415 ( .A(n482), .B(n12501), .Z(n12500) );
  XOR U12416 ( .A(p_input[377]), .B(p_input[361]), .Z(n12501) );
  XNOR U12417 ( .A(n12338), .B(n12496), .Z(n12498) );
  XOR U12418 ( .A(n12502), .B(n12503), .Z(n12338) );
  AND U12419 ( .A(n480), .B(n12504), .Z(n12503) );
  XOR U12420 ( .A(p_input[345]), .B(p_input[329]), .Z(n12504) );
  XOR U12421 ( .A(n12505), .B(n12506), .Z(n12496) );
  AND U12422 ( .A(n12507), .B(n12508), .Z(n12506) );
  XOR U12423 ( .A(n12505), .B(n12353), .Z(n12508) );
  XNOR U12424 ( .A(p_input[360]), .B(n12509), .Z(n12353) );
  AND U12425 ( .A(n482), .B(n12510), .Z(n12509) );
  XOR U12426 ( .A(p_input[376]), .B(p_input[360]), .Z(n12510) );
  XNOR U12427 ( .A(n12350), .B(n12505), .Z(n12507) );
  XOR U12428 ( .A(n12511), .B(n12512), .Z(n12350) );
  AND U12429 ( .A(n480), .B(n12513), .Z(n12512) );
  XOR U12430 ( .A(p_input[344]), .B(p_input[328]), .Z(n12513) );
  XOR U12431 ( .A(n12514), .B(n12515), .Z(n12505) );
  AND U12432 ( .A(n12516), .B(n12517), .Z(n12515) );
  XOR U12433 ( .A(n12514), .B(n12365), .Z(n12517) );
  XNOR U12434 ( .A(p_input[359]), .B(n12518), .Z(n12365) );
  AND U12435 ( .A(n482), .B(n12519), .Z(n12518) );
  XOR U12436 ( .A(p_input[375]), .B(p_input[359]), .Z(n12519) );
  XNOR U12437 ( .A(n12362), .B(n12514), .Z(n12516) );
  XOR U12438 ( .A(n12520), .B(n12521), .Z(n12362) );
  AND U12439 ( .A(n480), .B(n12522), .Z(n12521) );
  XOR U12440 ( .A(p_input[343]), .B(p_input[327]), .Z(n12522) );
  XOR U12441 ( .A(n12523), .B(n12524), .Z(n12514) );
  AND U12442 ( .A(n12525), .B(n12526), .Z(n12524) );
  XOR U12443 ( .A(n12523), .B(n12377), .Z(n12526) );
  XNOR U12444 ( .A(p_input[358]), .B(n12527), .Z(n12377) );
  AND U12445 ( .A(n482), .B(n12528), .Z(n12527) );
  XOR U12446 ( .A(p_input[374]), .B(p_input[358]), .Z(n12528) );
  XNOR U12447 ( .A(n12374), .B(n12523), .Z(n12525) );
  XOR U12448 ( .A(n12529), .B(n12530), .Z(n12374) );
  AND U12449 ( .A(n480), .B(n12531), .Z(n12530) );
  XOR U12450 ( .A(p_input[342]), .B(p_input[326]), .Z(n12531) );
  XOR U12451 ( .A(n12532), .B(n12533), .Z(n12523) );
  AND U12452 ( .A(n12534), .B(n12535), .Z(n12533) );
  XOR U12453 ( .A(n12532), .B(n12389), .Z(n12535) );
  XNOR U12454 ( .A(p_input[357]), .B(n12536), .Z(n12389) );
  AND U12455 ( .A(n482), .B(n12537), .Z(n12536) );
  XOR U12456 ( .A(p_input[373]), .B(p_input[357]), .Z(n12537) );
  XNOR U12457 ( .A(n12386), .B(n12532), .Z(n12534) );
  XOR U12458 ( .A(n12538), .B(n12539), .Z(n12386) );
  AND U12459 ( .A(n480), .B(n12540), .Z(n12539) );
  XOR U12460 ( .A(p_input[341]), .B(p_input[325]), .Z(n12540) );
  XOR U12461 ( .A(n12541), .B(n12542), .Z(n12532) );
  AND U12462 ( .A(n12543), .B(n12544), .Z(n12542) );
  XOR U12463 ( .A(n12541), .B(n12401), .Z(n12544) );
  XNOR U12464 ( .A(p_input[356]), .B(n12545), .Z(n12401) );
  AND U12465 ( .A(n482), .B(n12546), .Z(n12545) );
  XOR U12466 ( .A(p_input[372]), .B(p_input[356]), .Z(n12546) );
  XNOR U12467 ( .A(n12398), .B(n12541), .Z(n12543) );
  XOR U12468 ( .A(n12547), .B(n12548), .Z(n12398) );
  AND U12469 ( .A(n480), .B(n12549), .Z(n12548) );
  XOR U12470 ( .A(p_input[340]), .B(p_input[324]), .Z(n12549) );
  XOR U12471 ( .A(n12550), .B(n12551), .Z(n12541) );
  AND U12472 ( .A(n12552), .B(n12553), .Z(n12551) );
  XOR U12473 ( .A(n12550), .B(n12413), .Z(n12553) );
  XNOR U12474 ( .A(p_input[355]), .B(n12554), .Z(n12413) );
  AND U12475 ( .A(n482), .B(n12555), .Z(n12554) );
  XOR U12476 ( .A(p_input[371]), .B(p_input[355]), .Z(n12555) );
  XNOR U12477 ( .A(n12410), .B(n12550), .Z(n12552) );
  XOR U12478 ( .A(n12556), .B(n12557), .Z(n12410) );
  AND U12479 ( .A(n480), .B(n12558), .Z(n12557) );
  XOR U12480 ( .A(p_input[339]), .B(p_input[323]), .Z(n12558) );
  XOR U12481 ( .A(n12559), .B(n12560), .Z(n12550) );
  AND U12482 ( .A(n12561), .B(n12562), .Z(n12560) );
  XOR U12483 ( .A(n12425), .B(n12559), .Z(n12562) );
  XNOR U12484 ( .A(p_input[354]), .B(n12563), .Z(n12425) );
  AND U12485 ( .A(n482), .B(n12564), .Z(n12563) );
  XOR U12486 ( .A(p_input[370]), .B(p_input[354]), .Z(n12564) );
  XNOR U12487 ( .A(n12559), .B(n12422), .Z(n12561) );
  XOR U12488 ( .A(n12565), .B(n12566), .Z(n12422) );
  AND U12489 ( .A(n480), .B(n12567), .Z(n12566) );
  XOR U12490 ( .A(p_input[338]), .B(p_input[322]), .Z(n12567) );
  XOR U12491 ( .A(n12568), .B(n12569), .Z(n12559) );
  AND U12492 ( .A(n12570), .B(n12571), .Z(n12569) );
  XNOR U12493 ( .A(n12572), .B(n12438), .Z(n12571) );
  XNOR U12494 ( .A(p_input[353]), .B(n12573), .Z(n12438) );
  AND U12495 ( .A(n482), .B(n12574), .Z(n12573) );
  XNOR U12496 ( .A(p_input[369]), .B(n12575), .Z(n12574) );
  IV U12497 ( .A(p_input[353]), .Z(n12575) );
  XNOR U12498 ( .A(n12435), .B(n12568), .Z(n12570) );
  XNOR U12499 ( .A(p_input[321]), .B(n12576), .Z(n12435) );
  AND U12500 ( .A(n480), .B(n12577), .Z(n12576) );
  XOR U12501 ( .A(p_input[337]), .B(p_input[321]), .Z(n12577) );
  IV U12502 ( .A(n12572), .Z(n12568) );
  AND U12503 ( .A(n12443), .B(n12446), .Z(n12572) );
  XOR U12504 ( .A(p_input[352]), .B(n12578), .Z(n12446) );
  AND U12505 ( .A(n482), .B(n12579), .Z(n12578) );
  XOR U12506 ( .A(p_input[368]), .B(p_input[352]), .Z(n12579) );
  XOR U12507 ( .A(n12580), .B(n12581), .Z(n482) );
  AND U12508 ( .A(n12582), .B(n12583), .Z(n12581) );
  XNOR U12509 ( .A(p_input[383]), .B(n12580), .Z(n12583) );
  XOR U12510 ( .A(n12580), .B(p_input[367]), .Z(n12582) );
  XOR U12511 ( .A(n12584), .B(n12585), .Z(n12580) );
  AND U12512 ( .A(n12586), .B(n12587), .Z(n12585) );
  XNOR U12513 ( .A(p_input[382]), .B(n12584), .Z(n12587) );
  XOR U12514 ( .A(n12584), .B(p_input[366]), .Z(n12586) );
  XOR U12515 ( .A(n12588), .B(n12589), .Z(n12584) );
  AND U12516 ( .A(n12590), .B(n12591), .Z(n12589) );
  XNOR U12517 ( .A(p_input[381]), .B(n12588), .Z(n12591) );
  XOR U12518 ( .A(n12588), .B(p_input[365]), .Z(n12590) );
  XOR U12519 ( .A(n12592), .B(n12593), .Z(n12588) );
  AND U12520 ( .A(n12594), .B(n12595), .Z(n12593) );
  XNOR U12521 ( .A(p_input[380]), .B(n12592), .Z(n12595) );
  XOR U12522 ( .A(n12592), .B(p_input[364]), .Z(n12594) );
  XOR U12523 ( .A(n12596), .B(n12597), .Z(n12592) );
  AND U12524 ( .A(n12598), .B(n12599), .Z(n12597) );
  XNOR U12525 ( .A(p_input[379]), .B(n12596), .Z(n12599) );
  XOR U12526 ( .A(n12596), .B(p_input[363]), .Z(n12598) );
  XOR U12527 ( .A(n12600), .B(n12601), .Z(n12596) );
  AND U12528 ( .A(n12602), .B(n12603), .Z(n12601) );
  XNOR U12529 ( .A(p_input[378]), .B(n12600), .Z(n12603) );
  XOR U12530 ( .A(n12600), .B(p_input[362]), .Z(n12602) );
  XOR U12531 ( .A(n12604), .B(n12605), .Z(n12600) );
  AND U12532 ( .A(n12606), .B(n12607), .Z(n12605) );
  XNOR U12533 ( .A(p_input[377]), .B(n12604), .Z(n12607) );
  XOR U12534 ( .A(n12604), .B(p_input[361]), .Z(n12606) );
  XOR U12535 ( .A(n12608), .B(n12609), .Z(n12604) );
  AND U12536 ( .A(n12610), .B(n12611), .Z(n12609) );
  XNOR U12537 ( .A(p_input[376]), .B(n12608), .Z(n12611) );
  XOR U12538 ( .A(n12608), .B(p_input[360]), .Z(n12610) );
  XOR U12539 ( .A(n12612), .B(n12613), .Z(n12608) );
  AND U12540 ( .A(n12614), .B(n12615), .Z(n12613) );
  XNOR U12541 ( .A(p_input[375]), .B(n12612), .Z(n12615) );
  XOR U12542 ( .A(n12612), .B(p_input[359]), .Z(n12614) );
  XOR U12543 ( .A(n12616), .B(n12617), .Z(n12612) );
  AND U12544 ( .A(n12618), .B(n12619), .Z(n12617) );
  XNOR U12545 ( .A(p_input[374]), .B(n12616), .Z(n12619) );
  XOR U12546 ( .A(n12616), .B(p_input[358]), .Z(n12618) );
  XOR U12547 ( .A(n12620), .B(n12621), .Z(n12616) );
  AND U12548 ( .A(n12622), .B(n12623), .Z(n12621) );
  XNOR U12549 ( .A(p_input[373]), .B(n12620), .Z(n12623) );
  XOR U12550 ( .A(n12620), .B(p_input[357]), .Z(n12622) );
  XOR U12551 ( .A(n12624), .B(n12625), .Z(n12620) );
  AND U12552 ( .A(n12626), .B(n12627), .Z(n12625) );
  XNOR U12553 ( .A(p_input[372]), .B(n12624), .Z(n12627) );
  XOR U12554 ( .A(n12624), .B(p_input[356]), .Z(n12626) );
  XOR U12555 ( .A(n12628), .B(n12629), .Z(n12624) );
  AND U12556 ( .A(n12630), .B(n12631), .Z(n12629) );
  XNOR U12557 ( .A(p_input[371]), .B(n12628), .Z(n12631) );
  XOR U12558 ( .A(n12628), .B(p_input[355]), .Z(n12630) );
  XOR U12559 ( .A(n12632), .B(n12633), .Z(n12628) );
  AND U12560 ( .A(n12634), .B(n12635), .Z(n12633) );
  XNOR U12561 ( .A(p_input[370]), .B(n12632), .Z(n12635) );
  XOR U12562 ( .A(n12632), .B(p_input[354]), .Z(n12634) );
  XNOR U12563 ( .A(n12636), .B(n12637), .Z(n12632) );
  AND U12564 ( .A(n12638), .B(n12639), .Z(n12637) );
  XOR U12565 ( .A(p_input[369]), .B(n12636), .Z(n12639) );
  XNOR U12566 ( .A(p_input[353]), .B(n12636), .Z(n12638) );
  AND U12567 ( .A(p_input[368]), .B(n12640), .Z(n12636) );
  IV U12568 ( .A(p_input[352]), .Z(n12640) );
  XNOR U12569 ( .A(p_input[320]), .B(n12641), .Z(n12443) );
  AND U12570 ( .A(n480), .B(n12642), .Z(n12641) );
  XOR U12571 ( .A(p_input[336]), .B(p_input[320]), .Z(n12642) );
  XOR U12572 ( .A(n12643), .B(n12644), .Z(n480) );
  AND U12573 ( .A(n12645), .B(n12646), .Z(n12644) );
  XNOR U12574 ( .A(p_input[351]), .B(n12643), .Z(n12646) );
  XOR U12575 ( .A(n12643), .B(p_input[335]), .Z(n12645) );
  XOR U12576 ( .A(n12647), .B(n12648), .Z(n12643) );
  AND U12577 ( .A(n12649), .B(n12650), .Z(n12648) );
  XNOR U12578 ( .A(p_input[350]), .B(n12647), .Z(n12650) );
  XNOR U12579 ( .A(n12647), .B(n12457), .Z(n12649) );
  IV U12580 ( .A(p_input[334]), .Z(n12457) );
  XOR U12581 ( .A(n12651), .B(n12652), .Z(n12647) );
  AND U12582 ( .A(n12653), .B(n12654), .Z(n12652) );
  XNOR U12583 ( .A(p_input[349]), .B(n12651), .Z(n12654) );
  XNOR U12584 ( .A(n12651), .B(n12466), .Z(n12653) );
  IV U12585 ( .A(p_input[333]), .Z(n12466) );
  XOR U12586 ( .A(n12655), .B(n12656), .Z(n12651) );
  AND U12587 ( .A(n12657), .B(n12658), .Z(n12656) );
  XNOR U12588 ( .A(p_input[348]), .B(n12655), .Z(n12658) );
  XNOR U12589 ( .A(n12655), .B(n12475), .Z(n12657) );
  IV U12590 ( .A(p_input[332]), .Z(n12475) );
  XOR U12591 ( .A(n12659), .B(n12660), .Z(n12655) );
  AND U12592 ( .A(n12661), .B(n12662), .Z(n12660) );
  XNOR U12593 ( .A(p_input[347]), .B(n12659), .Z(n12662) );
  XNOR U12594 ( .A(n12659), .B(n12484), .Z(n12661) );
  IV U12595 ( .A(p_input[331]), .Z(n12484) );
  XOR U12596 ( .A(n12663), .B(n12664), .Z(n12659) );
  AND U12597 ( .A(n12665), .B(n12666), .Z(n12664) );
  XNOR U12598 ( .A(p_input[346]), .B(n12663), .Z(n12666) );
  XNOR U12599 ( .A(n12663), .B(n12493), .Z(n12665) );
  IV U12600 ( .A(p_input[330]), .Z(n12493) );
  XOR U12601 ( .A(n12667), .B(n12668), .Z(n12663) );
  AND U12602 ( .A(n12669), .B(n12670), .Z(n12668) );
  XNOR U12603 ( .A(p_input[345]), .B(n12667), .Z(n12670) );
  XNOR U12604 ( .A(n12667), .B(n12502), .Z(n12669) );
  IV U12605 ( .A(p_input[329]), .Z(n12502) );
  XOR U12606 ( .A(n12671), .B(n12672), .Z(n12667) );
  AND U12607 ( .A(n12673), .B(n12674), .Z(n12672) );
  XNOR U12608 ( .A(p_input[344]), .B(n12671), .Z(n12674) );
  XNOR U12609 ( .A(n12671), .B(n12511), .Z(n12673) );
  IV U12610 ( .A(p_input[328]), .Z(n12511) );
  XOR U12611 ( .A(n12675), .B(n12676), .Z(n12671) );
  AND U12612 ( .A(n12677), .B(n12678), .Z(n12676) );
  XNOR U12613 ( .A(p_input[343]), .B(n12675), .Z(n12678) );
  XNOR U12614 ( .A(n12675), .B(n12520), .Z(n12677) );
  IV U12615 ( .A(p_input[327]), .Z(n12520) );
  XOR U12616 ( .A(n12679), .B(n12680), .Z(n12675) );
  AND U12617 ( .A(n12681), .B(n12682), .Z(n12680) );
  XNOR U12618 ( .A(p_input[342]), .B(n12679), .Z(n12682) );
  XNOR U12619 ( .A(n12679), .B(n12529), .Z(n12681) );
  IV U12620 ( .A(p_input[326]), .Z(n12529) );
  XOR U12621 ( .A(n12683), .B(n12684), .Z(n12679) );
  AND U12622 ( .A(n12685), .B(n12686), .Z(n12684) );
  XNOR U12623 ( .A(p_input[341]), .B(n12683), .Z(n12686) );
  XNOR U12624 ( .A(n12683), .B(n12538), .Z(n12685) );
  IV U12625 ( .A(p_input[325]), .Z(n12538) );
  XOR U12626 ( .A(n12687), .B(n12688), .Z(n12683) );
  AND U12627 ( .A(n12689), .B(n12690), .Z(n12688) );
  XNOR U12628 ( .A(p_input[340]), .B(n12687), .Z(n12690) );
  XNOR U12629 ( .A(n12687), .B(n12547), .Z(n12689) );
  IV U12630 ( .A(p_input[324]), .Z(n12547) );
  XOR U12631 ( .A(n12691), .B(n12692), .Z(n12687) );
  AND U12632 ( .A(n12693), .B(n12694), .Z(n12692) );
  XNOR U12633 ( .A(p_input[339]), .B(n12691), .Z(n12694) );
  XNOR U12634 ( .A(n12691), .B(n12556), .Z(n12693) );
  IV U12635 ( .A(p_input[323]), .Z(n12556) );
  XOR U12636 ( .A(n12695), .B(n12696), .Z(n12691) );
  AND U12637 ( .A(n12697), .B(n12698), .Z(n12696) );
  XNOR U12638 ( .A(p_input[338]), .B(n12695), .Z(n12698) );
  XNOR U12639 ( .A(n12695), .B(n12565), .Z(n12697) );
  IV U12640 ( .A(p_input[322]), .Z(n12565) );
  XNOR U12641 ( .A(n12699), .B(n12700), .Z(n12695) );
  AND U12642 ( .A(n12701), .B(n12702), .Z(n12700) );
  XOR U12643 ( .A(p_input[337]), .B(n12699), .Z(n12702) );
  XNOR U12644 ( .A(p_input[321]), .B(n12699), .Z(n12701) );
  AND U12645 ( .A(p_input[336]), .B(n12703), .Z(n12699) );
  IV U12646 ( .A(p_input[320]), .Z(n12703) );
  XOR U12647 ( .A(n12704), .B(n12705), .Z(n12262) );
  AND U12648 ( .A(n315), .B(n12706), .Z(n12705) );
  XNOR U12649 ( .A(n12707), .B(n12704), .Z(n12706) );
  XOR U12650 ( .A(n12708), .B(n12709), .Z(n315) );
  AND U12651 ( .A(n12710), .B(n12711), .Z(n12709) );
  XNOR U12652 ( .A(n12273), .B(n12708), .Z(n12711) );
  AND U12653 ( .A(p_input[319]), .B(p_input[303]), .Z(n12273) );
  XOR U12654 ( .A(n12708), .B(n12272), .Z(n12710) );
  AND U12655 ( .A(p_input[271]), .B(p_input[287]), .Z(n12272) );
  XOR U12656 ( .A(n12712), .B(n12713), .Z(n12708) );
  AND U12657 ( .A(n12714), .B(n12715), .Z(n12713) );
  XOR U12658 ( .A(n12712), .B(n12285), .Z(n12715) );
  XNOR U12659 ( .A(p_input[302]), .B(n12716), .Z(n12285) );
  AND U12660 ( .A(n486), .B(n12717), .Z(n12716) );
  XOR U12661 ( .A(p_input[318]), .B(p_input[302]), .Z(n12717) );
  XNOR U12662 ( .A(n12282), .B(n12712), .Z(n12714) );
  XOR U12663 ( .A(n12718), .B(n12719), .Z(n12282) );
  AND U12664 ( .A(n483), .B(n12720), .Z(n12719) );
  XOR U12665 ( .A(p_input[286]), .B(p_input[270]), .Z(n12720) );
  XOR U12666 ( .A(n12721), .B(n12722), .Z(n12712) );
  AND U12667 ( .A(n12723), .B(n12724), .Z(n12722) );
  XOR U12668 ( .A(n12721), .B(n12297), .Z(n12724) );
  XNOR U12669 ( .A(p_input[301]), .B(n12725), .Z(n12297) );
  AND U12670 ( .A(n486), .B(n12726), .Z(n12725) );
  XOR U12671 ( .A(p_input[317]), .B(p_input[301]), .Z(n12726) );
  XNOR U12672 ( .A(n12294), .B(n12721), .Z(n12723) );
  XOR U12673 ( .A(n12727), .B(n12728), .Z(n12294) );
  AND U12674 ( .A(n483), .B(n12729), .Z(n12728) );
  XOR U12675 ( .A(p_input[285]), .B(p_input[269]), .Z(n12729) );
  XOR U12676 ( .A(n12730), .B(n12731), .Z(n12721) );
  AND U12677 ( .A(n12732), .B(n12733), .Z(n12731) );
  XOR U12678 ( .A(n12730), .B(n12309), .Z(n12733) );
  XNOR U12679 ( .A(p_input[300]), .B(n12734), .Z(n12309) );
  AND U12680 ( .A(n486), .B(n12735), .Z(n12734) );
  XOR U12681 ( .A(p_input[316]), .B(p_input[300]), .Z(n12735) );
  XNOR U12682 ( .A(n12306), .B(n12730), .Z(n12732) );
  XOR U12683 ( .A(n12736), .B(n12737), .Z(n12306) );
  AND U12684 ( .A(n483), .B(n12738), .Z(n12737) );
  XOR U12685 ( .A(p_input[284]), .B(p_input[268]), .Z(n12738) );
  XOR U12686 ( .A(n12739), .B(n12740), .Z(n12730) );
  AND U12687 ( .A(n12741), .B(n12742), .Z(n12740) );
  XOR U12688 ( .A(n12739), .B(n12321), .Z(n12742) );
  XNOR U12689 ( .A(p_input[299]), .B(n12743), .Z(n12321) );
  AND U12690 ( .A(n486), .B(n12744), .Z(n12743) );
  XOR U12691 ( .A(p_input[315]), .B(p_input[299]), .Z(n12744) );
  XNOR U12692 ( .A(n12318), .B(n12739), .Z(n12741) );
  XOR U12693 ( .A(n12745), .B(n12746), .Z(n12318) );
  AND U12694 ( .A(n483), .B(n12747), .Z(n12746) );
  XOR U12695 ( .A(p_input[283]), .B(p_input[267]), .Z(n12747) );
  XOR U12696 ( .A(n12748), .B(n12749), .Z(n12739) );
  AND U12697 ( .A(n12750), .B(n12751), .Z(n12749) );
  XOR U12698 ( .A(n12748), .B(n12333), .Z(n12751) );
  XNOR U12699 ( .A(p_input[298]), .B(n12752), .Z(n12333) );
  AND U12700 ( .A(n486), .B(n12753), .Z(n12752) );
  XOR U12701 ( .A(p_input[314]), .B(p_input[298]), .Z(n12753) );
  XNOR U12702 ( .A(n12330), .B(n12748), .Z(n12750) );
  XOR U12703 ( .A(n12754), .B(n12755), .Z(n12330) );
  AND U12704 ( .A(n483), .B(n12756), .Z(n12755) );
  XOR U12705 ( .A(p_input[282]), .B(p_input[266]), .Z(n12756) );
  XOR U12706 ( .A(n12757), .B(n12758), .Z(n12748) );
  AND U12707 ( .A(n12759), .B(n12760), .Z(n12758) );
  XOR U12708 ( .A(n12757), .B(n12345), .Z(n12760) );
  XNOR U12709 ( .A(p_input[297]), .B(n12761), .Z(n12345) );
  AND U12710 ( .A(n486), .B(n12762), .Z(n12761) );
  XOR U12711 ( .A(p_input[313]), .B(p_input[297]), .Z(n12762) );
  XNOR U12712 ( .A(n12342), .B(n12757), .Z(n12759) );
  XOR U12713 ( .A(n12763), .B(n12764), .Z(n12342) );
  AND U12714 ( .A(n483), .B(n12765), .Z(n12764) );
  XOR U12715 ( .A(p_input[281]), .B(p_input[265]), .Z(n12765) );
  XOR U12716 ( .A(n12766), .B(n12767), .Z(n12757) );
  AND U12717 ( .A(n12768), .B(n12769), .Z(n12767) );
  XOR U12718 ( .A(n12766), .B(n12357), .Z(n12769) );
  XNOR U12719 ( .A(p_input[296]), .B(n12770), .Z(n12357) );
  AND U12720 ( .A(n486), .B(n12771), .Z(n12770) );
  XOR U12721 ( .A(p_input[312]), .B(p_input[296]), .Z(n12771) );
  XNOR U12722 ( .A(n12354), .B(n12766), .Z(n12768) );
  XOR U12723 ( .A(n12772), .B(n12773), .Z(n12354) );
  AND U12724 ( .A(n483), .B(n12774), .Z(n12773) );
  XOR U12725 ( .A(p_input[280]), .B(p_input[264]), .Z(n12774) );
  XOR U12726 ( .A(n12775), .B(n12776), .Z(n12766) );
  AND U12727 ( .A(n12777), .B(n12778), .Z(n12776) );
  XOR U12728 ( .A(n12775), .B(n12369), .Z(n12778) );
  XNOR U12729 ( .A(p_input[295]), .B(n12779), .Z(n12369) );
  AND U12730 ( .A(n486), .B(n12780), .Z(n12779) );
  XOR U12731 ( .A(p_input[311]), .B(p_input[295]), .Z(n12780) );
  XNOR U12732 ( .A(n12366), .B(n12775), .Z(n12777) );
  XOR U12733 ( .A(n12781), .B(n12782), .Z(n12366) );
  AND U12734 ( .A(n483), .B(n12783), .Z(n12782) );
  XOR U12735 ( .A(p_input[279]), .B(p_input[263]), .Z(n12783) );
  XOR U12736 ( .A(n12784), .B(n12785), .Z(n12775) );
  AND U12737 ( .A(n12786), .B(n12787), .Z(n12785) );
  XOR U12738 ( .A(n12784), .B(n12381), .Z(n12787) );
  XNOR U12739 ( .A(p_input[294]), .B(n12788), .Z(n12381) );
  AND U12740 ( .A(n486), .B(n12789), .Z(n12788) );
  XOR U12741 ( .A(p_input[310]), .B(p_input[294]), .Z(n12789) );
  XNOR U12742 ( .A(n12378), .B(n12784), .Z(n12786) );
  XOR U12743 ( .A(n12790), .B(n12791), .Z(n12378) );
  AND U12744 ( .A(n483), .B(n12792), .Z(n12791) );
  XOR U12745 ( .A(p_input[278]), .B(p_input[262]), .Z(n12792) );
  XOR U12746 ( .A(n12793), .B(n12794), .Z(n12784) );
  AND U12747 ( .A(n12795), .B(n12796), .Z(n12794) );
  XOR U12748 ( .A(n12793), .B(n12393), .Z(n12796) );
  XNOR U12749 ( .A(p_input[293]), .B(n12797), .Z(n12393) );
  AND U12750 ( .A(n486), .B(n12798), .Z(n12797) );
  XOR U12751 ( .A(p_input[309]), .B(p_input[293]), .Z(n12798) );
  XNOR U12752 ( .A(n12390), .B(n12793), .Z(n12795) );
  XOR U12753 ( .A(n12799), .B(n12800), .Z(n12390) );
  AND U12754 ( .A(n483), .B(n12801), .Z(n12800) );
  XOR U12755 ( .A(p_input[277]), .B(p_input[261]), .Z(n12801) );
  XOR U12756 ( .A(n12802), .B(n12803), .Z(n12793) );
  AND U12757 ( .A(n12804), .B(n12805), .Z(n12803) );
  XOR U12758 ( .A(n12802), .B(n12405), .Z(n12805) );
  XNOR U12759 ( .A(p_input[292]), .B(n12806), .Z(n12405) );
  AND U12760 ( .A(n486), .B(n12807), .Z(n12806) );
  XOR U12761 ( .A(p_input[308]), .B(p_input[292]), .Z(n12807) );
  XNOR U12762 ( .A(n12402), .B(n12802), .Z(n12804) );
  XOR U12763 ( .A(n12808), .B(n12809), .Z(n12402) );
  AND U12764 ( .A(n483), .B(n12810), .Z(n12809) );
  XOR U12765 ( .A(p_input[276]), .B(p_input[260]), .Z(n12810) );
  XOR U12766 ( .A(n12811), .B(n12812), .Z(n12802) );
  AND U12767 ( .A(n12813), .B(n12814), .Z(n12812) );
  XOR U12768 ( .A(n12811), .B(n12417), .Z(n12814) );
  XNOR U12769 ( .A(p_input[291]), .B(n12815), .Z(n12417) );
  AND U12770 ( .A(n486), .B(n12816), .Z(n12815) );
  XOR U12771 ( .A(p_input[307]), .B(p_input[291]), .Z(n12816) );
  XNOR U12772 ( .A(n12414), .B(n12811), .Z(n12813) );
  XOR U12773 ( .A(n12817), .B(n12818), .Z(n12414) );
  AND U12774 ( .A(n483), .B(n12819), .Z(n12818) );
  XOR U12775 ( .A(p_input[275]), .B(p_input[259]), .Z(n12819) );
  XOR U12776 ( .A(n12820), .B(n12821), .Z(n12811) );
  AND U12777 ( .A(n12822), .B(n12823), .Z(n12821) );
  XOR U12778 ( .A(n12429), .B(n12820), .Z(n12823) );
  XNOR U12779 ( .A(p_input[290]), .B(n12824), .Z(n12429) );
  AND U12780 ( .A(n486), .B(n12825), .Z(n12824) );
  XOR U12781 ( .A(p_input[306]), .B(p_input[290]), .Z(n12825) );
  XNOR U12782 ( .A(n12820), .B(n12426), .Z(n12822) );
  XOR U12783 ( .A(n12826), .B(n12827), .Z(n12426) );
  AND U12784 ( .A(n483), .B(n12828), .Z(n12827) );
  XOR U12785 ( .A(p_input[274]), .B(p_input[258]), .Z(n12828) );
  XOR U12786 ( .A(n12829), .B(n12830), .Z(n12820) );
  AND U12787 ( .A(n12831), .B(n12832), .Z(n12830) );
  XNOR U12788 ( .A(n12833), .B(n12442), .Z(n12832) );
  XNOR U12789 ( .A(p_input[289]), .B(n12834), .Z(n12442) );
  AND U12790 ( .A(n486), .B(n12835), .Z(n12834) );
  XNOR U12791 ( .A(p_input[305]), .B(n12836), .Z(n12835) );
  IV U12792 ( .A(p_input[289]), .Z(n12836) );
  XNOR U12793 ( .A(n12439), .B(n12829), .Z(n12831) );
  XNOR U12794 ( .A(p_input[257]), .B(n12837), .Z(n12439) );
  AND U12795 ( .A(n483), .B(n12838), .Z(n12837) );
  XOR U12796 ( .A(p_input[273]), .B(p_input[257]), .Z(n12838) );
  IV U12797 ( .A(n12833), .Z(n12829) );
  AND U12798 ( .A(n12704), .B(n12707), .Z(n12833) );
  XOR U12799 ( .A(p_input[288]), .B(n12839), .Z(n12707) );
  AND U12800 ( .A(n486), .B(n12840), .Z(n12839) );
  XOR U12801 ( .A(p_input[304]), .B(p_input[288]), .Z(n12840) );
  XOR U12802 ( .A(n12841), .B(n12842), .Z(n486) );
  AND U12803 ( .A(n12843), .B(n12844), .Z(n12842) );
  XNOR U12804 ( .A(p_input[319]), .B(n12841), .Z(n12844) );
  XOR U12805 ( .A(n12841), .B(p_input[303]), .Z(n12843) );
  XOR U12806 ( .A(n12845), .B(n12846), .Z(n12841) );
  AND U12807 ( .A(n12847), .B(n12848), .Z(n12846) );
  XNOR U12808 ( .A(p_input[318]), .B(n12845), .Z(n12848) );
  XOR U12809 ( .A(n12845), .B(p_input[302]), .Z(n12847) );
  XOR U12810 ( .A(n12849), .B(n12850), .Z(n12845) );
  AND U12811 ( .A(n12851), .B(n12852), .Z(n12850) );
  XNOR U12812 ( .A(p_input[317]), .B(n12849), .Z(n12852) );
  XOR U12813 ( .A(n12849), .B(p_input[301]), .Z(n12851) );
  XOR U12814 ( .A(n12853), .B(n12854), .Z(n12849) );
  AND U12815 ( .A(n12855), .B(n12856), .Z(n12854) );
  XNOR U12816 ( .A(p_input[316]), .B(n12853), .Z(n12856) );
  XOR U12817 ( .A(n12853), .B(p_input[300]), .Z(n12855) );
  XOR U12818 ( .A(n12857), .B(n12858), .Z(n12853) );
  AND U12819 ( .A(n12859), .B(n12860), .Z(n12858) );
  XNOR U12820 ( .A(p_input[315]), .B(n12857), .Z(n12860) );
  XOR U12821 ( .A(n12857), .B(p_input[299]), .Z(n12859) );
  XOR U12822 ( .A(n12861), .B(n12862), .Z(n12857) );
  AND U12823 ( .A(n12863), .B(n12864), .Z(n12862) );
  XNOR U12824 ( .A(p_input[314]), .B(n12861), .Z(n12864) );
  XOR U12825 ( .A(n12861), .B(p_input[298]), .Z(n12863) );
  XOR U12826 ( .A(n12865), .B(n12866), .Z(n12861) );
  AND U12827 ( .A(n12867), .B(n12868), .Z(n12866) );
  XNOR U12828 ( .A(p_input[313]), .B(n12865), .Z(n12868) );
  XOR U12829 ( .A(n12865), .B(p_input[297]), .Z(n12867) );
  XOR U12830 ( .A(n12869), .B(n12870), .Z(n12865) );
  AND U12831 ( .A(n12871), .B(n12872), .Z(n12870) );
  XNOR U12832 ( .A(p_input[312]), .B(n12869), .Z(n12872) );
  XOR U12833 ( .A(n12869), .B(p_input[296]), .Z(n12871) );
  XOR U12834 ( .A(n12873), .B(n12874), .Z(n12869) );
  AND U12835 ( .A(n12875), .B(n12876), .Z(n12874) );
  XNOR U12836 ( .A(p_input[311]), .B(n12873), .Z(n12876) );
  XOR U12837 ( .A(n12873), .B(p_input[295]), .Z(n12875) );
  XOR U12838 ( .A(n12877), .B(n12878), .Z(n12873) );
  AND U12839 ( .A(n12879), .B(n12880), .Z(n12878) );
  XNOR U12840 ( .A(p_input[310]), .B(n12877), .Z(n12880) );
  XOR U12841 ( .A(n12877), .B(p_input[294]), .Z(n12879) );
  XOR U12842 ( .A(n12881), .B(n12882), .Z(n12877) );
  AND U12843 ( .A(n12883), .B(n12884), .Z(n12882) );
  XNOR U12844 ( .A(p_input[309]), .B(n12881), .Z(n12884) );
  XOR U12845 ( .A(n12881), .B(p_input[293]), .Z(n12883) );
  XOR U12846 ( .A(n12885), .B(n12886), .Z(n12881) );
  AND U12847 ( .A(n12887), .B(n12888), .Z(n12886) );
  XNOR U12848 ( .A(p_input[308]), .B(n12885), .Z(n12888) );
  XOR U12849 ( .A(n12885), .B(p_input[292]), .Z(n12887) );
  XOR U12850 ( .A(n12889), .B(n12890), .Z(n12885) );
  AND U12851 ( .A(n12891), .B(n12892), .Z(n12890) );
  XNOR U12852 ( .A(p_input[307]), .B(n12889), .Z(n12892) );
  XOR U12853 ( .A(n12889), .B(p_input[291]), .Z(n12891) );
  XOR U12854 ( .A(n12893), .B(n12894), .Z(n12889) );
  AND U12855 ( .A(n12895), .B(n12896), .Z(n12894) );
  XNOR U12856 ( .A(p_input[306]), .B(n12893), .Z(n12896) );
  XOR U12857 ( .A(n12893), .B(p_input[290]), .Z(n12895) );
  XNOR U12858 ( .A(n12897), .B(n12898), .Z(n12893) );
  AND U12859 ( .A(n12899), .B(n12900), .Z(n12898) );
  XOR U12860 ( .A(p_input[305]), .B(n12897), .Z(n12900) );
  XNOR U12861 ( .A(p_input[289]), .B(n12897), .Z(n12899) );
  AND U12862 ( .A(p_input[304]), .B(n12901), .Z(n12897) );
  IV U12863 ( .A(p_input[288]), .Z(n12901) );
  XNOR U12864 ( .A(p_input[256]), .B(n12902), .Z(n12704) );
  AND U12865 ( .A(n483), .B(n12903), .Z(n12902) );
  XOR U12866 ( .A(p_input[272]), .B(p_input[256]), .Z(n12903) );
  XOR U12867 ( .A(n12904), .B(n12905), .Z(n483) );
  AND U12868 ( .A(n12906), .B(n12907), .Z(n12905) );
  XNOR U12869 ( .A(p_input[287]), .B(n12904), .Z(n12907) );
  XOR U12870 ( .A(n12904), .B(p_input[271]), .Z(n12906) );
  XOR U12871 ( .A(n12908), .B(n12909), .Z(n12904) );
  AND U12872 ( .A(n12910), .B(n12911), .Z(n12909) );
  XNOR U12873 ( .A(p_input[286]), .B(n12908), .Z(n12911) );
  XNOR U12874 ( .A(n12908), .B(n12718), .Z(n12910) );
  IV U12875 ( .A(p_input[270]), .Z(n12718) );
  XOR U12876 ( .A(n12912), .B(n12913), .Z(n12908) );
  AND U12877 ( .A(n12914), .B(n12915), .Z(n12913) );
  XNOR U12878 ( .A(p_input[285]), .B(n12912), .Z(n12915) );
  XNOR U12879 ( .A(n12912), .B(n12727), .Z(n12914) );
  IV U12880 ( .A(p_input[269]), .Z(n12727) );
  XOR U12881 ( .A(n12916), .B(n12917), .Z(n12912) );
  AND U12882 ( .A(n12918), .B(n12919), .Z(n12917) );
  XNOR U12883 ( .A(p_input[284]), .B(n12916), .Z(n12919) );
  XNOR U12884 ( .A(n12916), .B(n12736), .Z(n12918) );
  IV U12885 ( .A(p_input[268]), .Z(n12736) );
  XOR U12886 ( .A(n12920), .B(n12921), .Z(n12916) );
  AND U12887 ( .A(n12922), .B(n12923), .Z(n12921) );
  XNOR U12888 ( .A(p_input[283]), .B(n12920), .Z(n12923) );
  XNOR U12889 ( .A(n12920), .B(n12745), .Z(n12922) );
  IV U12890 ( .A(p_input[267]), .Z(n12745) );
  XOR U12891 ( .A(n12924), .B(n12925), .Z(n12920) );
  AND U12892 ( .A(n12926), .B(n12927), .Z(n12925) );
  XNOR U12893 ( .A(p_input[282]), .B(n12924), .Z(n12927) );
  XNOR U12894 ( .A(n12924), .B(n12754), .Z(n12926) );
  IV U12895 ( .A(p_input[266]), .Z(n12754) );
  XOR U12896 ( .A(n12928), .B(n12929), .Z(n12924) );
  AND U12897 ( .A(n12930), .B(n12931), .Z(n12929) );
  XNOR U12898 ( .A(p_input[281]), .B(n12928), .Z(n12931) );
  XNOR U12899 ( .A(n12928), .B(n12763), .Z(n12930) );
  IV U12900 ( .A(p_input[265]), .Z(n12763) );
  XOR U12901 ( .A(n12932), .B(n12933), .Z(n12928) );
  AND U12902 ( .A(n12934), .B(n12935), .Z(n12933) );
  XNOR U12903 ( .A(p_input[280]), .B(n12932), .Z(n12935) );
  XNOR U12904 ( .A(n12932), .B(n12772), .Z(n12934) );
  IV U12905 ( .A(p_input[264]), .Z(n12772) );
  XOR U12906 ( .A(n12936), .B(n12937), .Z(n12932) );
  AND U12907 ( .A(n12938), .B(n12939), .Z(n12937) );
  XNOR U12908 ( .A(p_input[279]), .B(n12936), .Z(n12939) );
  XNOR U12909 ( .A(n12936), .B(n12781), .Z(n12938) );
  IV U12910 ( .A(p_input[263]), .Z(n12781) );
  XOR U12911 ( .A(n12940), .B(n12941), .Z(n12936) );
  AND U12912 ( .A(n12942), .B(n12943), .Z(n12941) );
  XNOR U12913 ( .A(p_input[278]), .B(n12940), .Z(n12943) );
  XNOR U12914 ( .A(n12940), .B(n12790), .Z(n12942) );
  IV U12915 ( .A(p_input[262]), .Z(n12790) );
  XOR U12916 ( .A(n12944), .B(n12945), .Z(n12940) );
  AND U12917 ( .A(n12946), .B(n12947), .Z(n12945) );
  XNOR U12918 ( .A(p_input[277]), .B(n12944), .Z(n12947) );
  XNOR U12919 ( .A(n12944), .B(n12799), .Z(n12946) );
  IV U12920 ( .A(p_input[261]), .Z(n12799) );
  XOR U12921 ( .A(n12948), .B(n12949), .Z(n12944) );
  AND U12922 ( .A(n12950), .B(n12951), .Z(n12949) );
  XNOR U12923 ( .A(p_input[276]), .B(n12948), .Z(n12951) );
  XNOR U12924 ( .A(n12948), .B(n12808), .Z(n12950) );
  IV U12925 ( .A(p_input[260]), .Z(n12808) );
  XOR U12926 ( .A(n12952), .B(n12953), .Z(n12948) );
  AND U12927 ( .A(n12954), .B(n12955), .Z(n12953) );
  XNOR U12928 ( .A(p_input[275]), .B(n12952), .Z(n12955) );
  XNOR U12929 ( .A(n12952), .B(n12817), .Z(n12954) );
  IV U12930 ( .A(p_input[259]), .Z(n12817) );
  XOR U12931 ( .A(n12956), .B(n12957), .Z(n12952) );
  AND U12932 ( .A(n12958), .B(n12959), .Z(n12957) );
  XNOR U12933 ( .A(p_input[274]), .B(n12956), .Z(n12959) );
  XNOR U12934 ( .A(n12956), .B(n12826), .Z(n12958) );
  IV U12935 ( .A(p_input[258]), .Z(n12826) );
  XNOR U12936 ( .A(n12960), .B(n12961), .Z(n12956) );
  AND U12937 ( .A(n12962), .B(n12963), .Z(n12961) );
  XOR U12938 ( .A(p_input[273]), .B(n12960), .Z(n12963) );
  XNOR U12939 ( .A(p_input[257]), .B(n12960), .Z(n12962) );
  AND U12940 ( .A(p_input[272]), .B(n12964), .Z(n12960) );
  IV U12941 ( .A(p_input[256]), .Z(n12964) );
  XOR U12942 ( .A(n12965), .B(n12966), .Z(n11192) );
  AND U12943 ( .A(n511), .B(n12967), .Z(n12966) );
  XNOR U12944 ( .A(n12968), .B(n12965), .Z(n12967) );
  XOR U12945 ( .A(n12969), .B(n12970), .Z(n511) );
  AND U12946 ( .A(n12971), .B(n12972), .Z(n12970) );
  XNOR U12947 ( .A(n11207), .B(n12969), .Z(n12972) );
  AND U12948 ( .A(n12973), .B(n12974), .Z(n11207) );
  XNOR U12949 ( .A(n12969), .B(n11204), .Z(n12971) );
  IV U12950 ( .A(n12975), .Z(n11204) );
  AND U12951 ( .A(n12976), .B(n12977), .Z(n12975) );
  XOR U12952 ( .A(n12978), .B(n12979), .Z(n12969) );
  AND U12953 ( .A(n12980), .B(n12981), .Z(n12979) );
  XOR U12954 ( .A(n12978), .B(n11219), .Z(n12981) );
  XOR U12955 ( .A(n12982), .B(n12983), .Z(n11219) );
  AND U12956 ( .A(n454), .B(n12984), .Z(n12983) );
  XOR U12957 ( .A(n12985), .B(n12982), .Z(n12984) );
  XNOR U12958 ( .A(n11216), .B(n12978), .Z(n12980) );
  XOR U12959 ( .A(n12986), .B(n12987), .Z(n11216) );
  AND U12960 ( .A(n451), .B(n12988), .Z(n12987) );
  XOR U12961 ( .A(n12989), .B(n12986), .Z(n12988) );
  XOR U12962 ( .A(n12990), .B(n12991), .Z(n12978) );
  AND U12963 ( .A(n12992), .B(n12993), .Z(n12991) );
  XOR U12964 ( .A(n12990), .B(n11231), .Z(n12993) );
  XOR U12965 ( .A(n12994), .B(n12995), .Z(n11231) );
  AND U12966 ( .A(n454), .B(n12996), .Z(n12995) );
  XOR U12967 ( .A(n12997), .B(n12994), .Z(n12996) );
  XNOR U12968 ( .A(n11228), .B(n12990), .Z(n12992) );
  XOR U12969 ( .A(n12998), .B(n12999), .Z(n11228) );
  AND U12970 ( .A(n451), .B(n13000), .Z(n12999) );
  XOR U12971 ( .A(n13001), .B(n12998), .Z(n13000) );
  XOR U12972 ( .A(n13002), .B(n13003), .Z(n12990) );
  AND U12973 ( .A(n13004), .B(n13005), .Z(n13003) );
  XOR U12974 ( .A(n13002), .B(n11243), .Z(n13005) );
  XOR U12975 ( .A(n13006), .B(n13007), .Z(n11243) );
  AND U12976 ( .A(n454), .B(n13008), .Z(n13007) );
  XOR U12977 ( .A(n13009), .B(n13006), .Z(n13008) );
  XNOR U12978 ( .A(n11240), .B(n13002), .Z(n13004) );
  XOR U12979 ( .A(n13010), .B(n13011), .Z(n11240) );
  AND U12980 ( .A(n451), .B(n13012), .Z(n13011) );
  XOR U12981 ( .A(n13013), .B(n13010), .Z(n13012) );
  XOR U12982 ( .A(n13014), .B(n13015), .Z(n13002) );
  AND U12983 ( .A(n13016), .B(n13017), .Z(n13015) );
  XOR U12984 ( .A(n13014), .B(n11255), .Z(n13017) );
  XOR U12985 ( .A(n13018), .B(n13019), .Z(n11255) );
  AND U12986 ( .A(n454), .B(n13020), .Z(n13019) );
  XOR U12987 ( .A(n13021), .B(n13018), .Z(n13020) );
  XNOR U12988 ( .A(n11252), .B(n13014), .Z(n13016) );
  XOR U12989 ( .A(n13022), .B(n13023), .Z(n11252) );
  AND U12990 ( .A(n451), .B(n13024), .Z(n13023) );
  XOR U12991 ( .A(n13025), .B(n13022), .Z(n13024) );
  XOR U12992 ( .A(n13026), .B(n13027), .Z(n13014) );
  AND U12993 ( .A(n13028), .B(n13029), .Z(n13027) );
  XOR U12994 ( .A(n13026), .B(n11267), .Z(n13029) );
  XOR U12995 ( .A(n13030), .B(n13031), .Z(n11267) );
  AND U12996 ( .A(n454), .B(n13032), .Z(n13031) );
  XOR U12997 ( .A(n13033), .B(n13030), .Z(n13032) );
  XNOR U12998 ( .A(n11264), .B(n13026), .Z(n13028) );
  XOR U12999 ( .A(n13034), .B(n13035), .Z(n11264) );
  AND U13000 ( .A(n451), .B(n13036), .Z(n13035) );
  XOR U13001 ( .A(n13037), .B(n13034), .Z(n13036) );
  XOR U13002 ( .A(n13038), .B(n13039), .Z(n13026) );
  AND U13003 ( .A(n13040), .B(n13041), .Z(n13039) );
  XOR U13004 ( .A(n13038), .B(n11279), .Z(n13041) );
  XOR U13005 ( .A(n13042), .B(n13043), .Z(n11279) );
  AND U13006 ( .A(n454), .B(n13044), .Z(n13043) );
  XOR U13007 ( .A(n13045), .B(n13042), .Z(n13044) );
  XNOR U13008 ( .A(n11276), .B(n13038), .Z(n13040) );
  XOR U13009 ( .A(n13046), .B(n13047), .Z(n11276) );
  AND U13010 ( .A(n451), .B(n13048), .Z(n13047) );
  XOR U13011 ( .A(n13049), .B(n13046), .Z(n13048) );
  XOR U13012 ( .A(n13050), .B(n13051), .Z(n13038) );
  AND U13013 ( .A(n13052), .B(n13053), .Z(n13051) );
  XOR U13014 ( .A(n13050), .B(n11291), .Z(n13053) );
  XOR U13015 ( .A(n13054), .B(n13055), .Z(n11291) );
  AND U13016 ( .A(n454), .B(n13056), .Z(n13055) );
  XOR U13017 ( .A(n13057), .B(n13054), .Z(n13056) );
  XNOR U13018 ( .A(n11288), .B(n13050), .Z(n13052) );
  XOR U13019 ( .A(n13058), .B(n13059), .Z(n11288) );
  AND U13020 ( .A(n451), .B(n13060), .Z(n13059) );
  XOR U13021 ( .A(n13061), .B(n13058), .Z(n13060) );
  XOR U13022 ( .A(n13062), .B(n13063), .Z(n13050) );
  AND U13023 ( .A(n13064), .B(n13065), .Z(n13063) );
  XOR U13024 ( .A(n13062), .B(n11303), .Z(n13065) );
  XOR U13025 ( .A(n13066), .B(n13067), .Z(n11303) );
  AND U13026 ( .A(n454), .B(n13068), .Z(n13067) );
  XOR U13027 ( .A(n13069), .B(n13066), .Z(n13068) );
  XNOR U13028 ( .A(n11300), .B(n13062), .Z(n13064) );
  XOR U13029 ( .A(n13070), .B(n13071), .Z(n11300) );
  AND U13030 ( .A(n451), .B(n13072), .Z(n13071) );
  XOR U13031 ( .A(n13073), .B(n13070), .Z(n13072) );
  XOR U13032 ( .A(n13074), .B(n13075), .Z(n13062) );
  AND U13033 ( .A(n13076), .B(n13077), .Z(n13075) );
  XOR U13034 ( .A(n13074), .B(n11315), .Z(n13077) );
  XOR U13035 ( .A(n13078), .B(n13079), .Z(n11315) );
  AND U13036 ( .A(n454), .B(n13080), .Z(n13079) );
  XOR U13037 ( .A(n13081), .B(n13078), .Z(n13080) );
  XNOR U13038 ( .A(n11312), .B(n13074), .Z(n13076) );
  XOR U13039 ( .A(n13082), .B(n13083), .Z(n11312) );
  AND U13040 ( .A(n451), .B(n13084), .Z(n13083) );
  XOR U13041 ( .A(n13085), .B(n13082), .Z(n13084) );
  XOR U13042 ( .A(n13086), .B(n13087), .Z(n13074) );
  AND U13043 ( .A(n13088), .B(n13089), .Z(n13087) );
  XOR U13044 ( .A(n13086), .B(n11327), .Z(n13089) );
  XOR U13045 ( .A(n13090), .B(n13091), .Z(n11327) );
  AND U13046 ( .A(n454), .B(n13092), .Z(n13091) );
  XOR U13047 ( .A(n13093), .B(n13090), .Z(n13092) );
  XNOR U13048 ( .A(n11324), .B(n13086), .Z(n13088) );
  XOR U13049 ( .A(n13094), .B(n13095), .Z(n11324) );
  AND U13050 ( .A(n451), .B(n13096), .Z(n13095) );
  XOR U13051 ( .A(n13097), .B(n13094), .Z(n13096) );
  XOR U13052 ( .A(n13098), .B(n13099), .Z(n13086) );
  AND U13053 ( .A(n13100), .B(n13101), .Z(n13099) );
  XOR U13054 ( .A(n13098), .B(n11339), .Z(n13101) );
  XOR U13055 ( .A(n13102), .B(n13103), .Z(n11339) );
  AND U13056 ( .A(n454), .B(n13104), .Z(n13103) );
  XOR U13057 ( .A(n13105), .B(n13102), .Z(n13104) );
  XNOR U13058 ( .A(n11336), .B(n13098), .Z(n13100) );
  XOR U13059 ( .A(n13106), .B(n13107), .Z(n11336) );
  AND U13060 ( .A(n451), .B(n13108), .Z(n13107) );
  XOR U13061 ( .A(n13109), .B(n13106), .Z(n13108) );
  XOR U13062 ( .A(n13110), .B(n13111), .Z(n13098) );
  AND U13063 ( .A(n13112), .B(n13113), .Z(n13111) );
  XOR U13064 ( .A(n13110), .B(n11351), .Z(n13113) );
  XOR U13065 ( .A(n13114), .B(n13115), .Z(n11351) );
  AND U13066 ( .A(n454), .B(n13116), .Z(n13115) );
  XOR U13067 ( .A(n13117), .B(n13114), .Z(n13116) );
  XNOR U13068 ( .A(n11348), .B(n13110), .Z(n13112) );
  XOR U13069 ( .A(n13118), .B(n13119), .Z(n11348) );
  AND U13070 ( .A(n451), .B(n13120), .Z(n13119) );
  XOR U13071 ( .A(n13121), .B(n13118), .Z(n13120) );
  XOR U13072 ( .A(n13122), .B(n13123), .Z(n13110) );
  AND U13073 ( .A(n13124), .B(n13125), .Z(n13123) );
  XOR U13074 ( .A(n11363), .B(n13122), .Z(n13125) );
  XOR U13075 ( .A(n13126), .B(n13127), .Z(n11363) );
  AND U13076 ( .A(n454), .B(n13128), .Z(n13127) );
  XOR U13077 ( .A(n13126), .B(n13129), .Z(n13128) );
  XNOR U13078 ( .A(n13122), .B(n11360), .Z(n13124) );
  XOR U13079 ( .A(n13130), .B(n13131), .Z(n11360) );
  AND U13080 ( .A(n451), .B(n13132), .Z(n13131) );
  XOR U13081 ( .A(n13130), .B(n13133), .Z(n13132) );
  XOR U13082 ( .A(n13134), .B(n13135), .Z(n13122) );
  AND U13083 ( .A(n13136), .B(n13137), .Z(n13135) );
  XNOR U13084 ( .A(n13138), .B(n11376), .Z(n13137) );
  XOR U13085 ( .A(n13139), .B(n13140), .Z(n11376) );
  AND U13086 ( .A(n454), .B(n13141), .Z(n13140) );
  XOR U13087 ( .A(n13142), .B(n13139), .Z(n13141) );
  XNOR U13088 ( .A(n11373), .B(n13134), .Z(n13136) );
  XOR U13089 ( .A(n13143), .B(n13144), .Z(n11373) );
  AND U13090 ( .A(n451), .B(n13145), .Z(n13144) );
  XOR U13091 ( .A(n13146), .B(n13143), .Z(n13145) );
  IV U13092 ( .A(n13138), .Z(n13134) );
  AND U13093 ( .A(n12965), .B(n12968), .Z(n13138) );
  XNOR U13094 ( .A(n13147), .B(n13148), .Z(n12968) );
  AND U13095 ( .A(n454), .B(n13149), .Z(n13148) );
  XNOR U13096 ( .A(n13150), .B(n13147), .Z(n13149) );
  XOR U13097 ( .A(n13151), .B(n13152), .Z(n454) );
  AND U13098 ( .A(n13153), .B(n13154), .Z(n13152) );
  XNOR U13099 ( .A(n12973), .B(n13151), .Z(n13154) );
  AND U13100 ( .A(n13155), .B(n13156), .Z(n12973) );
  XOR U13101 ( .A(n13151), .B(n12974), .Z(n13153) );
  AND U13102 ( .A(n13157), .B(n13158), .Z(n12974) );
  XOR U13103 ( .A(n13159), .B(n13160), .Z(n13151) );
  AND U13104 ( .A(n13161), .B(n13162), .Z(n13160) );
  XOR U13105 ( .A(n13159), .B(n12985), .Z(n13162) );
  XOR U13106 ( .A(n13163), .B(n13164), .Z(n12985) );
  AND U13107 ( .A(n326), .B(n13165), .Z(n13164) );
  XOR U13108 ( .A(n13166), .B(n13163), .Z(n13165) );
  XNOR U13109 ( .A(n12982), .B(n13159), .Z(n13161) );
  XOR U13110 ( .A(n13167), .B(n13168), .Z(n12982) );
  AND U13111 ( .A(n324), .B(n13169), .Z(n13168) );
  XOR U13112 ( .A(n13170), .B(n13167), .Z(n13169) );
  XOR U13113 ( .A(n13171), .B(n13172), .Z(n13159) );
  AND U13114 ( .A(n13173), .B(n13174), .Z(n13172) );
  XOR U13115 ( .A(n13171), .B(n12997), .Z(n13174) );
  XOR U13116 ( .A(n13175), .B(n13176), .Z(n12997) );
  AND U13117 ( .A(n326), .B(n13177), .Z(n13176) );
  XOR U13118 ( .A(n13178), .B(n13175), .Z(n13177) );
  XNOR U13119 ( .A(n12994), .B(n13171), .Z(n13173) );
  XOR U13120 ( .A(n13179), .B(n13180), .Z(n12994) );
  AND U13121 ( .A(n324), .B(n13181), .Z(n13180) );
  XOR U13122 ( .A(n13182), .B(n13179), .Z(n13181) );
  XOR U13123 ( .A(n13183), .B(n13184), .Z(n13171) );
  AND U13124 ( .A(n13185), .B(n13186), .Z(n13184) );
  XOR U13125 ( .A(n13183), .B(n13009), .Z(n13186) );
  XOR U13126 ( .A(n13187), .B(n13188), .Z(n13009) );
  AND U13127 ( .A(n326), .B(n13189), .Z(n13188) );
  XOR U13128 ( .A(n13190), .B(n13187), .Z(n13189) );
  XNOR U13129 ( .A(n13006), .B(n13183), .Z(n13185) );
  XOR U13130 ( .A(n13191), .B(n13192), .Z(n13006) );
  AND U13131 ( .A(n324), .B(n13193), .Z(n13192) );
  XOR U13132 ( .A(n13194), .B(n13191), .Z(n13193) );
  XOR U13133 ( .A(n13195), .B(n13196), .Z(n13183) );
  AND U13134 ( .A(n13197), .B(n13198), .Z(n13196) );
  XOR U13135 ( .A(n13195), .B(n13021), .Z(n13198) );
  XOR U13136 ( .A(n13199), .B(n13200), .Z(n13021) );
  AND U13137 ( .A(n326), .B(n13201), .Z(n13200) );
  XOR U13138 ( .A(n13202), .B(n13199), .Z(n13201) );
  XNOR U13139 ( .A(n13018), .B(n13195), .Z(n13197) );
  XOR U13140 ( .A(n13203), .B(n13204), .Z(n13018) );
  AND U13141 ( .A(n324), .B(n13205), .Z(n13204) );
  XOR U13142 ( .A(n13206), .B(n13203), .Z(n13205) );
  XOR U13143 ( .A(n13207), .B(n13208), .Z(n13195) );
  AND U13144 ( .A(n13209), .B(n13210), .Z(n13208) );
  XOR U13145 ( .A(n13207), .B(n13033), .Z(n13210) );
  XOR U13146 ( .A(n13211), .B(n13212), .Z(n13033) );
  AND U13147 ( .A(n326), .B(n13213), .Z(n13212) );
  XOR U13148 ( .A(n13214), .B(n13211), .Z(n13213) );
  XNOR U13149 ( .A(n13030), .B(n13207), .Z(n13209) );
  XOR U13150 ( .A(n13215), .B(n13216), .Z(n13030) );
  AND U13151 ( .A(n324), .B(n13217), .Z(n13216) );
  XOR U13152 ( .A(n13218), .B(n13215), .Z(n13217) );
  XOR U13153 ( .A(n13219), .B(n13220), .Z(n13207) );
  AND U13154 ( .A(n13221), .B(n13222), .Z(n13220) );
  XOR U13155 ( .A(n13219), .B(n13045), .Z(n13222) );
  XOR U13156 ( .A(n13223), .B(n13224), .Z(n13045) );
  AND U13157 ( .A(n326), .B(n13225), .Z(n13224) );
  XOR U13158 ( .A(n13226), .B(n13223), .Z(n13225) );
  XNOR U13159 ( .A(n13042), .B(n13219), .Z(n13221) );
  XOR U13160 ( .A(n13227), .B(n13228), .Z(n13042) );
  AND U13161 ( .A(n324), .B(n13229), .Z(n13228) );
  XOR U13162 ( .A(n13230), .B(n13227), .Z(n13229) );
  XOR U13163 ( .A(n13231), .B(n13232), .Z(n13219) );
  AND U13164 ( .A(n13233), .B(n13234), .Z(n13232) );
  XOR U13165 ( .A(n13231), .B(n13057), .Z(n13234) );
  XOR U13166 ( .A(n13235), .B(n13236), .Z(n13057) );
  AND U13167 ( .A(n326), .B(n13237), .Z(n13236) );
  XOR U13168 ( .A(n13238), .B(n13235), .Z(n13237) );
  XNOR U13169 ( .A(n13054), .B(n13231), .Z(n13233) );
  XOR U13170 ( .A(n13239), .B(n13240), .Z(n13054) );
  AND U13171 ( .A(n324), .B(n13241), .Z(n13240) );
  XOR U13172 ( .A(n13242), .B(n13239), .Z(n13241) );
  XOR U13173 ( .A(n13243), .B(n13244), .Z(n13231) );
  AND U13174 ( .A(n13245), .B(n13246), .Z(n13244) );
  XOR U13175 ( .A(n13243), .B(n13069), .Z(n13246) );
  XOR U13176 ( .A(n13247), .B(n13248), .Z(n13069) );
  AND U13177 ( .A(n326), .B(n13249), .Z(n13248) );
  XOR U13178 ( .A(n13250), .B(n13247), .Z(n13249) );
  XNOR U13179 ( .A(n13066), .B(n13243), .Z(n13245) );
  XOR U13180 ( .A(n13251), .B(n13252), .Z(n13066) );
  AND U13181 ( .A(n324), .B(n13253), .Z(n13252) );
  XOR U13182 ( .A(n13254), .B(n13251), .Z(n13253) );
  XOR U13183 ( .A(n13255), .B(n13256), .Z(n13243) );
  AND U13184 ( .A(n13257), .B(n13258), .Z(n13256) );
  XOR U13185 ( .A(n13255), .B(n13081), .Z(n13258) );
  XOR U13186 ( .A(n13259), .B(n13260), .Z(n13081) );
  AND U13187 ( .A(n326), .B(n13261), .Z(n13260) );
  XOR U13188 ( .A(n13262), .B(n13259), .Z(n13261) );
  XNOR U13189 ( .A(n13078), .B(n13255), .Z(n13257) );
  XOR U13190 ( .A(n13263), .B(n13264), .Z(n13078) );
  AND U13191 ( .A(n324), .B(n13265), .Z(n13264) );
  XOR U13192 ( .A(n13266), .B(n13263), .Z(n13265) );
  XOR U13193 ( .A(n13267), .B(n13268), .Z(n13255) );
  AND U13194 ( .A(n13269), .B(n13270), .Z(n13268) );
  XOR U13195 ( .A(n13267), .B(n13093), .Z(n13270) );
  XOR U13196 ( .A(n13271), .B(n13272), .Z(n13093) );
  AND U13197 ( .A(n326), .B(n13273), .Z(n13272) );
  XOR U13198 ( .A(n13274), .B(n13271), .Z(n13273) );
  XNOR U13199 ( .A(n13090), .B(n13267), .Z(n13269) );
  XOR U13200 ( .A(n13275), .B(n13276), .Z(n13090) );
  AND U13201 ( .A(n324), .B(n13277), .Z(n13276) );
  XOR U13202 ( .A(n13278), .B(n13275), .Z(n13277) );
  XOR U13203 ( .A(n13279), .B(n13280), .Z(n13267) );
  AND U13204 ( .A(n13281), .B(n13282), .Z(n13280) );
  XOR U13205 ( .A(n13279), .B(n13105), .Z(n13282) );
  XOR U13206 ( .A(n13283), .B(n13284), .Z(n13105) );
  AND U13207 ( .A(n326), .B(n13285), .Z(n13284) );
  XOR U13208 ( .A(n13286), .B(n13283), .Z(n13285) );
  XNOR U13209 ( .A(n13102), .B(n13279), .Z(n13281) );
  XOR U13210 ( .A(n13287), .B(n13288), .Z(n13102) );
  AND U13211 ( .A(n324), .B(n13289), .Z(n13288) );
  XOR U13212 ( .A(n13290), .B(n13287), .Z(n13289) );
  XOR U13213 ( .A(n13291), .B(n13292), .Z(n13279) );
  AND U13214 ( .A(n13293), .B(n13294), .Z(n13292) );
  XOR U13215 ( .A(n13291), .B(n13117), .Z(n13294) );
  XOR U13216 ( .A(n13295), .B(n13296), .Z(n13117) );
  AND U13217 ( .A(n326), .B(n13297), .Z(n13296) );
  XOR U13218 ( .A(n13298), .B(n13295), .Z(n13297) );
  XNOR U13219 ( .A(n13114), .B(n13291), .Z(n13293) );
  XOR U13220 ( .A(n13299), .B(n13300), .Z(n13114) );
  AND U13221 ( .A(n324), .B(n13301), .Z(n13300) );
  XOR U13222 ( .A(n13302), .B(n13299), .Z(n13301) );
  XOR U13223 ( .A(n13303), .B(n13304), .Z(n13291) );
  AND U13224 ( .A(n13305), .B(n13306), .Z(n13304) );
  XOR U13225 ( .A(n13129), .B(n13303), .Z(n13306) );
  XOR U13226 ( .A(n13307), .B(n13308), .Z(n13129) );
  AND U13227 ( .A(n326), .B(n13309), .Z(n13308) );
  XOR U13228 ( .A(n13307), .B(n13310), .Z(n13309) );
  XNOR U13229 ( .A(n13303), .B(n13126), .Z(n13305) );
  XOR U13230 ( .A(n13311), .B(n13312), .Z(n13126) );
  AND U13231 ( .A(n324), .B(n13313), .Z(n13312) );
  XOR U13232 ( .A(n13311), .B(n13314), .Z(n13313) );
  XOR U13233 ( .A(n13315), .B(n13316), .Z(n13303) );
  AND U13234 ( .A(n13317), .B(n13318), .Z(n13316) );
  XNOR U13235 ( .A(n13319), .B(n13142), .Z(n13318) );
  XOR U13236 ( .A(n13320), .B(n13321), .Z(n13142) );
  AND U13237 ( .A(n326), .B(n13322), .Z(n13321) );
  XOR U13238 ( .A(n13323), .B(n13320), .Z(n13322) );
  XNOR U13239 ( .A(n13139), .B(n13315), .Z(n13317) );
  XOR U13240 ( .A(n13324), .B(n13325), .Z(n13139) );
  AND U13241 ( .A(n324), .B(n13326), .Z(n13325) );
  XOR U13242 ( .A(n13327), .B(n13324), .Z(n13326) );
  IV U13243 ( .A(n13319), .Z(n13315) );
  AND U13244 ( .A(n13147), .B(n13150), .Z(n13319) );
  XNOR U13245 ( .A(n13328), .B(n13329), .Z(n13150) );
  AND U13246 ( .A(n326), .B(n13330), .Z(n13329) );
  XNOR U13247 ( .A(n13331), .B(n13328), .Z(n13330) );
  XOR U13248 ( .A(n13332), .B(n13333), .Z(n326) );
  AND U13249 ( .A(n13334), .B(n13335), .Z(n13333) );
  XNOR U13250 ( .A(n13155), .B(n13332), .Z(n13335) );
  AND U13251 ( .A(p_input[255]), .B(p_input[239]), .Z(n13155) );
  XOR U13252 ( .A(n13332), .B(n13156), .Z(n13334) );
  AND U13253 ( .A(p_input[223]), .B(p_input[207]), .Z(n13156) );
  XOR U13254 ( .A(n13336), .B(n13337), .Z(n13332) );
  AND U13255 ( .A(n13338), .B(n13339), .Z(n13337) );
  XOR U13256 ( .A(n13336), .B(n13166), .Z(n13339) );
  XNOR U13257 ( .A(p_input[238]), .B(n13340), .Z(n13166) );
  AND U13258 ( .A(n526), .B(n13341), .Z(n13340) );
  XOR U13259 ( .A(p_input[254]), .B(p_input[238]), .Z(n13341) );
  XNOR U13260 ( .A(n13163), .B(n13336), .Z(n13338) );
  XOR U13261 ( .A(n13342), .B(n13343), .Z(n13163) );
  AND U13262 ( .A(n524), .B(n13344), .Z(n13343) );
  XOR U13263 ( .A(p_input[222]), .B(p_input[206]), .Z(n13344) );
  XOR U13264 ( .A(n13345), .B(n13346), .Z(n13336) );
  AND U13265 ( .A(n13347), .B(n13348), .Z(n13346) );
  XOR U13266 ( .A(n13345), .B(n13178), .Z(n13348) );
  XNOR U13267 ( .A(p_input[237]), .B(n13349), .Z(n13178) );
  AND U13268 ( .A(n526), .B(n13350), .Z(n13349) );
  XOR U13269 ( .A(p_input[253]), .B(p_input[237]), .Z(n13350) );
  XNOR U13270 ( .A(n13175), .B(n13345), .Z(n13347) );
  XOR U13271 ( .A(n13351), .B(n13352), .Z(n13175) );
  AND U13272 ( .A(n524), .B(n13353), .Z(n13352) );
  XOR U13273 ( .A(p_input[221]), .B(p_input[205]), .Z(n13353) );
  XOR U13274 ( .A(n13354), .B(n13355), .Z(n13345) );
  AND U13275 ( .A(n13356), .B(n13357), .Z(n13355) );
  XOR U13276 ( .A(n13354), .B(n13190), .Z(n13357) );
  XNOR U13277 ( .A(p_input[236]), .B(n13358), .Z(n13190) );
  AND U13278 ( .A(n526), .B(n13359), .Z(n13358) );
  XOR U13279 ( .A(p_input[252]), .B(p_input[236]), .Z(n13359) );
  XNOR U13280 ( .A(n13187), .B(n13354), .Z(n13356) );
  XOR U13281 ( .A(n13360), .B(n13361), .Z(n13187) );
  AND U13282 ( .A(n524), .B(n13362), .Z(n13361) );
  XOR U13283 ( .A(p_input[220]), .B(p_input[204]), .Z(n13362) );
  XOR U13284 ( .A(n13363), .B(n13364), .Z(n13354) );
  AND U13285 ( .A(n13365), .B(n13366), .Z(n13364) );
  XOR U13286 ( .A(n13363), .B(n13202), .Z(n13366) );
  XNOR U13287 ( .A(p_input[235]), .B(n13367), .Z(n13202) );
  AND U13288 ( .A(n526), .B(n13368), .Z(n13367) );
  XOR U13289 ( .A(p_input[251]), .B(p_input[235]), .Z(n13368) );
  XNOR U13290 ( .A(n13199), .B(n13363), .Z(n13365) );
  XOR U13291 ( .A(n13369), .B(n13370), .Z(n13199) );
  AND U13292 ( .A(n524), .B(n13371), .Z(n13370) );
  XOR U13293 ( .A(p_input[219]), .B(p_input[203]), .Z(n13371) );
  XOR U13294 ( .A(n13372), .B(n13373), .Z(n13363) );
  AND U13295 ( .A(n13374), .B(n13375), .Z(n13373) );
  XOR U13296 ( .A(n13372), .B(n13214), .Z(n13375) );
  XNOR U13297 ( .A(p_input[234]), .B(n13376), .Z(n13214) );
  AND U13298 ( .A(n526), .B(n13377), .Z(n13376) );
  XOR U13299 ( .A(p_input[250]), .B(p_input[234]), .Z(n13377) );
  XNOR U13300 ( .A(n13211), .B(n13372), .Z(n13374) );
  XOR U13301 ( .A(n13378), .B(n13379), .Z(n13211) );
  AND U13302 ( .A(n524), .B(n13380), .Z(n13379) );
  XOR U13303 ( .A(p_input[218]), .B(p_input[202]), .Z(n13380) );
  XOR U13304 ( .A(n13381), .B(n13382), .Z(n13372) );
  AND U13305 ( .A(n13383), .B(n13384), .Z(n13382) );
  XOR U13306 ( .A(n13381), .B(n13226), .Z(n13384) );
  XNOR U13307 ( .A(p_input[233]), .B(n13385), .Z(n13226) );
  AND U13308 ( .A(n526), .B(n13386), .Z(n13385) );
  XOR U13309 ( .A(p_input[249]), .B(p_input[233]), .Z(n13386) );
  XNOR U13310 ( .A(n13223), .B(n13381), .Z(n13383) );
  XOR U13311 ( .A(n13387), .B(n13388), .Z(n13223) );
  AND U13312 ( .A(n524), .B(n13389), .Z(n13388) );
  XOR U13313 ( .A(p_input[217]), .B(p_input[201]), .Z(n13389) );
  XOR U13314 ( .A(n13390), .B(n13391), .Z(n13381) );
  AND U13315 ( .A(n13392), .B(n13393), .Z(n13391) );
  XOR U13316 ( .A(n13390), .B(n13238), .Z(n13393) );
  XNOR U13317 ( .A(p_input[232]), .B(n13394), .Z(n13238) );
  AND U13318 ( .A(n526), .B(n13395), .Z(n13394) );
  XOR U13319 ( .A(p_input[248]), .B(p_input[232]), .Z(n13395) );
  XNOR U13320 ( .A(n13235), .B(n13390), .Z(n13392) );
  XOR U13321 ( .A(n13396), .B(n13397), .Z(n13235) );
  AND U13322 ( .A(n524), .B(n13398), .Z(n13397) );
  XOR U13323 ( .A(p_input[216]), .B(p_input[200]), .Z(n13398) );
  XOR U13324 ( .A(n13399), .B(n13400), .Z(n13390) );
  AND U13325 ( .A(n13401), .B(n13402), .Z(n13400) );
  XOR U13326 ( .A(n13399), .B(n13250), .Z(n13402) );
  XNOR U13327 ( .A(p_input[231]), .B(n13403), .Z(n13250) );
  AND U13328 ( .A(n526), .B(n13404), .Z(n13403) );
  XOR U13329 ( .A(p_input[247]), .B(p_input[231]), .Z(n13404) );
  XNOR U13330 ( .A(n13247), .B(n13399), .Z(n13401) );
  XOR U13331 ( .A(n13405), .B(n13406), .Z(n13247) );
  AND U13332 ( .A(n524), .B(n13407), .Z(n13406) );
  XOR U13333 ( .A(p_input[215]), .B(p_input[199]), .Z(n13407) );
  XOR U13334 ( .A(n13408), .B(n13409), .Z(n13399) );
  AND U13335 ( .A(n13410), .B(n13411), .Z(n13409) );
  XOR U13336 ( .A(n13408), .B(n13262), .Z(n13411) );
  XNOR U13337 ( .A(p_input[230]), .B(n13412), .Z(n13262) );
  AND U13338 ( .A(n526), .B(n13413), .Z(n13412) );
  XOR U13339 ( .A(p_input[246]), .B(p_input[230]), .Z(n13413) );
  XNOR U13340 ( .A(n13259), .B(n13408), .Z(n13410) );
  XOR U13341 ( .A(n13414), .B(n13415), .Z(n13259) );
  AND U13342 ( .A(n524), .B(n13416), .Z(n13415) );
  XOR U13343 ( .A(p_input[214]), .B(p_input[198]), .Z(n13416) );
  XOR U13344 ( .A(n13417), .B(n13418), .Z(n13408) );
  AND U13345 ( .A(n13419), .B(n13420), .Z(n13418) );
  XOR U13346 ( .A(n13417), .B(n13274), .Z(n13420) );
  XNOR U13347 ( .A(p_input[229]), .B(n13421), .Z(n13274) );
  AND U13348 ( .A(n526), .B(n13422), .Z(n13421) );
  XOR U13349 ( .A(p_input[245]), .B(p_input[229]), .Z(n13422) );
  XNOR U13350 ( .A(n13271), .B(n13417), .Z(n13419) );
  XOR U13351 ( .A(n13423), .B(n13424), .Z(n13271) );
  AND U13352 ( .A(n524), .B(n13425), .Z(n13424) );
  XOR U13353 ( .A(p_input[213]), .B(p_input[197]), .Z(n13425) );
  XOR U13354 ( .A(n13426), .B(n13427), .Z(n13417) );
  AND U13355 ( .A(n13428), .B(n13429), .Z(n13427) );
  XOR U13356 ( .A(n13426), .B(n13286), .Z(n13429) );
  XNOR U13357 ( .A(p_input[228]), .B(n13430), .Z(n13286) );
  AND U13358 ( .A(n526), .B(n13431), .Z(n13430) );
  XOR U13359 ( .A(p_input[244]), .B(p_input[228]), .Z(n13431) );
  XNOR U13360 ( .A(n13283), .B(n13426), .Z(n13428) );
  XOR U13361 ( .A(n13432), .B(n13433), .Z(n13283) );
  AND U13362 ( .A(n524), .B(n13434), .Z(n13433) );
  XOR U13363 ( .A(p_input[212]), .B(p_input[196]), .Z(n13434) );
  XOR U13364 ( .A(n13435), .B(n13436), .Z(n13426) );
  AND U13365 ( .A(n13437), .B(n13438), .Z(n13436) );
  XOR U13366 ( .A(n13435), .B(n13298), .Z(n13438) );
  XNOR U13367 ( .A(p_input[227]), .B(n13439), .Z(n13298) );
  AND U13368 ( .A(n526), .B(n13440), .Z(n13439) );
  XOR U13369 ( .A(p_input[243]), .B(p_input[227]), .Z(n13440) );
  XNOR U13370 ( .A(n13295), .B(n13435), .Z(n13437) );
  XOR U13371 ( .A(n13441), .B(n13442), .Z(n13295) );
  AND U13372 ( .A(n524), .B(n13443), .Z(n13442) );
  XOR U13373 ( .A(p_input[211]), .B(p_input[195]), .Z(n13443) );
  XOR U13374 ( .A(n13444), .B(n13445), .Z(n13435) );
  AND U13375 ( .A(n13446), .B(n13447), .Z(n13445) );
  XOR U13376 ( .A(n13310), .B(n13444), .Z(n13447) );
  XNOR U13377 ( .A(p_input[226]), .B(n13448), .Z(n13310) );
  AND U13378 ( .A(n526), .B(n13449), .Z(n13448) );
  XOR U13379 ( .A(p_input[242]), .B(p_input[226]), .Z(n13449) );
  XNOR U13380 ( .A(n13444), .B(n13307), .Z(n13446) );
  XOR U13381 ( .A(n13450), .B(n13451), .Z(n13307) );
  AND U13382 ( .A(n524), .B(n13452), .Z(n13451) );
  XOR U13383 ( .A(p_input[210]), .B(p_input[194]), .Z(n13452) );
  XOR U13384 ( .A(n13453), .B(n13454), .Z(n13444) );
  AND U13385 ( .A(n13455), .B(n13456), .Z(n13454) );
  XNOR U13386 ( .A(n13457), .B(n13323), .Z(n13456) );
  XNOR U13387 ( .A(p_input[225]), .B(n13458), .Z(n13323) );
  AND U13388 ( .A(n526), .B(n13459), .Z(n13458) );
  XNOR U13389 ( .A(p_input[241]), .B(n13460), .Z(n13459) );
  IV U13390 ( .A(p_input[225]), .Z(n13460) );
  XNOR U13391 ( .A(n13320), .B(n13453), .Z(n13455) );
  XNOR U13392 ( .A(p_input[193]), .B(n13461), .Z(n13320) );
  AND U13393 ( .A(n524), .B(n13462), .Z(n13461) );
  XOR U13394 ( .A(p_input[209]), .B(p_input[193]), .Z(n13462) );
  IV U13395 ( .A(n13457), .Z(n13453) );
  AND U13396 ( .A(n13328), .B(n13331), .Z(n13457) );
  XOR U13397 ( .A(p_input[224]), .B(n13463), .Z(n13331) );
  AND U13398 ( .A(n526), .B(n13464), .Z(n13463) );
  XOR U13399 ( .A(p_input[240]), .B(p_input[224]), .Z(n13464) );
  XOR U13400 ( .A(n13465), .B(n13466), .Z(n526) );
  AND U13401 ( .A(n13467), .B(n13468), .Z(n13466) );
  XNOR U13402 ( .A(p_input[255]), .B(n13465), .Z(n13468) );
  XOR U13403 ( .A(n13465), .B(p_input[239]), .Z(n13467) );
  XOR U13404 ( .A(n13469), .B(n13470), .Z(n13465) );
  AND U13405 ( .A(n13471), .B(n13472), .Z(n13470) );
  XNOR U13406 ( .A(p_input[254]), .B(n13469), .Z(n13472) );
  XOR U13407 ( .A(n13469), .B(p_input[238]), .Z(n13471) );
  XOR U13408 ( .A(n13473), .B(n13474), .Z(n13469) );
  AND U13409 ( .A(n13475), .B(n13476), .Z(n13474) );
  XNOR U13410 ( .A(p_input[253]), .B(n13473), .Z(n13476) );
  XOR U13411 ( .A(n13473), .B(p_input[237]), .Z(n13475) );
  XOR U13412 ( .A(n13477), .B(n13478), .Z(n13473) );
  AND U13413 ( .A(n13479), .B(n13480), .Z(n13478) );
  XNOR U13414 ( .A(p_input[252]), .B(n13477), .Z(n13480) );
  XOR U13415 ( .A(n13477), .B(p_input[236]), .Z(n13479) );
  XOR U13416 ( .A(n13481), .B(n13482), .Z(n13477) );
  AND U13417 ( .A(n13483), .B(n13484), .Z(n13482) );
  XNOR U13418 ( .A(p_input[251]), .B(n13481), .Z(n13484) );
  XOR U13419 ( .A(n13481), .B(p_input[235]), .Z(n13483) );
  XOR U13420 ( .A(n13485), .B(n13486), .Z(n13481) );
  AND U13421 ( .A(n13487), .B(n13488), .Z(n13486) );
  XNOR U13422 ( .A(p_input[250]), .B(n13485), .Z(n13488) );
  XOR U13423 ( .A(n13485), .B(p_input[234]), .Z(n13487) );
  XOR U13424 ( .A(n13489), .B(n13490), .Z(n13485) );
  AND U13425 ( .A(n13491), .B(n13492), .Z(n13490) );
  XNOR U13426 ( .A(p_input[249]), .B(n13489), .Z(n13492) );
  XOR U13427 ( .A(n13489), .B(p_input[233]), .Z(n13491) );
  XOR U13428 ( .A(n13493), .B(n13494), .Z(n13489) );
  AND U13429 ( .A(n13495), .B(n13496), .Z(n13494) );
  XNOR U13430 ( .A(p_input[248]), .B(n13493), .Z(n13496) );
  XOR U13431 ( .A(n13493), .B(p_input[232]), .Z(n13495) );
  XOR U13432 ( .A(n13497), .B(n13498), .Z(n13493) );
  AND U13433 ( .A(n13499), .B(n13500), .Z(n13498) );
  XNOR U13434 ( .A(p_input[247]), .B(n13497), .Z(n13500) );
  XOR U13435 ( .A(n13497), .B(p_input[231]), .Z(n13499) );
  XOR U13436 ( .A(n13501), .B(n13502), .Z(n13497) );
  AND U13437 ( .A(n13503), .B(n13504), .Z(n13502) );
  XNOR U13438 ( .A(p_input[246]), .B(n13501), .Z(n13504) );
  XOR U13439 ( .A(n13501), .B(p_input[230]), .Z(n13503) );
  XOR U13440 ( .A(n13505), .B(n13506), .Z(n13501) );
  AND U13441 ( .A(n13507), .B(n13508), .Z(n13506) );
  XNOR U13442 ( .A(p_input[245]), .B(n13505), .Z(n13508) );
  XOR U13443 ( .A(n13505), .B(p_input[229]), .Z(n13507) );
  XOR U13444 ( .A(n13509), .B(n13510), .Z(n13505) );
  AND U13445 ( .A(n13511), .B(n13512), .Z(n13510) );
  XNOR U13446 ( .A(p_input[244]), .B(n13509), .Z(n13512) );
  XOR U13447 ( .A(n13509), .B(p_input[228]), .Z(n13511) );
  XOR U13448 ( .A(n13513), .B(n13514), .Z(n13509) );
  AND U13449 ( .A(n13515), .B(n13516), .Z(n13514) );
  XNOR U13450 ( .A(p_input[243]), .B(n13513), .Z(n13516) );
  XOR U13451 ( .A(n13513), .B(p_input[227]), .Z(n13515) );
  XOR U13452 ( .A(n13517), .B(n13518), .Z(n13513) );
  AND U13453 ( .A(n13519), .B(n13520), .Z(n13518) );
  XNOR U13454 ( .A(p_input[242]), .B(n13517), .Z(n13520) );
  XOR U13455 ( .A(n13517), .B(p_input[226]), .Z(n13519) );
  XNOR U13456 ( .A(n13521), .B(n13522), .Z(n13517) );
  AND U13457 ( .A(n13523), .B(n13524), .Z(n13522) );
  XOR U13458 ( .A(p_input[241]), .B(n13521), .Z(n13524) );
  XNOR U13459 ( .A(p_input[225]), .B(n13521), .Z(n13523) );
  AND U13460 ( .A(p_input[240]), .B(n13525), .Z(n13521) );
  IV U13461 ( .A(p_input[224]), .Z(n13525) );
  XNOR U13462 ( .A(p_input[192]), .B(n13526), .Z(n13328) );
  AND U13463 ( .A(n524), .B(n13527), .Z(n13526) );
  XOR U13464 ( .A(p_input[208]), .B(p_input[192]), .Z(n13527) );
  XOR U13465 ( .A(n13528), .B(n13529), .Z(n524) );
  AND U13466 ( .A(n13530), .B(n13531), .Z(n13529) );
  XNOR U13467 ( .A(p_input[223]), .B(n13528), .Z(n13531) );
  XOR U13468 ( .A(n13528), .B(p_input[207]), .Z(n13530) );
  XOR U13469 ( .A(n13532), .B(n13533), .Z(n13528) );
  AND U13470 ( .A(n13534), .B(n13535), .Z(n13533) );
  XNOR U13471 ( .A(p_input[222]), .B(n13532), .Z(n13535) );
  XNOR U13472 ( .A(n13532), .B(n13342), .Z(n13534) );
  IV U13473 ( .A(p_input[206]), .Z(n13342) );
  XOR U13474 ( .A(n13536), .B(n13537), .Z(n13532) );
  AND U13475 ( .A(n13538), .B(n13539), .Z(n13537) );
  XNOR U13476 ( .A(p_input[221]), .B(n13536), .Z(n13539) );
  XNOR U13477 ( .A(n13536), .B(n13351), .Z(n13538) );
  IV U13478 ( .A(p_input[205]), .Z(n13351) );
  XOR U13479 ( .A(n13540), .B(n13541), .Z(n13536) );
  AND U13480 ( .A(n13542), .B(n13543), .Z(n13541) );
  XNOR U13481 ( .A(p_input[220]), .B(n13540), .Z(n13543) );
  XNOR U13482 ( .A(n13540), .B(n13360), .Z(n13542) );
  IV U13483 ( .A(p_input[204]), .Z(n13360) );
  XOR U13484 ( .A(n13544), .B(n13545), .Z(n13540) );
  AND U13485 ( .A(n13546), .B(n13547), .Z(n13545) );
  XNOR U13486 ( .A(p_input[219]), .B(n13544), .Z(n13547) );
  XNOR U13487 ( .A(n13544), .B(n13369), .Z(n13546) );
  IV U13488 ( .A(p_input[203]), .Z(n13369) );
  XOR U13489 ( .A(n13548), .B(n13549), .Z(n13544) );
  AND U13490 ( .A(n13550), .B(n13551), .Z(n13549) );
  XNOR U13491 ( .A(p_input[218]), .B(n13548), .Z(n13551) );
  XNOR U13492 ( .A(n13548), .B(n13378), .Z(n13550) );
  IV U13493 ( .A(p_input[202]), .Z(n13378) );
  XOR U13494 ( .A(n13552), .B(n13553), .Z(n13548) );
  AND U13495 ( .A(n13554), .B(n13555), .Z(n13553) );
  XNOR U13496 ( .A(p_input[217]), .B(n13552), .Z(n13555) );
  XNOR U13497 ( .A(n13552), .B(n13387), .Z(n13554) );
  IV U13498 ( .A(p_input[201]), .Z(n13387) );
  XOR U13499 ( .A(n13556), .B(n13557), .Z(n13552) );
  AND U13500 ( .A(n13558), .B(n13559), .Z(n13557) );
  XNOR U13501 ( .A(p_input[216]), .B(n13556), .Z(n13559) );
  XNOR U13502 ( .A(n13556), .B(n13396), .Z(n13558) );
  IV U13503 ( .A(p_input[200]), .Z(n13396) );
  XOR U13504 ( .A(n13560), .B(n13561), .Z(n13556) );
  AND U13505 ( .A(n13562), .B(n13563), .Z(n13561) );
  XNOR U13506 ( .A(p_input[215]), .B(n13560), .Z(n13563) );
  XNOR U13507 ( .A(n13560), .B(n13405), .Z(n13562) );
  IV U13508 ( .A(p_input[199]), .Z(n13405) );
  XOR U13509 ( .A(n13564), .B(n13565), .Z(n13560) );
  AND U13510 ( .A(n13566), .B(n13567), .Z(n13565) );
  XNOR U13511 ( .A(p_input[214]), .B(n13564), .Z(n13567) );
  XNOR U13512 ( .A(n13564), .B(n13414), .Z(n13566) );
  IV U13513 ( .A(p_input[198]), .Z(n13414) );
  XOR U13514 ( .A(n13568), .B(n13569), .Z(n13564) );
  AND U13515 ( .A(n13570), .B(n13571), .Z(n13569) );
  XNOR U13516 ( .A(p_input[213]), .B(n13568), .Z(n13571) );
  XNOR U13517 ( .A(n13568), .B(n13423), .Z(n13570) );
  IV U13518 ( .A(p_input[197]), .Z(n13423) );
  XOR U13519 ( .A(n13572), .B(n13573), .Z(n13568) );
  AND U13520 ( .A(n13574), .B(n13575), .Z(n13573) );
  XNOR U13521 ( .A(p_input[212]), .B(n13572), .Z(n13575) );
  XNOR U13522 ( .A(n13572), .B(n13432), .Z(n13574) );
  IV U13523 ( .A(p_input[196]), .Z(n13432) );
  XOR U13524 ( .A(n13576), .B(n13577), .Z(n13572) );
  AND U13525 ( .A(n13578), .B(n13579), .Z(n13577) );
  XNOR U13526 ( .A(p_input[211]), .B(n13576), .Z(n13579) );
  XNOR U13527 ( .A(n13576), .B(n13441), .Z(n13578) );
  IV U13528 ( .A(p_input[195]), .Z(n13441) );
  XOR U13529 ( .A(n13580), .B(n13581), .Z(n13576) );
  AND U13530 ( .A(n13582), .B(n13583), .Z(n13581) );
  XNOR U13531 ( .A(p_input[210]), .B(n13580), .Z(n13583) );
  XNOR U13532 ( .A(n13580), .B(n13450), .Z(n13582) );
  IV U13533 ( .A(p_input[194]), .Z(n13450) );
  XNOR U13534 ( .A(n13584), .B(n13585), .Z(n13580) );
  AND U13535 ( .A(n13586), .B(n13587), .Z(n13585) );
  XOR U13536 ( .A(p_input[209]), .B(n13584), .Z(n13587) );
  XNOR U13537 ( .A(p_input[193]), .B(n13584), .Z(n13586) );
  AND U13538 ( .A(p_input[208]), .B(n13588), .Z(n13584) );
  IV U13539 ( .A(p_input[192]), .Z(n13588) );
  XOR U13540 ( .A(n13589), .B(n13590), .Z(n13147) );
  AND U13541 ( .A(n324), .B(n13591), .Z(n13590) );
  XNOR U13542 ( .A(n13592), .B(n13589), .Z(n13591) );
  XOR U13543 ( .A(n13593), .B(n13594), .Z(n324) );
  AND U13544 ( .A(n13595), .B(n13596), .Z(n13594) );
  XNOR U13545 ( .A(n13157), .B(n13593), .Z(n13596) );
  AND U13546 ( .A(p_input[191]), .B(p_input[175]), .Z(n13157) );
  XOR U13547 ( .A(n13593), .B(n13158), .Z(n13595) );
  AND U13548 ( .A(p_input[159]), .B(p_input[143]), .Z(n13158) );
  XOR U13549 ( .A(n13597), .B(n13598), .Z(n13593) );
  AND U13550 ( .A(n13599), .B(n13600), .Z(n13598) );
  XOR U13551 ( .A(n13597), .B(n13170), .Z(n13600) );
  XNOR U13552 ( .A(p_input[174]), .B(n13601), .Z(n13170) );
  AND U13553 ( .A(n530), .B(n13602), .Z(n13601) );
  XOR U13554 ( .A(p_input[190]), .B(p_input[174]), .Z(n13602) );
  XNOR U13555 ( .A(n13167), .B(n13597), .Z(n13599) );
  XOR U13556 ( .A(n13603), .B(n13604), .Z(n13167) );
  AND U13557 ( .A(n527), .B(n13605), .Z(n13604) );
  XOR U13558 ( .A(p_input[158]), .B(p_input[142]), .Z(n13605) );
  XOR U13559 ( .A(n13606), .B(n13607), .Z(n13597) );
  AND U13560 ( .A(n13608), .B(n13609), .Z(n13607) );
  XOR U13561 ( .A(n13606), .B(n13182), .Z(n13609) );
  XNOR U13562 ( .A(p_input[173]), .B(n13610), .Z(n13182) );
  AND U13563 ( .A(n530), .B(n13611), .Z(n13610) );
  XOR U13564 ( .A(p_input[189]), .B(p_input[173]), .Z(n13611) );
  XNOR U13565 ( .A(n13179), .B(n13606), .Z(n13608) );
  XOR U13566 ( .A(n13612), .B(n13613), .Z(n13179) );
  AND U13567 ( .A(n527), .B(n13614), .Z(n13613) );
  XOR U13568 ( .A(p_input[157]), .B(p_input[141]), .Z(n13614) );
  XOR U13569 ( .A(n13615), .B(n13616), .Z(n13606) );
  AND U13570 ( .A(n13617), .B(n13618), .Z(n13616) );
  XOR U13571 ( .A(n13615), .B(n13194), .Z(n13618) );
  XNOR U13572 ( .A(p_input[172]), .B(n13619), .Z(n13194) );
  AND U13573 ( .A(n530), .B(n13620), .Z(n13619) );
  XOR U13574 ( .A(p_input[188]), .B(p_input[172]), .Z(n13620) );
  XNOR U13575 ( .A(n13191), .B(n13615), .Z(n13617) );
  XOR U13576 ( .A(n13621), .B(n13622), .Z(n13191) );
  AND U13577 ( .A(n527), .B(n13623), .Z(n13622) );
  XOR U13578 ( .A(p_input[156]), .B(p_input[140]), .Z(n13623) );
  XOR U13579 ( .A(n13624), .B(n13625), .Z(n13615) );
  AND U13580 ( .A(n13626), .B(n13627), .Z(n13625) );
  XOR U13581 ( .A(n13624), .B(n13206), .Z(n13627) );
  XNOR U13582 ( .A(p_input[171]), .B(n13628), .Z(n13206) );
  AND U13583 ( .A(n530), .B(n13629), .Z(n13628) );
  XOR U13584 ( .A(p_input[187]), .B(p_input[171]), .Z(n13629) );
  XNOR U13585 ( .A(n13203), .B(n13624), .Z(n13626) );
  XOR U13586 ( .A(n13630), .B(n13631), .Z(n13203) );
  AND U13587 ( .A(n527), .B(n13632), .Z(n13631) );
  XOR U13588 ( .A(p_input[155]), .B(p_input[139]), .Z(n13632) );
  XOR U13589 ( .A(n13633), .B(n13634), .Z(n13624) );
  AND U13590 ( .A(n13635), .B(n13636), .Z(n13634) );
  XOR U13591 ( .A(n13633), .B(n13218), .Z(n13636) );
  XNOR U13592 ( .A(p_input[170]), .B(n13637), .Z(n13218) );
  AND U13593 ( .A(n530), .B(n13638), .Z(n13637) );
  XOR U13594 ( .A(p_input[186]), .B(p_input[170]), .Z(n13638) );
  XNOR U13595 ( .A(n13215), .B(n13633), .Z(n13635) );
  XOR U13596 ( .A(n13639), .B(n13640), .Z(n13215) );
  AND U13597 ( .A(n527), .B(n13641), .Z(n13640) );
  XOR U13598 ( .A(p_input[154]), .B(p_input[138]), .Z(n13641) );
  XOR U13599 ( .A(n13642), .B(n13643), .Z(n13633) );
  AND U13600 ( .A(n13644), .B(n13645), .Z(n13643) );
  XOR U13601 ( .A(n13642), .B(n13230), .Z(n13645) );
  XNOR U13602 ( .A(p_input[169]), .B(n13646), .Z(n13230) );
  AND U13603 ( .A(n530), .B(n13647), .Z(n13646) );
  XOR U13604 ( .A(p_input[185]), .B(p_input[169]), .Z(n13647) );
  XNOR U13605 ( .A(n13227), .B(n13642), .Z(n13644) );
  XOR U13606 ( .A(n13648), .B(n13649), .Z(n13227) );
  AND U13607 ( .A(n527), .B(n13650), .Z(n13649) );
  XOR U13608 ( .A(p_input[153]), .B(p_input[137]), .Z(n13650) );
  XOR U13609 ( .A(n13651), .B(n13652), .Z(n13642) );
  AND U13610 ( .A(n13653), .B(n13654), .Z(n13652) );
  XOR U13611 ( .A(n13651), .B(n13242), .Z(n13654) );
  XNOR U13612 ( .A(p_input[168]), .B(n13655), .Z(n13242) );
  AND U13613 ( .A(n530), .B(n13656), .Z(n13655) );
  XOR U13614 ( .A(p_input[184]), .B(p_input[168]), .Z(n13656) );
  XNOR U13615 ( .A(n13239), .B(n13651), .Z(n13653) );
  XOR U13616 ( .A(n13657), .B(n13658), .Z(n13239) );
  AND U13617 ( .A(n527), .B(n13659), .Z(n13658) );
  XOR U13618 ( .A(p_input[152]), .B(p_input[136]), .Z(n13659) );
  XOR U13619 ( .A(n13660), .B(n13661), .Z(n13651) );
  AND U13620 ( .A(n13662), .B(n13663), .Z(n13661) );
  XOR U13621 ( .A(n13660), .B(n13254), .Z(n13663) );
  XNOR U13622 ( .A(p_input[167]), .B(n13664), .Z(n13254) );
  AND U13623 ( .A(n530), .B(n13665), .Z(n13664) );
  XOR U13624 ( .A(p_input[183]), .B(p_input[167]), .Z(n13665) );
  XNOR U13625 ( .A(n13251), .B(n13660), .Z(n13662) );
  XOR U13626 ( .A(n13666), .B(n13667), .Z(n13251) );
  AND U13627 ( .A(n527), .B(n13668), .Z(n13667) );
  XOR U13628 ( .A(p_input[151]), .B(p_input[135]), .Z(n13668) );
  XOR U13629 ( .A(n13669), .B(n13670), .Z(n13660) );
  AND U13630 ( .A(n13671), .B(n13672), .Z(n13670) );
  XOR U13631 ( .A(n13669), .B(n13266), .Z(n13672) );
  XNOR U13632 ( .A(p_input[166]), .B(n13673), .Z(n13266) );
  AND U13633 ( .A(n530), .B(n13674), .Z(n13673) );
  XOR U13634 ( .A(p_input[182]), .B(p_input[166]), .Z(n13674) );
  XNOR U13635 ( .A(n13263), .B(n13669), .Z(n13671) );
  XOR U13636 ( .A(n13675), .B(n13676), .Z(n13263) );
  AND U13637 ( .A(n527), .B(n13677), .Z(n13676) );
  XOR U13638 ( .A(p_input[150]), .B(p_input[134]), .Z(n13677) );
  XOR U13639 ( .A(n13678), .B(n13679), .Z(n13669) );
  AND U13640 ( .A(n13680), .B(n13681), .Z(n13679) );
  XOR U13641 ( .A(n13678), .B(n13278), .Z(n13681) );
  XNOR U13642 ( .A(p_input[165]), .B(n13682), .Z(n13278) );
  AND U13643 ( .A(n530), .B(n13683), .Z(n13682) );
  XOR U13644 ( .A(p_input[181]), .B(p_input[165]), .Z(n13683) );
  XNOR U13645 ( .A(n13275), .B(n13678), .Z(n13680) );
  XOR U13646 ( .A(n13684), .B(n13685), .Z(n13275) );
  AND U13647 ( .A(n527), .B(n13686), .Z(n13685) );
  XOR U13648 ( .A(p_input[149]), .B(p_input[133]), .Z(n13686) );
  XOR U13649 ( .A(n13687), .B(n13688), .Z(n13678) );
  AND U13650 ( .A(n13689), .B(n13690), .Z(n13688) );
  XOR U13651 ( .A(n13687), .B(n13290), .Z(n13690) );
  XNOR U13652 ( .A(p_input[164]), .B(n13691), .Z(n13290) );
  AND U13653 ( .A(n530), .B(n13692), .Z(n13691) );
  XOR U13654 ( .A(p_input[180]), .B(p_input[164]), .Z(n13692) );
  XNOR U13655 ( .A(n13287), .B(n13687), .Z(n13689) );
  XOR U13656 ( .A(n13693), .B(n13694), .Z(n13287) );
  AND U13657 ( .A(n527), .B(n13695), .Z(n13694) );
  XOR U13658 ( .A(p_input[148]), .B(p_input[132]), .Z(n13695) );
  XOR U13659 ( .A(n13696), .B(n13697), .Z(n13687) );
  AND U13660 ( .A(n13698), .B(n13699), .Z(n13697) );
  XOR U13661 ( .A(n13696), .B(n13302), .Z(n13699) );
  XNOR U13662 ( .A(p_input[163]), .B(n13700), .Z(n13302) );
  AND U13663 ( .A(n530), .B(n13701), .Z(n13700) );
  XOR U13664 ( .A(p_input[179]), .B(p_input[163]), .Z(n13701) );
  XNOR U13665 ( .A(n13299), .B(n13696), .Z(n13698) );
  XOR U13666 ( .A(n13702), .B(n13703), .Z(n13299) );
  AND U13667 ( .A(n527), .B(n13704), .Z(n13703) );
  XOR U13668 ( .A(p_input[147]), .B(p_input[131]), .Z(n13704) );
  XOR U13669 ( .A(n13705), .B(n13706), .Z(n13696) );
  AND U13670 ( .A(n13707), .B(n13708), .Z(n13706) );
  XOR U13671 ( .A(n13314), .B(n13705), .Z(n13708) );
  XNOR U13672 ( .A(p_input[162]), .B(n13709), .Z(n13314) );
  AND U13673 ( .A(n530), .B(n13710), .Z(n13709) );
  XOR U13674 ( .A(p_input[178]), .B(p_input[162]), .Z(n13710) );
  XNOR U13675 ( .A(n13705), .B(n13311), .Z(n13707) );
  XOR U13676 ( .A(n13711), .B(n13712), .Z(n13311) );
  AND U13677 ( .A(n527), .B(n13713), .Z(n13712) );
  XOR U13678 ( .A(p_input[146]), .B(p_input[130]), .Z(n13713) );
  XOR U13679 ( .A(n13714), .B(n13715), .Z(n13705) );
  AND U13680 ( .A(n13716), .B(n13717), .Z(n13715) );
  XNOR U13681 ( .A(n13718), .B(n13327), .Z(n13717) );
  XNOR U13682 ( .A(p_input[161]), .B(n13719), .Z(n13327) );
  AND U13683 ( .A(n530), .B(n13720), .Z(n13719) );
  XNOR U13684 ( .A(p_input[177]), .B(n13721), .Z(n13720) );
  IV U13685 ( .A(p_input[161]), .Z(n13721) );
  XNOR U13686 ( .A(n13324), .B(n13714), .Z(n13716) );
  XNOR U13687 ( .A(p_input[129]), .B(n13722), .Z(n13324) );
  AND U13688 ( .A(n527), .B(n13723), .Z(n13722) );
  XOR U13689 ( .A(p_input[145]), .B(p_input[129]), .Z(n13723) );
  IV U13690 ( .A(n13718), .Z(n13714) );
  AND U13691 ( .A(n13589), .B(n13592), .Z(n13718) );
  XOR U13692 ( .A(p_input[160]), .B(n13724), .Z(n13592) );
  AND U13693 ( .A(n530), .B(n13725), .Z(n13724) );
  XOR U13694 ( .A(p_input[176]), .B(p_input[160]), .Z(n13725) );
  XOR U13695 ( .A(n13726), .B(n13727), .Z(n530) );
  AND U13696 ( .A(n13728), .B(n13729), .Z(n13727) );
  XNOR U13697 ( .A(p_input[191]), .B(n13726), .Z(n13729) );
  XOR U13698 ( .A(n13726), .B(p_input[175]), .Z(n13728) );
  XOR U13699 ( .A(n13730), .B(n13731), .Z(n13726) );
  AND U13700 ( .A(n13732), .B(n13733), .Z(n13731) );
  XNOR U13701 ( .A(p_input[190]), .B(n13730), .Z(n13733) );
  XOR U13702 ( .A(n13730), .B(p_input[174]), .Z(n13732) );
  XOR U13703 ( .A(n13734), .B(n13735), .Z(n13730) );
  AND U13704 ( .A(n13736), .B(n13737), .Z(n13735) );
  XNOR U13705 ( .A(p_input[189]), .B(n13734), .Z(n13737) );
  XOR U13706 ( .A(n13734), .B(p_input[173]), .Z(n13736) );
  XOR U13707 ( .A(n13738), .B(n13739), .Z(n13734) );
  AND U13708 ( .A(n13740), .B(n13741), .Z(n13739) );
  XNOR U13709 ( .A(p_input[188]), .B(n13738), .Z(n13741) );
  XOR U13710 ( .A(n13738), .B(p_input[172]), .Z(n13740) );
  XOR U13711 ( .A(n13742), .B(n13743), .Z(n13738) );
  AND U13712 ( .A(n13744), .B(n13745), .Z(n13743) );
  XNOR U13713 ( .A(p_input[187]), .B(n13742), .Z(n13745) );
  XOR U13714 ( .A(n13742), .B(p_input[171]), .Z(n13744) );
  XOR U13715 ( .A(n13746), .B(n13747), .Z(n13742) );
  AND U13716 ( .A(n13748), .B(n13749), .Z(n13747) );
  XNOR U13717 ( .A(p_input[186]), .B(n13746), .Z(n13749) );
  XOR U13718 ( .A(n13746), .B(p_input[170]), .Z(n13748) );
  XOR U13719 ( .A(n13750), .B(n13751), .Z(n13746) );
  AND U13720 ( .A(n13752), .B(n13753), .Z(n13751) );
  XNOR U13721 ( .A(p_input[185]), .B(n13750), .Z(n13753) );
  XOR U13722 ( .A(n13750), .B(p_input[169]), .Z(n13752) );
  XOR U13723 ( .A(n13754), .B(n13755), .Z(n13750) );
  AND U13724 ( .A(n13756), .B(n13757), .Z(n13755) );
  XNOR U13725 ( .A(p_input[184]), .B(n13754), .Z(n13757) );
  XOR U13726 ( .A(n13754), .B(p_input[168]), .Z(n13756) );
  XOR U13727 ( .A(n13758), .B(n13759), .Z(n13754) );
  AND U13728 ( .A(n13760), .B(n13761), .Z(n13759) );
  XNOR U13729 ( .A(p_input[183]), .B(n13758), .Z(n13761) );
  XOR U13730 ( .A(n13758), .B(p_input[167]), .Z(n13760) );
  XOR U13731 ( .A(n13762), .B(n13763), .Z(n13758) );
  AND U13732 ( .A(n13764), .B(n13765), .Z(n13763) );
  XNOR U13733 ( .A(p_input[182]), .B(n13762), .Z(n13765) );
  XOR U13734 ( .A(n13762), .B(p_input[166]), .Z(n13764) );
  XOR U13735 ( .A(n13766), .B(n13767), .Z(n13762) );
  AND U13736 ( .A(n13768), .B(n13769), .Z(n13767) );
  XNOR U13737 ( .A(p_input[181]), .B(n13766), .Z(n13769) );
  XOR U13738 ( .A(n13766), .B(p_input[165]), .Z(n13768) );
  XOR U13739 ( .A(n13770), .B(n13771), .Z(n13766) );
  AND U13740 ( .A(n13772), .B(n13773), .Z(n13771) );
  XNOR U13741 ( .A(p_input[180]), .B(n13770), .Z(n13773) );
  XOR U13742 ( .A(n13770), .B(p_input[164]), .Z(n13772) );
  XOR U13743 ( .A(n13774), .B(n13775), .Z(n13770) );
  AND U13744 ( .A(n13776), .B(n13777), .Z(n13775) );
  XNOR U13745 ( .A(p_input[179]), .B(n13774), .Z(n13777) );
  XOR U13746 ( .A(n13774), .B(p_input[163]), .Z(n13776) );
  XOR U13747 ( .A(n13778), .B(n13779), .Z(n13774) );
  AND U13748 ( .A(n13780), .B(n13781), .Z(n13779) );
  XNOR U13749 ( .A(p_input[178]), .B(n13778), .Z(n13781) );
  XOR U13750 ( .A(n13778), .B(p_input[162]), .Z(n13780) );
  XNOR U13751 ( .A(n13782), .B(n13783), .Z(n13778) );
  AND U13752 ( .A(n13784), .B(n13785), .Z(n13783) );
  XOR U13753 ( .A(p_input[177]), .B(n13782), .Z(n13785) );
  XNOR U13754 ( .A(p_input[161]), .B(n13782), .Z(n13784) );
  AND U13755 ( .A(p_input[176]), .B(n13786), .Z(n13782) );
  IV U13756 ( .A(p_input[160]), .Z(n13786) );
  XNOR U13757 ( .A(p_input[128]), .B(n13787), .Z(n13589) );
  AND U13758 ( .A(n527), .B(n13788), .Z(n13787) );
  XOR U13759 ( .A(p_input[144]), .B(p_input[128]), .Z(n13788) );
  XOR U13760 ( .A(n13789), .B(n13790), .Z(n527) );
  AND U13761 ( .A(n13791), .B(n13792), .Z(n13790) );
  XNOR U13762 ( .A(p_input[159]), .B(n13789), .Z(n13792) );
  XOR U13763 ( .A(n13789), .B(p_input[143]), .Z(n13791) );
  XOR U13764 ( .A(n13793), .B(n13794), .Z(n13789) );
  AND U13765 ( .A(n13795), .B(n13796), .Z(n13794) );
  XNOR U13766 ( .A(p_input[158]), .B(n13793), .Z(n13796) );
  XNOR U13767 ( .A(n13793), .B(n13603), .Z(n13795) );
  IV U13768 ( .A(p_input[142]), .Z(n13603) );
  XOR U13769 ( .A(n13797), .B(n13798), .Z(n13793) );
  AND U13770 ( .A(n13799), .B(n13800), .Z(n13798) );
  XNOR U13771 ( .A(p_input[157]), .B(n13797), .Z(n13800) );
  XNOR U13772 ( .A(n13797), .B(n13612), .Z(n13799) );
  IV U13773 ( .A(p_input[141]), .Z(n13612) );
  XOR U13774 ( .A(n13801), .B(n13802), .Z(n13797) );
  AND U13775 ( .A(n13803), .B(n13804), .Z(n13802) );
  XNOR U13776 ( .A(p_input[156]), .B(n13801), .Z(n13804) );
  XNOR U13777 ( .A(n13801), .B(n13621), .Z(n13803) );
  IV U13778 ( .A(p_input[140]), .Z(n13621) );
  XOR U13779 ( .A(n13805), .B(n13806), .Z(n13801) );
  AND U13780 ( .A(n13807), .B(n13808), .Z(n13806) );
  XNOR U13781 ( .A(p_input[155]), .B(n13805), .Z(n13808) );
  XNOR U13782 ( .A(n13805), .B(n13630), .Z(n13807) );
  IV U13783 ( .A(p_input[139]), .Z(n13630) );
  XOR U13784 ( .A(n13809), .B(n13810), .Z(n13805) );
  AND U13785 ( .A(n13811), .B(n13812), .Z(n13810) );
  XNOR U13786 ( .A(p_input[154]), .B(n13809), .Z(n13812) );
  XNOR U13787 ( .A(n13809), .B(n13639), .Z(n13811) );
  IV U13788 ( .A(p_input[138]), .Z(n13639) );
  XOR U13789 ( .A(n13813), .B(n13814), .Z(n13809) );
  AND U13790 ( .A(n13815), .B(n13816), .Z(n13814) );
  XNOR U13791 ( .A(p_input[153]), .B(n13813), .Z(n13816) );
  XNOR U13792 ( .A(n13813), .B(n13648), .Z(n13815) );
  IV U13793 ( .A(p_input[137]), .Z(n13648) );
  XOR U13794 ( .A(n13817), .B(n13818), .Z(n13813) );
  AND U13795 ( .A(n13819), .B(n13820), .Z(n13818) );
  XNOR U13796 ( .A(p_input[152]), .B(n13817), .Z(n13820) );
  XNOR U13797 ( .A(n13817), .B(n13657), .Z(n13819) );
  IV U13798 ( .A(p_input[136]), .Z(n13657) );
  XOR U13799 ( .A(n13821), .B(n13822), .Z(n13817) );
  AND U13800 ( .A(n13823), .B(n13824), .Z(n13822) );
  XNOR U13801 ( .A(p_input[151]), .B(n13821), .Z(n13824) );
  XNOR U13802 ( .A(n13821), .B(n13666), .Z(n13823) );
  IV U13803 ( .A(p_input[135]), .Z(n13666) );
  XOR U13804 ( .A(n13825), .B(n13826), .Z(n13821) );
  AND U13805 ( .A(n13827), .B(n13828), .Z(n13826) );
  XNOR U13806 ( .A(p_input[150]), .B(n13825), .Z(n13828) );
  XNOR U13807 ( .A(n13825), .B(n13675), .Z(n13827) );
  IV U13808 ( .A(p_input[134]), .Z(n13675) );
  XOR U13809 ( .A(n13829), .B(n13830), .Z(n13825) );
  AND U13810 ( .A(n13831), .B(n13832), .Z(n13830) );
  XNOR U13811 ( .A(p_input[149]), .B(n13829), .Z(n13832) );
  XNOR U13812 ( .A(n13829), .B(n13684), .Z(n13831) );
  IV U13813 ( .A(p_input[133]), .Z(n13684) );
  XOR U13814 ( .A(n13833), .B(n13834), .Z(n13829) );
  AND U13815 ( .A(n13835), .B(n13836), .Z(n13834) );
  XNOR U13816 ( .A(p_input[148]), .B(n13833), .Z(n13836) );
  XNOR U13817 ( .A(n13833), .B(n13693), .Z(n13835) );
  IV U13818 ( .A(p_input[132]), .Z(n13693) );
  XOR U13819 ( .A(n13837), .B(n13838), .Z(n13833) );
  AND U13820 ( .A(n13839), .B(n13840), .Z(n13838) );
  XNOR U13821 ( .A(p_input[147]), .B(n13837), .Z(n13840) );
  XNOR U13822 ( .A(n13837), .B(n13702), .Z(n13839) );
  IV U13823 ( .A(p_input[131]), .Z(n13702) );
  XOR U13824 ( .A(n13841), .B(n13842), .Z(n13837) );
  AND U13825 ( .A(n13843), .B(n13844), .Z(n13842) );
  XNOR U13826 ( .A(p_input[146]), .B(n13841), .Z(n13844) );
  XNOR U13827 ( .A(n13841), .B(n13711), .Z(n13843) );
  IV U13828 ( .A(p_input[130]), .Z(n13711) );
  XNOR U13829 ( .A(n13845), .B(n13846), .Z(n13841) );
  AND U13830 ( .A(n13847), .B(n13848), .Z(n13846) );
  XOR U13831 ( .A(p_input[145]), .B(n13845), .Z(n13848) );
  XNOR U13832 ( .A(p_input[129]), .B(n13845), .Z(n13847) );
  AND U13833 ( .A(p_input[144]), .B(n13849), .Z(n13845) );
  IV U13834 ( .A(p_input[128]), .Z(n13849) );
  XOR U13835 ( .A(n13850), .B(n13851), .Z(n12965) );
  AND U13836 ( .A(n451), .B(n13852), .Z(n13851) );
  XNOR U13837 ( .A(n13853), .B(n13850), .Z(n13852) );
  XOR U13838 ( .A(n13854), .B(n13855), .Z(n451) );
  AND U13839 ( .A(n13856), .B(n13857), .Z(n13855) );
  XNOR U13840 ( .A(n12977), .B(n13854), .Z(n13857) );
  AND U13841 ( .A(n13858), .B(n13859), .Z(n12977) );
  XOR U13842 ( .A(n13854), .B(n12976), .Z(n13856) );
  AND U13843 ( .A(n13860), .B(n13861), .Z(n12976) );
  XOR U13844 ( .A(n13862), .B(n13863), .Z(n13854) );
  AND U13845 ( .A(n13864), .B(n13865), .Z(n13863) );
  XOR U13846 ( .A(n13862), .B(n12989), .Z(n13865) );
  XOR U13847 ( .A(n13866), .B(n13867), .Z(n12989) );
  AND U13848 ( .A(n330), .B(n13868), .Z(n13867) );
  XOR U13849 ( .A(n13869), .B(n13866), .Z(n13868) );
  XNOR U13850 ( .A(n12986), .B(n13862), .Z(n13864) );
  XOR U13851 ( .A(n13870), .B(n13871), .Z(n12986) );
  AND U13852 ( .A(n327), .B(n13872), .Z(n13871) );
  XOR U13853 ( .A(n13873), .B(n13870), .Z(n13872) );
  XOR U13854 ( .A(n13874), .B(n13875), .Z(n13862) );
  AND U13855 ( .A(n13876), .B(n13877), .Z(n13875) );
  XOR U13856 ( .A(n13874), .B(n13001), .Z(n13877) );
  XOR U13857 ( .A(n13878), .B(n13879), .Z(n13001) );
  AND U13858 ( .A(n330), .B(n13880), .Z(n13879) );
  XOR U13859 ( .A(n13881), .B(n13878), .Z(n13880) );
  XNOR U13860 ( .A(n12998), .B(n13874), .Z(n13876) );
  XOR U13861 ( .A(n13882), .B(n13883), .Z(n12998) );
  AND U13862 ( .A(n327), .B(n13884), .Z(n13883) );
  XOR U13863 ( .A(n13885), .B(n13882), .Z(n13884) );
  XOR U13864 ( .A(n13886), .B(n13887), .Z(n13874) );
  AND U13865 ( .A(n13888), .B(n13889), .Z(n13887) );
  XOR U13866 ( .A(n13886), .B(n13013), .Z(n13889) );
  XOR U13867 ( .A(n13890), .B(n13891), .Z(n13013) );
  AND U13868 ( .A(n330), .B(n13892), .Z(n13891) );
  XOR U13869 ( .A(n13893), .B(n13890), .Z(n13892) );
  XNOR U13870 ( .A(n13010), .B(n13886), .Z(n13888) );
  XOR U13871 ( .A(n13894), .B(n13895), .Z(n13010) );
  AND U13872 ( .A(n327), .B(n13896), .Z(n13895) );
  XOR U13873 ( .A(n13897), .B(n13894), .Z(n13896) );
  XOR U13874 ( .A(n13898), .B(n13899), .Z(n13886) );
  AND U13875 ( .A(n13900), .B(n13901), .Z(n13899) );
  XOR U13876 ( .A(n13898), .B(n13025), .Z(n13901) );
  XOR U13877 ( .A(n13902), .B(n13903), .Z(n13025) );
  AND U13878 ( .A(n330), .B(n13904), .Z(n13903) );
  XOR U13879 ( .A(n13905), .B(n13902), .Z(n13904) );
  XNOR U13880 ( .A(n13022), .B(n13898), .Z(n13900) );
  XOR U13881 ( .A(n13906), .B(n13907), .Z(n13022) );
  AND U13882 ( .A(n327), .B(n13908), .Z(n13907) );
  XOR U13883 ( .A(n13909), .B(n13906), .Z(n13908) );
  XOR U13884 ( .A(n13910), .B(n13911), .Z(n13898) );
  AND U13885 ( .A(n13912), .B(n13913), .Z(n13911) );
  XOR U13886 ( .A(n13910), .B(n13037), .Z(n13913) );
  XOR U13887 ( .A(n13914), .B(n13915), .Z(n13037) );
  AND U13888 ( .A(n330), .B(n13916), .Z(n13915) );
  XOR U13889 ( .A(n13917), .B(n13914), .Z(n13916) );
  XNOR U13890 ( .A(n13034), .B(n13910), .Z(n13912) );
  XOR U13891 ( .A(n13918), .B(n13919), .Z(n13034) );
  AND U13892 ( .A(n327), .B(n13920), .Z(n13919) );
  XOR U13893 ( .A(n13921), .B(n13918), .Z(n13920) );
  XOR U13894 ( .A(n13922), .B(n13923), .Z(n13910) );
  AND U13895 ( .A(n13924), .B(n13925), .Z(n13923) );
  XOR U13896 ( .A(n13922), .B(n13049), .Z(n13925) );
  XOR U13897 ( .A(n13926), .B(n13927), .Z(n13049) );
  AND U13898 ( .A(n330), .B(n13928), .Z(n13927) );
  XOR U13899 ( .A(n13929), .B(n13926), .Z(n13928) );
  XNOR U13900 ( .A(n13046), .B(n13922), .Z(n13924) );
  XOR U13901 ( .A(n13930), .B(n13931), .Z(n13046) );
  AND U13902 ( .A(n327), .B(n13932), .Z(n13931) );
  XOR U13903 ( .A(n13933), .B(n13930), .Z(n13932) );
  XOR U13904 ( .A(n13934), .B(n13935), .Z(n13922) );
  AND U13905 ( .A(n13936), .B(n13937), .Z(n13935) );
  XOR U13906 ( .A(n13934), .B(n13061), .Z(n13937) );
  XOR U13907 ( .A(n13938), .B(n13939), .Z(n13061) );
  AND U13908 ( .A(n330), .B(n13940), .Z(n13939) );
  XOR U13909 ( .A(n13941), .B(n13938), .Z(n13940) );
  XNOR U13910 ( .A(n13058), .B(n13934), .Z(n13936) );
  XOR U13911 ( .A(n13942), .B(n13943), .Z(n13058) );
  AND U13912 ( .A(n327), .B(n13944), .Z(n13943) );
  XOR U13913 ( .A(n13945), .B(n13942), .Z(n13944) );
  XOR U13914 ( .A(n13946), .B(n13947), .Z(n13934) );
  AND U13915 ( .A(n13948), .B(n13949), .Z(n13947) );
  XOR U13916 ( .A(n13946), .B(n13073), .Z(n13949) );
  XOR U13917 ( .A(n13950), .B(n13951), .Z(n13073) );
  AND U13918 ( .A(n330), .B(n13952), .Z(n13951) );
  XOR U13919 ( .A(n13953), .B(n13950), .Z(n13952) );
  XNOR U13920 ( .A(n13070), .B(n13946), .Z(n13948) );
  XOR U13921 ( .A(n13954), .B(n13955), .Z(n13070) );
  AND U13922 ( .A(n327), .B(n13956), .Z(n13955) );
  XOR U13923 ( .A(n13957), .B(n13954), .Z(n13956) );
  XOR U13924 ( .A(n13958), .B(n13959), .Z(n13946) );
  AND U13925 ( .A(n13960), .B(n13961), .Z(n13959) );
  XOR U13926 ( .A(n13958), .B(n13085), .Z(n13961) );
  XOR U13927 ( .A(n13962), .B(n13963), .Z(n13085) );
  AND U13928 ( .A(n330), .B(n13964), .Z(n13963) );
  XOR U13929 ( .A(n13965), .B(n13962), .Z(n13964) );
  XNOR U13930 ( .A(n13082), .B(n13958), .Z(n13960) );
  XOR U13931 ( .A(n13966), .B(n13967), .Z(n13082) );
  AND U13932 ( .A(n327), .B(n13968), .Z(n13967) );
  XOR U13933 ( .A(n13969), .B(n13966), .Z(n13968) );
  XOR U13934 ( .A(n13970), .B(n13971), .Z(n13958) );
  AND U13935 ( .A(n13972), .B(n13973), .Z(n13971) );
  XOR U13936 ( .A(n13970), .B(n13097), .Z(n13973) );
  XOR U13937 ( .A(n13974), .B(n13975), .Z(n13097) );
  AND U13938 ( .A(n330), .B(n13976), .Z(n13975) );
  XOR U13939 ( .A(n13977), .B(n13974), .Z(n13976) );
  XNOR U13940 ( .A(n13094), .B(n13970), .Z(n13972) );
  XOR U13941 ( .A(n13978), .B(n13979), .Z(n13094) );
  AND U13942 ( .A(n327), .B(n13980), .Z(n13979) );
  XOR U13943 ( .A(n13981), .B(n13978), .Z(n13980) );
  XOR U13944 ( .A(n13982), .B(n13983), .Z(n13970) );
  AND U13945 ( .A(n13984), .B(n13985), .Z(n13983) );
  XOR U13946 ( .A(n13982), .B(n13109), .Z(n13985) );
  XOR U13947 ( .A(n13986), .B(n13987), .Z(n13109) );
  AND U13948 ( .A(n330), .B(n13988), .Z(n13987) );
  XOR U13949 ( .A(n13989), .B(n13986), .Z(n13988) );
  XNOR U13950 ( .A(n13106), .B(n13982), .Z(n13984) );
  XOR U13951 ( .A(n13990), .B(n13991), .Z(n13106) );
  AND U13952 ( .A(n327), .B(n13992), .Z(n13991) );
  XOR U13953 ( .A(n13993), .B(n13990), .Z(n13992) );
  XOR U13954 ( .A(n13994), .B(n13995), .Z(n13982) );
  AND U13955 ( .A(n13996), .B(n13997), .Z(n13995) );
  XOR U13956 ( .A(n13994), .B(n13121), .Z(n13997) );
  XOR U13957 ( .A(n13998), .B(n13999), .Z(n13121) );
  AND U13958 ( .A(n330), .B(n14000), .Z(n13999) );
  XOR U13959 ( .A(n14001), .B(n13998), .Z(n14000) );
  XNOR U13960 ( .A(n13118), .B(n13994), .Z(n13996) );
  XOR U13961 ( .A(n14002), .B(n14003), .Z(n13118) );
  AND U13962 ( .A(n327), .B(n14004), .Z(n14003) );
  XOR U13963 ( .A(n14005), .B(n14002), .Z(n14004) );
  XOR U13964 ( .A(n14006), .B(n14007), .Z(n13994) );
  AND U13965 ( .A(n14008), .B(n14009), .Z(n14007) );
  XOR U13966 ( .A(n13133), .B(n14006), .Z(n14009) );
  XOR U13967 ( .A(n14010), .B(n14011), .Z(n13133) );
  AND U13968 ( .A(n330), .B(n14012), .Z(n14011) );
  XOR U13969 ( .A(n14010), .B(n14013), .Z(n14012) );
  XNOR U13970 ( .A(n14006), .B(n13130), .Z(n14008) );
  XOR U13971 ( .A(n14014), .B(n14015), .Z(n13130) );
  AND U13972 ( .A(n327), .B(n14016), .Z(n14015) );
  XOR U13973 ( .A(n14014), .B(n14017), .Z(n14016) );
  XOR U13974 ( .A(n14018), .B(n14019), .Z(n14006) );
  AND U13975 ( .A(n14020), .B(n14021), .Z(n14019) );
  XNOR U13976 ( .A(n14022), .B(n13146), .Z(n14021) );
  XOR U13977 ( .A(n14023), .B(n14024), .Z(n13146) );
  AND U13978 ( .A(n330), .B(n14025), .Z(n14024) );
  XOR U13979 ( .A(n14026), .B(n14023), .Z(n14025) );
  XNOR U13980 ( .A(n13143), .B(n14018), .Z(n14020) );
  XOR U13981 ( .A(n14027), .B(n14028), .Z(n13143) );
  AND U13982 ( .A(n327), .B(n14029), .Z(n14028) );
  XOR U13983 ( .A(n14030), .B(n14027), .Z(n14029) );
  IV U13984 ( .A(n14022), .Z(n14018) );
  AND U13985 ( .A(n13850), .B(n13853), .Z(n14022) );
  XNOR U13986 ( .A(n14031), .B(n14032), .Z(n13853) );
  AND U13987 ( .A(n330), .B(n14033), .Z(n14032) );
  XNOR U13988 ( .A(n14034), .B(n14031), .Z(n14033) );
  XOR U13989 ( .A(n14035), .B(n14036), .Z(n330) );
  AND U13990 ( .A(n14037), .B(n14038), .Z(n14036) );
  XNOR U13991 ( .A(n13858), .B(n14035), .Z(n14038) );
  AND U13992 ( .A(p_input[127]), .B(p_input[111]), .Z(n13858) );
  XOR U13993 ( .A(n14035), .B(n13859), .Z(n14037) );
  AND U13994 ( .A(p_input[95]), .B(p_input[79]), .Z(n13859) );
  XOR U13995 ( .A(n14039), .B(n14040), .Z(n14035) );
  AND U13996 ( .A(n14041), .B(n14042), .Z(n14040) );
  XOR U13997 ( .A(n14039), .B(n13869), .Z(n14042) );
  XNOR U13998 ( .A(p_input[110]), .B(n14043), .Z(n13869) );
  AND U13999 ( .A(n550), .B(n14044), .Z(n14043) );
  XOR U14000 ( .A(p_input[126]), .B(p_input[110]), .Z(n14044) );
  XNOR U14001 ( .A(n13866), .B(n14039), .Z(n14041) );
  XOR U14002 ( .A(n14045), .B(n14046), .Z(n13866) );
  AND U14003 ( .A(n548), .B(n14047), .Z(n14046) );
  XOR U14004 ( .A(p_input[94]), .B(p_input[78]), .Z(n14047) );
  XOR U14005 ( .A(n14048), .B(n14049), .Z(n14039) );
  AND U14006 ( .A(n14050), .B(n14051), .Z(n14049) );
  XOR U14007 ( .A(n14048), .B(n13881), .Z(n14051) );
  XNOR U14008 ( .A(p_input[109]), .B(n14052), .Z(n13881) );
  AND U14009 ( .A(n550), .B(n14053), .Z(n14052) );
  XOR U14010 ( .A(p_input[125]), .B(p_input[109]), .Z(n14053) );
  XNOR U14011 ( .A(n13878), .B(n14048), .Z(n14050) );
  XOR U14012 ( .A(n14054), .B(n14055), .Z(n13878) );
  AND U14013 ( .A(n548), .B(n14056), .Z(n14055) );
  XOR U14014 ( .A(p_input[93]), .B(p_input[77]), .Z(n14056) );
  XOR U14015 ( .A(n14057), .B(n14058), .Z(n14048) );
  AND U14016 ( .A(n14059), .B(n14060), .Z(n14058) );
  XOR U14017 ( .A(n14057), .B(n13893), .Z(n14060) );
  XNOR U14018 ( .A(p_input[108]), .B(n14061), .Z(n13893) );
  AND U14019 ( .A(n550), .B(n14062), .Z(n14061) );
  XOR U14020 ( .A(p_input[124]), .B(p_input[108]), .Z(n14062) );
  XNOR U14021 ( .A(n13890), .B(n14057), .Z(n14059) );
  XOR U14022 ( .A(n14063), .B(n14064), .Z(n13890) );
  AND U14023 ( .A(n548), .B(n14065), .Z(n14064) );
  XOR U14024 ( .A(p_input[92]), .B(p_input[76]), .Z(n14065) );
  XOR U14025 ( .A(n14066), .B(n14067), .Z(n14057) );
  AND U14026 ( .A(n14068), .B(n14069), .Z(n14067) );
  XOR U14027 ( .A(n14066), .B(n13905), .Z(n14069) );
  XNOR U14028 ( .A(p_input[107]), .B(n14070), .Z(n13905) );
  AND U14029 ( .A(n550), .B(n14071), .Z(n14070) );
  XOR U14030 ( .A(p_input[123]), .B(p_input[107]), .Z(n14071) );
  XNOR U14031 ( .A(n13902), .B(n14066), .Z(n14068) );
  XOR U14032 ( .A(n14072), .B(n14073), .Z(n13902) );
  AND U14033 ( .A(n548), .B(n14074), .Z(n14073) );
  XOR U14034 ( .A(p_input[91]), .B(p_input[75]), .Z(n14074) );
  XOR U14035 ( .A(n14075), .B(n14076), .Z(n14066) );
  AND U14036 ( .A(n14077), .B(n14078), .Z(n14076) );
  XOR U14037 ( .A(n14075), .B(n13917), .Z(n14078) );
  XNOR U14038 ( .A(p_input[106]), .B(n14079), .Z(n13917) );
  AND U14039 ( .A(n550), .B(n14080), .Z(n14079) );
  XOR U14040 ( .A(p_input[122]), .B(p_input[106]), .Z(n14080) );
  XNOR U14041 ( .A(n13914), .B(n14075), .Z(n14077) );
  XOR U14042 ( .A(n14081), .B(n14082), .Z(n13914) );
  AND U14043 ( .A(n548), .B(n14083), .Z(n14082) );
  XOR U14044 ( .A(p_input[90]), .B(p_input[74]), .Z(n14083) );
  XOR U14045 ( .A(n14084), .B(n14085), .Z(n14075) );
  AND U14046 ( .A(n14086), .B(n14087), .Z(n14085) );
  XOR U14047 ( .A(n14084), .B(n13929), .Z(n14087) );
  XNOR U14048 ( .A(p_input[105]), .B(n14088), .Z(n13929) );
  AND U14049 ( .A(n550), .B(n14089), .Z(n14088) );
  XOR U14050 ( .A(p_input[121]), .B(p_input[105]), .Z(n14089) );
  XNOR U14051 ( .A(n13926), .B(n14084), .Z(n14086) );
  XOR U14052 ( .A(n14090), .B(n14091), .Z(n13926) );
  AND U14053 ( .A(n548), .B(n14092), .Z(n14091) );
  XOR U14054 ( .A(p_input[89]), .B(p_input[73]), .Z(n14092) );
  XOR U14055 ( .A(n14093), .B(n14094), .Z(n14084) );
  AND U14056 ( .A(n14095), .B(n14096), .Z(n14094) );
  XOR U14057 ( .A(n14093), .B(n13941), .Z(n14096) );
  XNOR U14058 ( .A(p_input[104]), .B(n14097), .Z(n13941) );
  AND U14059 ( .A(n550), .B(n14098), .Z(n14097) );
  XOR U14060 ( .A(p_input[120]), .B(p_input[104]), .Z(n14098) );
  XNOR U14061 ( .A(n13938), .B(n14093), .Z(n14095) );
  XOR U14062 ( .A(n14099), .B(n14100), .Z(n13938) );
  AND U14063 ( .A(n548), .B(n14101), .Z(n14100) );
  XOR U14064 ( .A(p_input[88]), .B(p_input[72]), .Z(n14101) );
  XOR U14065 ( .A(n14102), .B(n14103), .Z(n14093) );
  AND U14066 ( .A(n14104), .B(n14105), .Z(n14103) );
  XOR U14067 ( .A(n14102), .B(n13953), .Z(n14105) );
  XNOR U14068 ( .A(p_input[103]), .B(n14106), .Z(n13953) );
  AND U14069 ( .A(n550), .B(n14107), .Z(n14106) );
  XOR U14070 ( .A(p_input[119]), .B(p_input[103]), .Z(n14107) );
  XNOR U14071 ( .A(n13950), .B(n14102), .Z(n14104) );
  XOR U14072 ( .A(n14108), .B(n14109), .Z(n13950) );
  AND U14073 ( .A(n548), .B(n14110), .Z(n14109) );
  XOR U14074 ( .A(p_input[87]), .B(p_input[71]), .Z(n14110) );
  XOR U14075 ( .A(n14111), .B(n14112), .Z(n14102) );
  AND U14076 ( .A(n14113), .B(n14114), .Z(n14112) );
  XOR U14077 ( .A(n14111), .B(n13965), .Z(n14114) );
  XNOR U14078 ( .A(p_input[102]), .B(n14115), .Z(n13965) );
  AND U14079 ( .A(n550), .B(n14116), .Z(n14115) );
  XOR U14080 ( .A(p_input[118]), .B(p_input[102]), .Z(n14116) );
  XNOR U14081 ( .A(n13962), .B(n14111), .Z(n14113) );
  XOR U14082 ( .A(n14117), .B(n14118), .Z(n13962) );
  AND U14083 ( .A(n548), .B(n14119), .Z(n14118) );
  XOR U14084 ( .A(p_input[86]), .B(p_input[70]), .Z(n14119) );
  XOR U14085 ( .A(n14120), .B(n14121), .Z(n14111) );
  AND U14086 ( .A(n14122), .B(n14123), .Z(n14121) );
  XOR U14087 ( .A(n14120), .B(n13977), .Z(n14123) );
  XNOR U14088 ( .A(p_input[101]), .B(n14124), .Z(n13977) );
  AND U14089 ( .A(n550), .B(n14125), .Z(n14124) );
  XOR U14090 ( .A(p_input[117]), .B(p_input[101]), .Z(n14125) );
  XNOR U14091 ( .A(n13974), .B(n14120), .Z(n14122) );
  XOR U14092 ( .A(n14126), .B(n14127), .Z(n13974) );
  AND U14093 ( .A(n548), .B(n14128), .Z(n14127) );
  XOR U14094 ( .A(p_input[85]), .B(p_input[69]), .Z(n14128) );
  XOR U14095 ( .A(n14129), .B(n14130), .Z(n14120) );
  AND U14096 ( .A(n14131), .B(n14132), .Z(n14130) );
  XOR U14097 ( .A(n14129), .B(n13989), .Z(n14132) );
  XNOR U14098 ( .A(p_input[100]), .B(n14133), .Z(n13989) );
  AND U14099 ( .A(n550), .B(n14134), .Z(n14133) );
  XOR U14100 ( .A(p_input[116]), .B(p_input[100]), .Z(n14134) );
  XNOR U14101 ( .A(n13986), .B(n14129), .Z(n14131) );
  XOR U14102 ( .A(n14135), .B(n14136), .Z(n13986) );
  AND U14103 ( .A(n548), .B(n14137), .Z(n14136) );
  XOR U14104 ( .A(p_input[84]), .B(p_input[68]), .Z(n14137) );
  XOR U14105 ( .A(n14138), .B(n14139), .Z(n14129) );
  AND U14106 ( .A(n14140), .B(n14141), .Z(n14139) );
  XOR U14107 ( .A(n14138), .B(n14001), .Z(n14141) );
  XNOR U14108 ( .A(p_input[99]), .B(n14142), .Z(n14001) );
  AND U14109 ( .A(n550), .B(n14143), .Z(n14142) );
  XOR U14110 ( .A(p_input[99]), .B(p_input[115]), .Z(n14143) );
  XNOR U14111 ( .A(n13998), .B(n14138), .Z(n14140) );
  XOR U14112 ( .A(n14144), .B(n14145), .Z(n13998) );
  AND U14113 ( .A(n548), .B(n14146), .Z(n14145) );
  XOR U14114 ( .A(p_input[83]), .B(p_input[67]), .Z(n14146) );
  XOR U14115 ( .A(n14147), .B(n14148), .Z(n14138) );
  AND U14116 ( .A(n14149), .B(n14150), .Z(n14148) );
  XOR U14117 ( .A(n14013), .B(n14147), .Z(n14150) );
  XNOR U14118 ( .A(p_input[98]), .B(n14151), .Z(n14013) );
  AND U14119 ( .A(n550), .B(n14152), .Z(n14151) );
  XOR U14120 ( .A(p_input[98]), .B(p_input[114]), .Z(n14152) );
  XNOR U14121 ( .A(n14147), .B(n14010), .Z(n14149) );
  XOR U14122 ( .A(n14153), .B(n14154), .Z(n14010) );
  AND U14123 ( .A(n548), .B(n14155), .Z(n14154) );
  XOR U14124 ( .A(p_input[82]), .B(p_input[66]), .Z(n14155) );
  XOR U14125 ( .A(n14156), .B(n14157), .Z(n14147) );
  AND U14126 ( .A(n14158), .B(n14159), .Z(n14157) );
  XNOR U14127 ( .A(n14160), .B(n14026), .Z(n14159) );
  XNOR U14128 ( .A(p_input[97]), .B(n14161), .Z(n14026) );
  AND U14129 ( .A(n550), .B(n14162), .Z(n14161) );
  XNOR U14130 ( .A(n14163), .B(p_input[113]), .Z(n14162) );
  IV U14131 ( .A(p_input[97]), .Z(n14163) );
  XNOR U14132 ( .A(n14023), .B(n14156), .Z(n14158) );
  XNOR U14133 ( .A(p_input[65]), .B(n14164), .Z(n14023) );
  AND U14134 ( .A(n548), .B(n14165), .Z(n14164) );
  XOR U14135 ( .A(p_input[81]), .B(p_input[65]), .Z(n14165) );
  IV U14136 ( .A(n14160), .Z(n14156) );
  AND U14137 ( .A(n14031), .B(n14034), .Z(n14160) );
  XOR U14138 ( .A(p_input[96]), .B(n14166), .Z(n14034) );
  AND U14139 ( .A(n550), .B(n14167), .Z(n14166) );
  XOR U14140 ( .A(p_input[96]), .B(p_input[112]), .Z(n14167) );
  XOR U14141 ( .A(n14168), .B(n14169), .Z(n550) );
  AND U14142 ( .A(n14170), .B(n14171), .Z(n14169) );
  XNOR U14143 ( .A(p_input[127]), .B(n14168), .Z(n14171) );
  XOR U14144 ( .A(n14168), .B(p_input[111]), .Z(n14170) );
  XOR U14145 ( .A(n14172), .B(n14173), .Z(n14168) );
  AND U14146 ( .A(n14174), .B(n14175), .Z(n14173) );
  XNOR U14147 ( .A(p_input[126]), .B(n14172), .Z(n14175) );
  XOR U14148 ( .A(n14172), .B(p_input[110]), .Z(n14174) );
  XOR U14149 ( .A(n14176), .B(n14177), .Z(n14172) );
  AND U14150 ( .A(n14178), .B(n14179), .Z(n14177) );
  XNOR U14151 ( .A(p_input[125]), .B(n14176), .Z(n14179) );
  XOR U14152 ( .A(n14176), .B(p_input[109]), .Z(n14178) );
  XOR U14153 ( .A(n14180), .B(n14181), .Z(n14176) );
  AND U14154 ( .A(n14182), .B(n14183), .Z(n14181) );
  XNOR U14155 ( .A(p_input[124]), .B(n14180), .Z(n14183) );
  XOR U14156 ( .A(n14180), .B(p_input[108]), .Z(n14182) );
  XOR U14157 ( .A(n14184), .B(n14185), .Z(n14180) );
  AND U14158 ( .A(n14186), .B(n14187), .Z(n14185) );
  XNOR U14159 ( .A(p_input[123]), .B(n14184), .Z(n14187) );
  XOR U14160 ( .A(n14184), .B(p_input[107]), .Z(n14186) );
  XOR U14161 ( .A(n14188), .B(n14189), .Z(n14184) );
  AND U14162 ( .A(n14190), .B(n14191), .Z(n14189) );
  XNOR U14163 ( .A(p_input[122]), .B(n14188), .Z(n14191) );
  XOR U14164 ( .A(n14188), .B(p_input[106]), .Z(n14190) );
  XOR U14165 ( .A(n14192), .B(n14193), .Z(n14188) );
  AND U14166 ( .A(n14194), .B(n14195), .Z(n14193) );
  XNOR U14167 ( .A(p_input[121]), .B(n14192), .Z(n14195) );
  XOR U14168 ( .A(n14192), .B(p_input[105]), .Z(n14194) );
  XOR U14169 ( .A(n14196), .B(n14197), .Z(n14192) );
  AND U14170 ( .A(n14198), .B(n14199), .Z(n14197) );
  XNOR U14171 ( .A(p_input[120]), .B(n14196), .Z(n14199) );
  XOR U14172 ( .A(n14196), .B(p_input[104]), .Z(n14198) );
  XOR U14173 ( .A(n14200), .B(n14201), .Z(n14196) );
  AND U14174 ( .A(n14202), .B(n14203), .Z(n14201) );
  XNOR U14175 ( .A(p_input[119]), .B(n14200), .Z(n14203) );
  XOR U14176 ( .A(n14200), .B(p_input[103]), .Z(n14202) );
  XOR U14177 ( .A(n14204), .B(n14205), .Z(n14200) );
  AND U14178 ( .A(n14206), .B(n14207), .Z(n14205) );
  XNOR U14179 ( .A(p_input[118]), .B(n14204), .Z(n14207) );
  XOR U14180 ( .A(n14204), .B(p_input[102]), .Z(n14206) );
  XOR U14181 ( .A(n14208), .B(n14209), .Z(n14204) );
  AND U14182 ( .A(n14210), .B(n14211), .Z(n14209) );
  XNOR U14183 ( .A(p_input[117]), .B(n14208), .Z(n14211) );
  XOR U14184 ( .A(n14208), .B(p_input[101]), .Z(n14210) );
  XOR U14185 ( .A(n14212), .B(n14213), .Z(n14208) );
  AND U14186 ( .A(n14214), .B(n14215), .Z(n14213) );
  XNOR U14187 ( .A(p_input[116]), .B(n14212), .Z(n14215) );
  XOR U14188 ( .A(n14212), .B(p_input[100]), .Z(n14214) );
  XOR U14189 ( .A(n14216), .B(n14217), .Z(n14212) );
  AND U14190 ( .A(n14218), .B(n14219), .Z(n14217) );
  XNOR U14191 ( .A(p_input[115]), .B(n14216), .Z(n14219) );
  XOR U14192 ( .A(n14216), .B(p_input[99]), .Z(n14218) );
  XOR U14193 ( .A(n14220), .B(n14221), .Z(n14216) );
  AND U14194 ( .A(n14222), .B(n14223), .Z(n14221) );
  XNOR U14195 ( .A(p_input[114]), .B(n14220), .Z(n14223) );
  XOR U14196 ( .A(n14220), .B(p_input[98]), .Z(n14222) );
  XNOR U14197 ( .A(n14224), .B(n14225), .Z(n14220) );
  AND U14198 ( .A(n14226), .B(n14227), .Z(n14225) );
  XOR U14199 ( .A(p_input[113]), .B(n14224), .Z(n14227) );
  XNOR U14200 ( .A(p_input[97]), .B(n14224), .Z(n14226) );
  AND U14201 ( .A(p_input[112]), .B(n14228), .Z(n14224) );
  IV U14202 ( .A(p_input[96]), .Z(n14228) );
  XNOR U14203 ( .A(p_input[64]), .B(n14229), .Z(n14031) );
  AND U14204 ( .A(n548), .B(n14230), .Z(n14229) );
  XOR U14205 ( .A(p_input[80]), .B(p_input[64]), .Z(n14230) );
  XOR U14206 ( .A(n14231), .B(n14232), .Z(n548) );
  AND U14207 ( .A(n14233), .B(n14234), .Z(n14232) );
  XNOR U14208 ( .A(p_input[95]), .B(n14231), .Z(n14234) );
  XOR U14209 ( .A(n14231), .B(p_input[79]), .Z(n14233) );
  XOR U14210 ( .A(n14235), .B(n14236), .Z(n14231) );
  AND U14211 ( .A(n14237), .B(n14238), .Z(n14236) );
  XNOR U14212 ( .A(p_input[94]), .B(n14235), .Z(n14238) );
  XNOR U14213 ( .A(n14235), .B(n14045), .Z(n14237) );
  IV U14214 ( .A(p_input[78]), .Z(n14045) );
  XOR U14215 ( .A(n14239), .B(n14240), .Z(n14235) );
  AND U14216 ( .A(n14241), .B(n14242), .Z(n14240) );
  XNOR U14217 ( .A(p_input[93]), .B(n14239), .Z(n14242) );
  XNOR U14218 ( .A(n14239), .B(n14054), .Z(n14241) );
  IV U14219 ( .A(p_input[77]), .Z(n14054) );
  XOR U14220 ( .A(n14243), .B(n14244), .Z(n14239) );
  AND U14221 ( .A(n14245), .B(n14246), .Z(n14244) );
  XNOR U14222 ( .A(p_input[92]), .B(n14243), .Z(n14246) );
  XNOR U14223 ( .A(n14243), .B(n14063), .Z(n14245) );
  IV U14224 ( .A(p_input[76]), .Z(n14063) );
  XOR U14225 ( .A(n14247), .B(n14248), .Z(n14243) );
  AND U14226 ( .A(n14249), .B(n14250), .Z(n14248) );
  XNOR U14227 ( .A(p_input[91]), .B(n14247), .Z(n14250) );
  XNOR U14228 ( .A(n14247), .B(n14072), .Z(n14249) );
  IV U14229 ( .A(p_input[75]), .Z(n14072) );
  XOR U14230 ( .A(n14251), .B(n14252), .Z(n14247) );
  AND U14231 ( .A(n14253), .B(n14254), .Z(n14252) );
  XNOR U14232 ( .A(p_input[90]), .B(n14251), .Z(n14254) );
  XNOR U14233 ( .A(n14251), .B(n14081), .Z(n14253) );
  IV U14234 ( .A(p_input[74]), .Z(n14081) );
  XOR U14235 ( .A(n14255), .B(n14256), .Z(n14251) );
  AND U14236 ( .A(n14257), .B(n14258), .Z(n14256) );
  XNOR U14237 ( .A(p_input[89]), .B(n14255), .Z(n14258) );
  XNOR U14238 ( .A(n14255), .B(n14090), .Z(n14257) );
  IV U14239 ( .A(p_input[73]), .Z(n14090) );
  XOR U14240 ( .A(n14259), .B(n14260), .Z(n14255) );
  AND U14241 ( .A(n14261), .B(n14262), .Z(n14260) );
  XNOR U14242 ( .A(p_input[88]), .B(n14259), .Z(n14262) );
  XNOR U14243 ( .A(n14259), .B(n14099), .Z(n14261) );
  IV U14244 ( .A(p_input[72]), .Z(n14099) );
  XOR U14245 ( .A(n14263), .B(n14264), .Z(n14259) );
  AND U14246 ( .A(n14265), .B(n14266), .Z(n14264) );
  XNOR U14247 ( .A(p_input[87]), .B(n14263), .Z(n14266) );
  XNOR U14248 ( .A(n14263), .B(n14108), .Z(n14265) );
  IV U14249 ( .A(p_input[71]), .Z(n14108) );
  XOR U14250 ( .A(n14267), .B(n14268), .Z(n14263) );
  AND U14251 ( .A(n14269), .B(n14270), .Z(n14268) );
  XNOR U14252 ( .A(p_input[86]), .B(n14267), .Z(n14270) );
  XNOR U14253 ( .A(n14267), .B(n14117), .Z(n14269) );
  IV U14254 ( .A(p_input[70]), .Z(n14117) );
  XOR U14255 ( .A(n14271), .B(n14272), .Z(n14267) );
  AND U14256 ( .A(n14273), .B(n14274), .Z(n14272) );
  XNOR U14257 ( .A(p_input[85]), .B(n14271), .Z(n14274) );
  XNOR U14258 ( .A(n14271), .B(n14126), .Z(n14273) );
  IV U14259 ( .A(p_input[69]), .Z(n14126) );
  XOR U14260 ( .A(n14275), .B(n14276), .Z(n14271) );
  AND U14261 ( .A(n14277), .B(n14278), .Z(n14276) );
  XNOR U14262 ( .A(p_input[84]), .B(n14275), .Z(n14278) );
  XNOR U14263 ( .A(n14275), .B(n14135), .Z(n14277) );
  IV U14264 ( .A(p_input[68]), .Z(n14135) );
  XOR U14265 ( .A(n14279), .B(n14280), .Z(n14275) );
  AND U14266 ( .A(n14281), .B(n14282), .Z(n14280) );
  XNOR U14267 ( .A(p_input[83]), .B(n14279), .Z(n14282) );
  XNOR U14268 ( .A(n14279), .B(n14144), .Z(n14281) );
  IV U14269 ( .A(p_input[67]), .Z(n14144) );
  XOR U14270 ( .A(n14283), .B(n14284), .Z(n14279) );
  AND U14271 ( .A(n14285), .B(n14286), .Z(n14284) );
  XNOR U14272 ( .A(p_input[82]), .B(n14283), .Z(n14286) );
  XNOR U14273 ( .A(n14283), .B(n14153), .Z(n14285) );
  IV U14274 ( .A(p_input[66]), .Z(n14153) );
  XNOR U14275 ( .A(n14287), .B(n14288), .Z(n14283) );
  AND U14276 ( .A(n14289), .B(n14290), .Z(n14288) );
  XOR U14277 ( .A(p_input[81]), .B(n14287), .Z(n14290) );
  XNOR U14278 ( .A(p_input[65]), .B(n14287), .Z(n14289) );
  AND U14279 ( .A(p_input[80]), .B(n14291), .Z(n14287) );
  IV U14280 ( .A(p_input[64]), .Z(n14291) );
  XOR U14281 ( .A(n14292), .B(n14293), .Z(n13850) );
  AND U14282 ( .A(n327), .B(n14294), .Z(n14293) );
  XNOR U14283 ( .A(n14295), .B(n14292), .Z(n14294) );
  XOR U14284 ( .A(n14296), .B(n14297), .Z(n327) );
  AND U14285 ( .A(n14298), .B(n14299), .Z(n14297) );
  XNOR U14286 ( .A(n13861), .B(n14296), .Z(n14299) );
  AND U14287 ( .A(p_input[63]), .B(p_input[47]), .Z(n13861) );
  XOR U14288 ( .A(n14296), .B(n13860), .Z(n14298) );
  AND U14289 ( .A(p_input[15]), .B(p_input[31]), .Z(n13860) );
  XOR U14290 ( .A(n14300), .B(n14301), .Z(n14296) );
  AND U14291 ( .A(n14302), .B(n14303), .Z(n14301) );
  XOR U14292 ( .A(n14300), .B(n13873), .Z(n14303) );
  XNOR U14293 ( .A(p_input[46]), .B(n14304), .Z(n13873) );
  AND U14294 ( .A(n558), .B(n14305), .Z(n14304) );
  XOR U14295 ( .A(p_input[62]), .B(p_input[46]), .Z(n14305) );
  XNOR U14296 ( .A(n13870), .B(n14300), .Z(n14302) );
  XOR U14297 ( .A(n14306), .B(n14307), .Z(n13870) );
  AND U14298 ( .A(n555), .B(n14308), .Z(n14307) );
  XOR U14299 ( .A(p_input[30]), .B(p_input[14]), .Z(n14308) );
  XOR U14300 ( .A(n14309), .B(n14310), .Z(n14300) );
  AND U14301 ( .A(n14311), .B(n14312), .Z(n14310) );
  XOR U14302 ( .A(n14309), .B(n13885), .Z(n14312) );
  XNOR U14303 ( .A(p_input[45]), .B(n14313), .Z(n13885) );
  AND U14304 ( .A(n558), .B(n14314), .Z(n14313) );
  XOR U14305 ( .A(p_input[61]), .B(p_input[45]), .Z(n14314) );
  XNOR U14306 ( .A(n13882), .B(n14309), .Z(n14311) );
  XOR U14307 ( .A(n14315), .B(n14316), .Z(n13882) );
  AND U14308 ( .A(n555), .B(n14317), .Z(n14316) );
  XOR U14309 ( .A(p_input[29]), .B(p_input[13]), .Z(n14317) );
  XOR U14310 ( .A(n14318), .B(n14319), .Z(n14309) );
  AND U14311 ( .A(n14320), .B(n14321), .Z(n14319) );
  XOR U14312 ( .A(n14318), .B(n13897), .Z(n14321) );
  XNOR U14313 ( .A(p_input[44]), .B(n14322), .Z(n13897) );
  AND U14314 ( .A(n558), .B(n14323), .Z(n14322) );
  XOR U14315 ( .A(p_input[60]), .B(p_input[44]), .Z(n14323) );
  XNOR U14316 ( .A(n13894), .B(n14318), .Z(n14320) );
  XOR U14317 ( .A(n14324), .B(n14325), .Z(n13894) );
  AND U14318 ( .A(n555), .B(n14326), .Z(n14325) );
  XOR U14319 ( .A(p_input[28]), .B(p_input[12]), .Z(n14326) );
  XOR U14320 ( .A(n14327), .B(n14328), .Z(n14318) );
  AND U14321 ( .A(n14329), .B(n14330), .Z(n14328) );
  XOR U14322 ( .A(n14327), .B(n13909), .Z(n14330) );
  XNOR U14323 ( .A(p_input[43]), .B(n14331), .Z(n13909) );
  AND U14324 ( .A(n558), .B(n14332), .Z(n14331) );
  XOR U14325 ( .A(p_input[59]), .B(p_input[43]), .Z(n14332) );
  XNOR U14326 ( .A(n13906), .B(n14327), .Z(n14329) );
  XOR U14327 ( .A(n14333), .B(n14334), .Z(n13906) );
  AND U14328 ( .A(n555), .B(n14335), .Z(n14334) );
  XOR U14329 ( .A(p_input[27]), .B(p_input[11]), .Z(n14335) );
  XOR U14330 ( .A(n14336), .B(n14337), .Z(n14327) );
  AND U14331 ( .A(n14338), .B(n14339), .Z(n14337) );
  XOR U14332 ( .A(n14336), .B(n13921), .Z(n14339) );
  XNOR U14333 ( .A(p_input[42]), .B(n14340), .Z(n13921) );
  AND U14334 ( .A(n558), .B(n14341), .Z(n14340) );
  XOR U14335 ( .A(p_input[58]), .B(p_input[42]), .Z(n14341) );
  XNOR U14336 ( .A(n13918), .B(n14336), .Z(n14338) );
  XOR U14337 ( .A(n14342), .B(n14343), .Z(n13918) );
  AND U14338 ( .A(n555), .B(n14344), .Z(n14343) );
  XOR U14339 ( .A(p_input[26]), .B(p_input[10]), .Z(n14344) );
  XOR U14340 ( .A(n14345), .B(n14346), .Z(n14336) );
  AND U14341 ( .A(n14347), .B(n14348), .Z(n14346) );
  XOR U14342 ( .A(n14345), .B(n13933), .Z(n14348) );
  XNOR U14343 ( .A(p_input[41]), .B(n14349), .Z(n13933) );
  AND U14344 ( .A(n558), .B(n14350), .Z(n14349) );
  XOR U14345 ( .A(p_input[57]), .B(p_input[41]), .Z(n14350) );
  XNOR U14346 ( .A(n13930), .B(n14345), .Z(n14347) );
  XOR U14347 ( .A(n14351), .B(n14352), .Z(n13930) );
  AND U14348 ( .A(n555), .B(n14353), .Z(n14352) );
  XOR U14349 ( .A(p_input[9]), .B(p_input[25]), .Z(n14353) );
  XOR U14350 ( .A(n14354), .B(n14355), .Z(n14345) );
  AND U14351 ( .A(n14356), .B(n14357), .Z(n14355) );
  XOR U14352 ( .A(n14354), .B(n13945), .Z(n14357) );
  XNOR U14353 ( .A(p_input[40]), .B(n14358), .Z(n13945) );
  AND U14354 ( .A(n558), .B(n14359), .Z(n14358) );
  XOR U14355 ( .A(p_input[56]), .B(p_input[40]), .Z(n14359) );
  XNOR U14356 ( .A(n13942), .B(n14354), .Z(n14356) );
  XOR U14357 ( .A(n14360), .B(n14361), .Z(n13942) );
  AND U14358 ( .A(n555), .B(n14362), .Z(n14361) );
  XOR U14359 ( .A(p_input[8]), .B(p_input[24]), .Z(n14362) );
  XOR U14360 ( .A(n14363), .B(n14364), .Z(n14354) );
  AND U14361 ( .A(n14365), .B(n14366), .Z(n14364) );
  XOR U14362 ( .A(n14363), .B(n13957), .Z(n14366) );
  XNOR U14363 ( .A(p_input[39]), .B(n14367), .Z(n13957) );
  AND U14364 ( .A(n558), .B(n14368), .Z(n14367) );
  XOR U14365 ( .A(p_input[55]), .B(p_input[39]), .Z(n14368) );
  XNOR U14366 ( .A(n13954), .B(n14363), .Z(n14365) );
  XOR U14367 ( .A(n14369), .B(n14370), .Z(n13954) );
  AND U14368 ( .A(n555), .B(n14371), .Z(n14370) );
  XOR U14369 ( .A(p_input[7]), .B(p_input[23]), .Z(n14371) );
  XOR U14370 ( .A(n14372), .B(n14373), .Z(n14363) );
  AND U14371 ( .A(n14374), .B(n14375), .Z(n14373) );
  XOR U14372 ( .A(n14372), .B(n13969), .Z(n14375) );
  XNOR U14373 ( .A(p_input[38]), .B(n14376), .Z(n13969) );
  AND U14374 ( .A(n558), .B(n14377), .Z(n14376) );
  XOR U14375 ( .A(p_input[54]), .B(p_input[38]), .Z(n14377) );
  XNOR U14376 ( .A(n13966), .B(n14372), .Z(n14374) );
  XOR U14377 ( .A(n14378), .B(n14379), .Z(n13966) );
  AND U14378 ( .A(n555), .B(n14380), .Z(n14379) );
  XOR U14379 ( .A(p_input[6]), .B(p_input[22]), .Z(n14380) );
  XOR U14380 ( .A(n14381), .B(n14382), .Z(n14372) );
  AND U14381 ( .A(n14383), .B(n14384), .Z(n14382) );
  XOR U14382 ( .A(n14381), .B(n13981), .Z(n14384) );
  XNOR U14383 ( .A(p_input[37]), .B(n14385), .Z(n13981) );
  AND U14384 ( .A(n558), .B(n14386), .Z(n14385) );
  XOR U14385 ( .A(p_input[53]), .B(p_input[37]), .Z(n14386) );
  XNOR U14386 ( .A(n13978), .B(n14381), .Z(n14383) );
  XOR U14387 ( .A(n14387), .B(n14388), .Z(n13978) );
  AND U14388 ( .A(n555), .B(n14389), .Z(n14388) );
  XOR U14389 ( .A(p_input[5]), .B(p_input[21]), .Z(n14389) );
  XOR U14390 ( .A(n14390), .B(n14391), .Z(n14381) );
  AND U14391 ( .A(n14392), .B(n14393), .Z(n14391) );
  XOR U14392 ( .A(n14390), .B(n13993), .Z(n14393) );
  XNOR U14393 ( .A(p_input[36]), .B(n14394), .Z(n13993) );
  AND U14394 ( .A(n558), .B(n14395), .Z(n14394) );
  XOR U14395 ( .A(p_input[52]), .B(p_input[36]), .Z(n14395) );
  XNOR U14396 ( .A(n13990), .B(n14390), .Z(n14392) );
  XOR U14397 ( .A(n14396), .B(n14397), .Z(n13990) );
  AND U14398 ( .A(n555), .B(n14398), .Z(n14397) );
  XOR U14399 ( .A(p_input[4]), .B(p_input[20]), .Z(n14398) );
  XOR U14400 ( .A(n14399), .B(n14400), .Z(n14390) );
  AND U14401 ( .A(n14401), .B(n14402), .Z(n14400) );
  XOR U14402 ( .A(n14399), .B(n14005), .Z(n14402) );
  XNOR U14403 ( .A(p_input[35]), .B(n14403), .Z(n14005) );
  AND U14404 ( .A(n558), .B(n14404), .Z(n14403) );
  XOR U14405 ( .A(p_input[51]), .B(p_input[35]), .Z(n14404) );
  XNOR U14406 ( .A(n14002), .B(n14399), .Z(n14401) );
  XOR U14407 ( .A(n14405), .B(n14406), .Z(n14002) );
  AND U14408 ( .A(n555), .B(n14407), .Z(n14406) );
  XOR U14409 ( .A(p_input[3]), .B(p_input[19]), .Z(n14407) );
  XOR U14410 ( .A(n14408), .B(n14409), .Z(n14399) );
  AND U14411 ( .A(n14410), .B(n14411), .Z(n14409) );
  XOR U14412 ( .A(n14017), .B(n14408), .Z(n14411) );
  XNOR U14413 ( .A(p_input[34]), .B(n14412), .Z(n14017) );
  AND U14414 ( .A(n558), .B(n14413), .Z(n14412) );
  XOR U14415 ( .A(p_input[50]), .B(p_input[34]), .Z(n14413) );
  XNOR U14416 ( .A(n14408), .B(n14014), .Z(n14410) );
  XOR U14417 ( .A(n14414), .B(n14415), .Z(n14014) );
  AND U14418 ( .A(n555), .B(n14416), .Z(n14415) );
  XOR U14419 ( .A(p_input[2]), .B(p_input[18]), .Z(n14416) );
  XOR U14420 ( .A(n14417), .B(n14418), .Z(n14408) );
  AND U14421 ( .A(n14419), .B(n14420), .Z(n14418) );
  XNOR U14422 ( .A(n14421), .B(n14030), .Z(n14420) );
  XNOR U14423 ( .A(p_input[33]), .B(n14422), .Z(n14030) );
  AND U14424 ( .A(n558), .B(n14423), .Z(n14422) );
  XNOR U14425 ( .A(p_input[49]), .B(n14424), .Z(n14423) );
  IV U14426 ( .A(p_input[33]), .Z(n14424) );
  XNOR U14427 ( .A(n14027), .B(n14417), .Z(n14419) );
  XNOR U14428 ( .A(p_input[1]), .B(n14425), .Z(n14027) );
  AND U14429 ( .A(n555), .B(n14426), .Z(n14425) );
  XOR U14430 ( .A(p_input[1]), .B(p_input[17]), .Z(n14426) );
  IV U14431 ( .A(n14421), .Z(n14417) );
  AND U14432 ( .A(n14292), .B(n14295), .Z(n14421) );
  XOR U14433 ( .A(p_input[32]), .B(n14427), .Z(n14295) );
  AND U14434 ( .A(n558), .B(n14428), .Z(n14427) );
  XOR U14435 ( .A(p_input[48]), .B(p_input[32]), .Z(n14428) );
  XOR U14436 ( .A(n14429), .B(n14430), .Z(n558) );
  AND U14437 ( .A(n14431), .B(n14432), .Z(n14430) );
  XNOR U14438 ( .A(p_input[63]), .B(n14429), .Z(n14432) );
  XOR U14439 ( .A(n14429), .B(p_input[47]), .Z(n14431) );
  XOR U14440 ( .A(n14433), .B(n14434), .Z(n14429) );
  AND U14441 ( .A(n14435), .B(n14436), .Z(n14434) );
  XNOR U14442 ( .A(p_input[62]), .B(n14433), .Z(n14436) );
  XOR U14443 ( .A(n14433), .B(p_input[46]), .Z(n14435) );
  XOR U14444 ( .A(n14437), .B(n14438), .Z(n14433) );
  AND U14445 ( .A(n14439), .B(n14440), .Z(n14438) );
  XNOR U14446 ( .A(p_input[61]), .B(n14437), .Z(n14440) );
  XOR U14447 ( .A(n14437), .B(p_input[45]), .Z(n14439) );
  XOR U14448 ( .A(n14441), .B(n14442), .Z(n14437) );
  AND U14449 ( .A(n14443), .B(n14444), .Z(n14442) );
  XNOR U14450 ( .A(p_input[60]), .B(n14441), .Z(n14444) );
  XOR U14451 ( .A(n14441), .B(p_input[44]), .Z(n14443) );
  XOR U14452 ( .A(n14445), .B(n14446), .Z(n14441) );
  AND U14453 ( .A(n14447), .B(n14448), .Z(n14446) );
  XNOR U14454 ( .A(p_input[59]), .B(n14445), .Z(n14448) );
  XOR U14455 ( .A(n14445), .B(p_input[43]), .Z(n14447) );
  XOR U14456 ( .A(n14449), .B(n14450), .Z(n14445) );
  AND U14457 ( .A(n14451), .B(n14452), .Z(n14450) );
  XNOR U14458 ( .A(p_input[58]), .B(n14449), .Z(n14452) );
  XOR U14459 ( .A(n14449), .B(p_input[42]), .Z(n14451) );
  XOR U14460 ( .A(n14453), .B(n14454), .Z(n14449) );
  AND U14461 ( .A(n14455), .B(n14456), .Z(n14454) );
  XNOR U14462 ( .A(p_input[57]), .B(n14453), .Z(n14456) );
  XOR U14463 ( .A(n14453), .B(p_input[41]), .Z(n14455) );
  XOR U14464 ( .A(n14457), .B(n14458), .Z(n14453) );
  AND U14465 ( .A(n14459), .B(n14460), .Z(n14458) );
  XNOR U14466 ( .A(p_input[56]), .B(n14457), .Z(n14460) );
  XOR U14467 ( .A(n14457), .B(p_input[40]), .Z(n14459) );
  XOR U14468 ( .A(n14461), .B(n14462), .Z(n14457) );
  AND U14469 ( .A(n14463), .B(n14464), .Z(n14462) );
  XNOR U14470 ( .A(p_input[55]), .B(n14461), .Z(n14464) );
  XOR U14471 ( .A(n14461), .B(p_input[39]), .Z(n14463) );
  XOR U14472 ( .A(n14465), .B(n14466), .Z(n14461) );
  AND U14473 ( .A(n14467), .B(n14468), .Z(n14466) );
  XNOR U14474 ( .A(p_input[54]), .B(n14465), .Z(n14468) );
  XOR U14475 ( .A(n14465), .B(p_input[38]), .Z(n14467) );
  XOR U14476 ( .A(n14469), .B(n14470), .Z(n14465) );
  AND U14477 ( .A(n14471), .B(n14472), .Z(n14470) );
  XNOR U14478 ( .A(p_input[53]), .B(n14469), .Z(n14472) );
  XOR U14479 ( .A(n14469), .B(p_input[37]), .Z(n14471) );
  XOR U14480 ( .A(n14473), .B(n14474), .Z(n14469) );
  AND U14481 ( .A(n14475), .B(n14476), .Z(n14474) );
  XNOR U14482 ( .A(p_input[52]), .B(n14473), .Z(n14476) );
  XOR U14483 ( .A(n14473), .B(p_input[36]), .Z(n14475) );
  XOR U14484 ( .A(n14477), .B(n14478), .Z(n14473) );
  AND U14485 ( .A(n14479), .B(n14480), .Z(n14478) );
  XNOR U14486 ( .A(p_input[51]), .B(n14477), .Z(n14480) );
  XOR U14487 ( .A(n14477), .B(p_input[35]), .Z(n14479) );
  XOR U14488 ( .A(n14481), .B(n14482), .Z(n14477) );
  AND U14489 ( .A(n14483), .B(n14484), .Z(n14482) );
  XNOR U14490 ( .A(p_input[50]), .B(n14481), .Z(n14484) );
  XOR U14491 ( .A(n14481), .B(p_input[34]), .Z(n14483) );
  XNOR U14492 ( .A(n14485), .B(n14486), .Z(n14481) );
  AND U14493 ( .A(n14487), .B(n14488), .Z(n14486) );
  XOR U14494 ( .A(p_input[49]), .B(n14485), .Z(n14488) );
  XNOR U14495 ( .A(p_input[33]), .B(n14485), .Z(n14487) );
  AND U14496 ( .A(p_input[48]), .B(n14489), .Z(n14485) );
  IV U14497 ( .A(p_input[32]), .Z(n14489) );
  XNOR U14498 ( .A(p_input[0]), .B(n14490), .Z(n14292) );
  AND U14499 ( .A(n555), .B(n14491), .Z(n14490) );
  XOR U14500 ( .A(p_input[16]), .B(p_input[0]), .Z(n14491) );
  XOR U14501 ( .A(n14492), .B(n14493), .Z(n555) );
  AND U14502 ( .A(n14494), .B(n14495), .Z(n14493) );
  XNOR U14503 ( .A(p_input[31]), .B(n14492), .Z(n14495) );
  XOR U14504 ( .A(n14492), .B(p_input[15]), .Z(n14494) );
  XOR U14505 ( .A(n14496), .B(n14497), .Z(n14492) );
  AND U14506 ( .A(n14498), .B(n14499), .Z(n14497) );
  XNOR U14507 ( .A(p_input[30]), .B(n14496), .Z(n14499) );
  XNOR U14508 ( .A(n14496), .B(n14306), .Z(n14498) );
  IV U14509 ( .A(p_input[14]), .Z(n14306) );
  XOR U14510 ( .A(n14500), .B(n14501), .Z(n14496) );
  AND U14511 ( .A(n14502), .B(n14503), .Z(n14501) );
  XNOR U14512 ( .A(p_input[29]), .B(n14500), .Z(n14503) );
  XNOR U14513 ( .A(n14500), .B(n14315), .Z(n14502) );
  IV U14514 ( .A(p_input[13]), .Z(n14315) );
  XOR U14515 ( .A(n14504), .B(n14505), .Z(n14500) );
  AND U14516 ( .A(n14506), .B(n14507), .Z(n14505) );
  XNOR U14517 ( .A(p_input[28]), .B(n14504), .Z(n14507) );
  XNOR U14518 ( .A(n14504), .B(n14324), .Z(n14506) );
  IV U14519 ( .A(p_input[12]), .Z(n14324) );
  XOR U14520 ( .A(n14508), .B(n14509), .Z(n14504) );
  AND U14521 ( .A(n14510), .B(n14511), .Z(n14509) );
  XNOR U14522 ( .A(p_input[27]), .B(n14508), .Z(n14511) );
  XNOR U14523 ( .A(n14508), .B(n14333), .Z(n14510) );
  IV U14524 ( .A(p_input[11]), .Z(n14333) );
  XOR U14525 ( .A(n14512), .B(n14513), .Z(n14508) );
  AND U14526 ( .A(n14514), .B(n14515), .Z(n14513) );
  XNOR U14527 ( .A(p_input[26]), .B(n14512), .Z(n14515) );
  XNOR U14528 ( .A(n14512), .B(n14342), .Z(n14514) );
  IV U14529 ( .A(p_input[10]), .Z(n14342) );
  XOR U14530 ( .A(n14516), .B(n14517), .Z(n14512) );
  AND U14531 ( .A(n14518), .B(n14519), .Z(n14517) );
  XNOR U14532 ( .A(p_input[25]), .B(n14516), .Z(n14519) );
  XNOR U14533 ( .A(n14516), .B(n14351), .Z(n14518) );
  IV U14534 ( .A(p_input[9]), .Z(n14351) );
  XOR U14535 ( .A(n14520), .B(n14521), .Z(n14516) );
  AND U14536 ( .A(n14522), .B(n14523), .Z(n14521) );
  XNOR U14537 ( .A(p_input[24]), .B(n14520), .Z(n14523) );
  XNOR U14538 ( .A(n14520), .B(n14360), .Z(n14522) );
  IV U14539 ( .A(p_input[8]), .Z(n14360) );
  XOR U14540 ( .A(n14524), .B(n14525), .Z(n14520) );
  AND U14541 ( .A(n14526), .B(n14527), .Z(n14525) );
  XNOR U14542 ( .A(p_input[23]), .B(n14524), .Z(n14527) );
  XNOR U14543 ( .A(n14524), .B(n14369), .Z(n14526) );
  IV U14544 ( .A(p_input[7]), .Z(n14369) );
  XOR U14545 ( .A(n14528), .B(n14529), .Z(n14524) );
  AND U14546 ( .A(n14530), .B(n14531), .Z(n14529) );
  XNOR U14547 ( .A(p_input[22]), .B(n14528), .Z(n14531) );
  XNOR U14548 ( .A(n14528), .B(n14378), .Z(n14530) );
  IV U14549 ( .A(p_input[6]), .Z(n14378) );
  XOR U14550 ( .A(n14532), .B(n14533), .Z(n14528) );
  AND U14551 ( .A(n14534), .B(n14535), .Z(n14533) );
  XNOR U14552 ( .A(p_input[21]), .B(n14532), .Z(n14535) );
  XNOR U14553 ( .A(n14532), .B(n14387), .Z(n14534) );
  IV U14554 ( .A(p_input[5]), .Z(n14387) );
  XOR U14555 ( .A(n14536), .B(n14537), .Z(n14532) );
  AND U14556 ( .A(n14538), .B(n14539), .Z(n14537) );
  XNOR U14557 ( .A(p_input[20]), .B(n14536), .Z(n14539) );
  XNOR U14558 ( .A(n14536), .B(n14396), .Z(n14538) );
  IV U14559 ( .A(p_input[4]), .Z(n14396) );
  XOR U14560 ( .A(n14540), .B(n14541), .Z(n14536) );
  AND U14561 ( .A(n14542), .B(n14543), .Z(n14541) );
  XNOR U14562 ( .A(p_input[19]), .B(n14540), .Z(n14543) );
  XNOR U14563 ( .A(n14540), .B(n14405), .Z(n14542) );
  IV U14564 ( .A(p_input[3]), .Z(n14405) );
  XOR U14565 ( .A(n14544), .B(n14545), .Z(n14540) );
  AND U14566 ( .A(n14546), .B(n14547), .Z(n14545) );
  XNOR U14567 ( .A(p_input[18]), .B(n14544), .Z(n14547) );
  XNOR U14568 ( .A(n14544), .B(n14414), .Z(n14546) );
  IV U14569 ( .A(p_input[2]), .Z(n14414) );
  XNOR U14570 ( .A(n14548), .B(n14549), .Z(n14544) );
  AND U14571 ( .A(n14550), .B(n14551), .Z(n14549) );
  XOR U14572 ( .A(p_input[17]), .B(n14548), .Z(n14551) );
  XNOR U14573 ( .A(p_input[1]), .B(n14548), .Z(n14550) );
  AND U14574 ( .A(p_input[16]), .B(n14552), .Z(n14548) );
  IV U14575 ( .A(p_input[0]), .Z(n14552) );
endmodule

