
module psi_BMR_b10_n10 ( p_input, o );
  input [99:0] p_input;
  output [9:0] o;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80;

  AND U1 ( .A(n1), .B(n2), .Z(o[9]) );
  AND U2 ( .A(n3), .B(n4), .Z(n2) );
  AND U3 ( .A(n5), .B(p_input[39]), .Z(n4) );
  AND U4 ( .A(p_input[29]), .B(p_input[19]), .Z(n5) );
  AND U5 ( .A(p_input[59]), .B(p_input[49]), .Z(n3) );
  AND U6 ( .A(n6), .B(n7), .Z(n1) );
  AND U7 ( .A(n8), .B(p_input[89]), .Z(n7) );
  AND U8 ( .A(p_input[79]), .B(p_input[69]), .Z(n8) );
  AND U9 ( .A(p_input[9]), .B(p_input[99]), .Z(n6) );
  AND U10 ( .A(n9), .B(n10), .Z(o[8]) );
  AND U11 ( .A(n11), .B(n12), .Z(n10) );
  AND U12 ( .A(n13), .B(p_input[38]), .Z(n12) );
  AND U13 ( .A(p_input[28]), .B(p_input[18]), .Z(n13) );
  AND U14 ( .A(p_input[58]), .B(p_input[48]), .Z(n11) );
  AND U15 ( .A(n14), .B(n15), .Z(n9) );
  AND U16 ( .A(n16), .B(p_input[88]), .Z(n15) );
  AND U17 ( .A(p_input[78]), .B(p_input[68]), .Z(n16) );
  AND U18 ( .A(p_input[98]), .B(p_input[8]), .Z(n14) );
  AND U19 ( .A(n17), .B(n18), .Z(o[7]) );
  AND U20 ( .A(n19), .B(n20), .Z(n18) );
  AND U21 ( .A(n21), .B(p_input[37]), .Z(n20) );
  AND U22 ( .A(p_input[27]), .B(p_input[17]), .Z(n21) );
  AND U23 ( .A(p_input[57]), .B(p_input[47]), .Z(n19) );
  AND U24 ( .A(n22), .B(n23), .Z(n17) );
  AND U25 ( .A(n24), .B(p_input[7]), .Z(n23) );
  AND U26 ( .A(p_input[77]), .B(p_input[67]), .Z(n24) );
  AND U27 ( .A(p_input[97]), .B(p_input[87]), .Z(n22) );
  AND U28 ( .A(n25), .B(n26), .Z(o[6]) );
  AND U29 ( .A(n27), .B(n28), .Z(n26) );
  AND U30 ( .A(n29), .B(p_input[36]), .Z(n28) );
  AND U31 ( .A(p_input[26]), .B(p_input[16]), .Z(n29) );
  AND U32 ( .A(p_input[56]), .B(p_input[46]), .Z(n27) );
  AND U33 ( .A(n30), .B(n31), .Z(n25) );
  AND U34 ( .A(n32), .B(p_input[76]), .Z(n31) );
  AND U35 ( .A(p_input[6]), .B(p_input[66]), .Z(n32) );
  AND U36 ( .A(p_input[96]), .B(p_input[86]), .Z(n30) );
  AND U37 ( .A(n33), .B(n34), .Z(o[5]) );
  AND U38 ( .A(n35), .B(n36), .Z(n34) );
  AND U39 ( .A(n37), .B(p_input[35]), .Z(n36) );
  AND U40 ( .A(p_input[25]), .B(p_input[15]), .Z(n37) );
  AND U41 ( .A(p_input[55]), .B(p_input[45]), .Z(n35) );
  AND U42 ( .A(n38), .B(n39), .Z(n33) );
  AND U43 ( .A(n40), .B(p_input[75]), .Z(n39) );
  AND U44 ( .A(p_input[65]), .B(p_input[5]), .Z(n40) );
  AND U45 ( .A(p_input[95]), .B(p_input[85]), .Z(n38) );
  AND U46 ( .A(n41), .B(n42), .Z(o[4]) );
  AND U47 ( .A(n43), .B(n44), .Z(n42) );
  AND U48 ( .A(n45), .B(p_input[34]), .Z(n44) );
  AND U49 ( .A(p_input[24]), .B(p_input[14]), .Z(n45) );
  AND U50 ( .A(p_input[4]), .B(p_input[44]), .Z(n43) );
  AND U51 ( .A(n46), .B(n47), .Z(n41) );
  AND U52 ( .A(n48), .B(p_input[74]), .Z(n47) );
  AND U53 ( .A(p_input[64]), .B(p_input[54]), .Z(n48) );
  AND U54 ( .A(p_input[94]), .B(p_input[84]), .Z(n46) );
  AND U55 ( .A(n49), .B(n50), .Z(o[3]) );
  AND U56 ( .A(n51), .B(n52), .Z(n50) );
  AND U57 ( .A(n53), .B(p_input[33]), .Z(n52) );
  AND U58 ( .A(p_input[23]), .B(p_input[13]), .Z(n53) );
  AND U59 ( .A(p_input[43]), .B(p_input[3]), .Z(n51) );
  AND U60 ( .A(n54), .B(n55), .Z(n49) );
  AND U61 ( .A(n56), .B(p_input[73]), .Z(n55) );
  AND U62 ( .A(p_input[63]), .B(p_input[53]), .Z(n56) );
  AND U63 ( .A(p_input[93]), .B(p_input[83]), .Z(n54) );
  AND U64 ( .A(n57), .B(n58), .Z(o[2]) );
  AND U65 ( .A(n59), .B(n60), .Z(n58) );
  AND U66 ( .A(n61), .B(p_input[2]), .Z(n60) );
  AND U67 ( .A(p_input[22]), .B(p_input[12]), .Z(n61) );
  AND U68 ( .A(p_input[42]), .B(p_input[32]), .Z(n59) );
  AND U69 ( .A(n62), .B(n63), .Z(n57) );
  AND U70 ( .A(n64), .B(p_input[72]), .Z(n63) );
  AND U71 ( .A(p_input[62]), .B(p_input[52]), .Z(n64) );
  AND U72 ( .A(p_input[92]), .B(p_input[82]), .Z(n62) );
  AND U73 ( .A(n65), .B(n66), .Z(o[1]) );
  AND U74 ( .A(n67), .B(n68), .Z(n66) );
  AND U75 ( .A(n69), .B(p_input[21]), .Z(n68) );
  AND U76 ( .A(p_input[1]), .B(p_input[11]), .Z(n69) );
  AND U77 ( .A(p_input[41]), .B(p_input[31]), .Z(n67) );
  AND U78 ( .A(n70), .B(n71), .Z(n65) );
  AND U79 ( .A(n72), .B(p_input[71]), .Z(n71) );
  AND U80 ( .A(p_input[61]), .B(p_input[51]), .Z(n72) );
  AND U81 ( .A(p_input[91]), .B(p_input[81]), .Z(n70) );
  AND U82 ( .A(n73), .B(n74), .Z(o[0]) );
  AND U83 ( .A(n75), .B(n76), .Z(n74) );
  AND U84 ( .A(n77), .B(p_input[20]), .Z(n76) );
  AND U85 ( .A(p_input[10]), .B(p_input[0]), .Z(n77) );
  AND U86 ( .A(p_input[40]), .B(p_input[30]), .Z(n75) );
  AND U87 ( .A(n78), .B(n79), .Z(n73) );
  AND U88 ( .A(n80), .B(p_input[70]), .Z(n79) );
  AND U89 ( .A(p_input[60]), .B(p_input[50]), .Z(n80) );
  AND U90 ( .A(p_input[90]), .B(p_input[80]), .Z(n78) );
endmodule

