
module auction_BMR_N6_W16 ( p_input, o );
  input [1023:0] p_input;
  output [21:0] o;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972,
         n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982,
         n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992,
         n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002,
         n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
         n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022,
         n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032,
         n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042,
         n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052,
         n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062,
         n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072,
         n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082,
         n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092,
         n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102,
         n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112,
         n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122,
         n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132,
         n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142,
         n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152,
         n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162,
         n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172,
         n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182,
         n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192,
         n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202,
         n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212,
         n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222,
         n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232,
         n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242,
         n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252,
         n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262,
         n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272,
         n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282,
         n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292,
         n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302,
         n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312,
         n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322,
         n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332,
         n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342,
         n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352,
         n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362,
         n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372,
         n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382,
         n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392,
         n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402,
         n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412,
         n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422,
         n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432,
         n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442,
         n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452,
         n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
         n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
         n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
         n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
         n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
         n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612,
         n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622,
         n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632,
         n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
         n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652,
         n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662,
         n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672,
         n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682,
         n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692,
         n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702,
         n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712,
         n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722,
         n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732,
         n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742,
         n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752,
         n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762,
         n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772,
         n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782,
         n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792,
         n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802,
         n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812,
         n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822,
         n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832,
         n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842,
         n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852,
         n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862,
         n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872,
         n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882,
         n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892,
         n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902,
         n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912,
         n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922,
         n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932,
         n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942,
         n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952,
         n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962,
         n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972,
         n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982,
         n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992,
         n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002,
         n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012,
         n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022,
         n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032,
         n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042,
         n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052,
         n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062,
         n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072,
         n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082,
         n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092,
         n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102,
         n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112,
         n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122,
         n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132,
         n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142,
         n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152,
         n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162,
         n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172,
         n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182,
         n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192,
         n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202,
         n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212,
         n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222,
         n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232,
         n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242,
         n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252,
         n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262,
         n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272,
         n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282,
         n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292,
         n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302,
         n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312,
         n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322,
         n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332,
         n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342,
         n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352,
         n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362,
         n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372,
         n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382,
         n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392,
         n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402,
         n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412,
         n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422,
         n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432,
         n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442,
         n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452,
         n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462,
         n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472,
         n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482,
         n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492,
         n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502,
         n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512,
         n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522,
         n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532,
         n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542,
         n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552,
         n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562,
         n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572,
         n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582,
         n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592,
         n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602,
         n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612,
         n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622,
         n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632,
         n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642,
         n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652,
         n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662,
         n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672,
         n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682,
         n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692,
         n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702,
         n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712,
         n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722,
         n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732,
         n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742,
         n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752,
         n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762,
         n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772,
         n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782,
         n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792,
         n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802,
         n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812,
         n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822,
         n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832,
         n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842,
         n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852,
         n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862,
         n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872,
         n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882,
         n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892,
         n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902,
         n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912,
         n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922,
         n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932,
         n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942,
         n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952,
         n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962,
         n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972,
         n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982,
         n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992,
         n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002,
         n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012,
         n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022,
         n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032,
         n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042,
         n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052,
         n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062,
         n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072,
         n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082,
         n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092,
         n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102,
         n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112,
         n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122,
         n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132,
         n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142,
         n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152,
         n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162,
         n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172,
         n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182,
         n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192,
         n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202,
         n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212,
         n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222,
         n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232,
         n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242,
         n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252,
         n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262,
         n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272,
         n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282,
         n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292,
         n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302,
         n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312,
         n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322,
         n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332,
         n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342,
         n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352,
         n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362,
         n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372,
         n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382,
         n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392,
         n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402,
         n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412,
         n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422,
         n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432,
         n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442,
         n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452,
         n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462,
         n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472,
         n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482,
         n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492,
         n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502,
         n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512,
         n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522,
         n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532,
         n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542,
         n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552,
         n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562,
         n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572,
         n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582,
         n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592,
         n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602,
         n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612,
         n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622,
         n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632,
         n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642,
         n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652,
         n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662,
         n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672,
         n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682,
         n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692,
         n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702,
         n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712,
         n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722,
         n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732,
         n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742,
         n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752,
         n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762,
         n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772,
         n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782,
         n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792,
         n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802,
         n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812,
         n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822,
         n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832,
         n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842,
         n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852,
         n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862,
         n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872,
         n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882,
         n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892,
         n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902,
         n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912,
         n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922,
         n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932,
         n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942,
         n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952,
         n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962,
         n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972,
         n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982,
         n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992,
         n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002,
         n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012,
         n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022,
         n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032,
         n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042,
         n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052,
         n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062,
         n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072,
         n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082,
         n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092,
         n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102,
         n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112,
         n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122,
         n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132,
         n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142,
         n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152,
         n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162,
         n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172,
         n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182,
         n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192,
         n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202,
         n7203, n7204, n7205, n7206, n7207, n7208;

  XNOR U1 ( .A(n1), .B(n2), .Z(o[9]) );
  AND U2 ( .A(o[5]), .B(n3), .Z(n1) );
  XOR U3 ( .A(n2), .B(n4), .Z(n3) );
  XOR U4 ( .A(n5), .B(n6), .Z(o[8]) );
  AND U5 ( .A(o[5]), .B(n7), .Z(n5) );
  XOR U6 ( .A(n8), .B(n9), .Z(n7) );
  XOR U7 ( .A(n10), .B(n11), .Z(o[7]) );
  AND U8 ( .A(o[5]), .B(n12), .Z(n10) );
  XOR U9 ( .A(n13), .B(n14), .Z(n12) );
  XNOR U10 ( .A(n15), .B(n16), .Z(o[6]) );
  AND U11 ( .A(o[5]), .B(n17), .Z(n15) );
  XNOR U12 ( .A(n18), .B(n16), .Z(n17) );
  XOR U13 ( .A(n19), .B(n20), .Z(o[21]) );
  AND U14 ( .A(o[5]), .B(n21), .Z(n19) );
  XOR U15 ( .A(n22), .B(n23), .Z(n21) );
  XOR U16 ( .A(n24), .B(n25), .Z(o[20]) );
  AND U17 ( .A(o[5]), .B(n26), .Z(n24) );
  XOR U18 ( .A(n27), .B(n28), .Z(n26) );
  XOR U19 ( .A(n29), .B(n30), .Z(o[19]) );
  AND U20 ( .A(o[5]), .B(n31), .Z(n29) );
  XOR U21 ( .A(n32), .B(n33), .Z(n31) );
  XOR U22 ( .A(n34), .B(n35), .Z(o[18]) );
  AND U23 ( .A(o[5]), .B(n36), .Z(n34) );
  XOR U24 ( .A(n37), .B(n38), .Z(n36) );
  XOR U25 ( .A(n39), .B(n40), .Z(o[17]) );
  AND U26 ( .A(o[5]), .B(n41), .Z(n39) );
  XOR U27 ( .A(n42), .B(n43), .Z(n41) );
  XOR U28 ( .A(n44), .B(n45), .Z(o[16]) );
  AND U29 ( .A(o[5]), .B(n46), .Z(n44) );
  XOR U30 ( .A(n47), .B(n48), .Z(n46) );
  XOR U31 ( .A(n49), .B(n50), .Z(o[15]) );
  AND U32 ( .A(o[5]), .B(n51), .Z(n49) );
  XOR U33 ( .A(n52), .B(n53), .Z(n51) );
  XOR U34 ( .A(n54), .B(n55), .Z(o[14]) );
  AND U35 ( .A(o[5]), .B(n56), .Z(n54) );
  XOR U36 ( .A(n57), .B(n58), .Z(n56) );
  XOR U37 ( .A(n59), .B(n60), .Z(o[13]) );
  AND U38 ( .A(o[5]), .B(n61), .Z(n59) );
  XOR U39 ( .A(n62), .B(n63), .Z(n61) );
  XOR U40 ( .A(n64), .B(n65), .Z(o[12]) );
  AND U41 ( .A(o[5]), .B(n66), .Z(n64) );
  XOR U42 ( .A(n67), .B(n68), .Z(n66) );
  XOR U43 ( .A(n69), .B(n70), .Z(o[11]) );
  AND U44 ( .A(o[5]), .B(n71), .Z(n69) );
  XOR U45 ( .A(n72), .B(n73), .Z(n71) );
  XOR U46 ( .A(n74), .B(n75), .Z(o[10]) );
  AND U47 ( .A(o[5]), .B(n76), .Z(n74) );
  XOR U48 ( .A(n77), .B(n78), .Z(n76) );
  XOR U49 ( .A(n79), .B(n80), .Z(o[0]) );
  AND U50 ( .A(o[1]), .B(n81), .Z(n80) );
  XNOR U51 ( .A(n82), .B(n83), .Z(n81) );
  XNOR U52 ( .A(n84), .B(n79), .Z(n83) );
  AND U53 ( .A(o[2]), .B(n85), .Z(n84) );
  XNOR U54 ( .A(n86), .B(n87), .Z(n85) );
  XNOR U55 ( .A(n88), .B(n82), .Z(n87) );
  AND U56 ( .A(o[3]), .B(n89), .Z(n88) );
  XNOR U57 ( .A(n90), .B(n91), .Z(n89) );
  XNOR U58 ( .A(n92), .B(n86), .Z(n91) );
  AND U59 ( .A(o[4]), .B(n93), .Z(n92) );
  XNOR U60 ( .A(n90), .B(n94), .Z(n93) );
  XNOR U61 ( .A(n95), .B(n96), .Z(n94) );
  AND U62 ( .A(o[5]), .B(n97), .Z(n95) );
  XOR U63 ( .A(n96), .B(n98), .Z(n97) );
  XOR U64 ( .A(n99), .B(n100), .Z(n90) );
  AND U65 ( .A(o[5]), .B(n101), .Z(n100) );
  XOR U66 ( .A(n99), .B(n102), .Z(n101) );
  XOR U67 ( .A(n103), .B(n104), .Z(n86) );
  AND U68 ( .A(o[4]), .B(n105), .Z(n104) );
  XNOR U69 ( .A(n103), .B(n106), .Z(n105) );
  XNOR U70 ( .A(n107), .B(n108), .Z(n106) );
  AND U71 ( .A(o[5]), .B(n109), .Z(n107) );
  XOR U72 ( .A(n108), .B(n110), .Z(n109) );
  XOR U73 ( .A(n111), .B(n112), .Z(n103) );
  AND U74 ( .A(o[5]), .B(n113), .Z(n112) );
  XOR U75 ( .A(n111), .B(n114), .Z(n113) );
  XOR U76 ( .A(n115), .B(n116), .Z(n82) );
  AND U77 ( .A(o[3]), .B(n117), .Z(n116) );
  XNOR U78 ( .A(n118), .B(n119), .Z(n117) );
  XNOR U79 ( .A(n120), .B(n115), .Z(n119) );
  AND U80 ( .A(o[4]), .B(n121), .Z(n120) );
  XNOR U81 ( .A(n118), .B(n122), .Z(n121) );
  XNOR U82 ( .A(n123), .B(n124), .Z(n122) );
  AND U83 ( .A(o[5]), .B(n125), .Z(n123) );
  XOR U84 ( .A(n124), .B(n126), .Z(n125) );
  XOR U85 ( .A(n127), .B(n128), .Z(n118) );
  AND U86 ( .A(o[5]), .B(n129), .Z(n128) );
  XOR U87 ( .A(n127), .B(n130), .Z(n129) );
  XOR U88 ( .A(n131), .B(n132), .Z(n115) );
  AND U89 ( .A(o[4]), .B(n133), .Z(n132) );
  XNOR U90 ( .A(n131), .B(n134), .Z(n133) );
  XNOR U91 ( .A(n135), .B(n136), .Z(n134) );
  AND U92 ( .A(o[5]), .B(n137), .Z(n135) );
  XOR U93 ( .A(n136), .B(n138), .Z(n137) );
  XOR U94 ( .A(n139), .B(n140), .Z(n131) );
  AND U95 ( .A(o[5]), .B(n141), .Z(n140) );
  XOR U96 ( .A(n139), .B(n142), .Z(n141) );
  XOR U97 ( .A(n143), .B(n144), .Z(o[1]) );
  AND U98 ( .A(o[2]), .B(n145), .Z(n144) );
  XNOR U99 ( .A(n146), .B(n147), .Z(n145) );
  XNOR U100 ( .A(n148), .B(n143), .Z(n147) );
  AND U101 ( .A(o[3]), .B(n149), .Z(n148) );
  XNOR U102 ( .A(n150), .B(n151), .Z(n149) );
  XNOR U103 ( .A(n152), .B(n146), .Z(n151) );
  AND U104 ( .A(o[4]), .B(n153), .Z(n152) );
  XNOR U105 ( .A(n150), .B(n154), .Z(n153) );
  XNOR U106 ( .A(n155), .B(n156), .Z(n154) );
  AND U107 ( .A(o[5]), .B(n157), .Z(n155) );
  XOR U108 ( .A(n156), .B(n158), .Z(n157) );
  XOR U109 ( .A(n159), .B(n160), .Z(n150) );
  AND U110 ( .A(o[5]), .B(n161), .Z(n160) );
  XOR U111 ( .A(n159), .B(n162), .Z(n161) );
  XOR U112 ( .A(n163), .B(n164), .Z(n146) );
  AND U113 ( .A(o[4]), .B(n165), .Z(n164) );
  XNOR U114 ( .A(n163), .B(n166), .Z(n165) );
  XNOR U115 ( .A(n167), .B(n168), .Z(n166) );
  AND U116 ( .A(o[5]), .B(n169), .Z(n167) );
  XOR U117 ( .A(n168), .B(n170), .Z(n169) );
  XOR U118 ( .A(n171), .B(n172), .Z(n163) );
  AND U119 ( .A(o[5]), .B(n173), .Z(n172) );
  XOR U120 ( .A(n171), .B(n174), .Z(n173) );
  XOR U121 ( .A(n175), .B(n176), .Z(n143) );
  AND U122 ( .A(o[3]), .B(n177), .Z(n176) );
  XNOR U123 ( .A(n178), .B(n179), .Z(n177) );
  XNOR U124 ( .A(n180), .B(n175), .Z(n179) );
  AND U125 ( .A(o[4]), .B(n181), .Z(n180) );
  XNOR U126 ( .A(n178), .B(n182), .Z(n181) );
  XNOR U127 ( .A(n183), .B(n184), .Z(n182) );
  AND U128 ( .A(o[5]), .B(n185), .Z(n183) );
  XOR U129 ( .A(n184), .B(n186), .Z(n185) );
  XOR U130 ( .A(n187), .B(n188), .Z(n178) );
  AND U131 ( .A(o[5]), .B(n189), .Z(n188) );
  XOR U132 ( .A(n187), .B(n190), .Z(n189) );
  XOR U133 ( .A(n191), .B(n192), .Z(n175) );
  AND U134 ( .A(o[4]), .B(n193), .Z(n192) );
  XNOR U135 ( .A(n191), .B(n194), .Z(n193) );
  XNOR U136 ( .A(n195), .B(n196), .Z(n194) );
  AND U137 ( .A(o[5]), .B(n197), .Z(n195) );
  XOR U138 ( .A(n196), .B(n198), .Z(n197) );
  XOR U139 ( .A(n199), .B(n200), .Z(n191) );
  AND U140 ( .A(o[5]), .B(n201), .Z(n200) );
  XOR U141 ( .A(n199), .B(n202), .Z(n201) );
  XOR U142 ( .A(n203), .B(n204), .Z(n79) );
  AND U143 ( .A(o[2]), .B(n205), .Z(n204) );
  XNOR U144 ( .A(n206), .B(n207), .Z(n205) );
  XNOR U145 ( .A(n208), .B(n203), .Z(n207) );
  AND U146 ( .A(o[3]), .B(n209), .Z(n208) );
  XNOR U147 ( .A(n210), .B(n211), .Z(n209) );
  XNOR U148 ( .A(n212), .B(n206), .Z(n211) );
  AND U149 ( .A(o[4]), .B(n213), .Z(n212) );
  XNOR U150 ( .A(n210), .B(n214), .Z(n213) );
  XNOR U151 ( .A(n215), .B(n216), .Z(n214) );
  AND U152 ( .A(o[5]), .B(n217), .Z(n215) );
  XOR U153 ( .A(n216), .B(n218), .Z(n217) );
  XOR U154 ( .A(n219), .B(n220), .Z(n210) );
  AND U155 ( .A(o[5]), .B(n221), .Z(n220) );
  XOR U156 ( .A(n219), .B(n222), .Z(n221) );
  XOR U157 ( .A(n223), .B(n224), .Z(n206) );
  AND U158 ( .A(o[4]), .B(n225), .Z(n224) );
  XNOR U159 ( .A(n223), .B(n226), .Z(n225) );
  XNOR U160 ( .A(n227), .B(n228), .Z(n226) );
  AND U161 ( .A(o[5]), .B(n229), .Z(n227) );
  XOR U162 ( .A(n228), .B(n230), .Z(n229) );
  XOR U163 ( .A(n231), .B(n232), .Z(n223) );
  AND U164 ( .A(o[5]), .B(n233), .Z(n232) );
  XOR U165 ( .A(n231), .B(n234), .Z(n233) );
  XOR U166 ( .A(n235), .B(n236), .Z(o[2]) );
  AND U167 ( .A(o[3]), .B(n237), .Z(n236) );
  XNOR U168 ( .A(n238), .B(n239), .Z(n237) );
  XNOR U169 ( .A(n240), .B(n235), .Z(n239) );
  AND U170 ( .A(o[4]), .B(n241), .Z(n240) );
  XNOR U171 ( .A(n238), .B(n242), .Z(n241) );
  XNOR U172 ( .A(n243), .B(n244), .Z(n242) );
  AND U173 ( .A(o[5]), .B(n245), .Z(n243) );
  XOR U174 ( .A(n244), .B(n246), .Z(n245) );
  XOR U175 ( .A(n247), .B(n248), .Z(n238) );
  AND U176 ( .A(o[5]), .B(n249), .Z(n248) );
  XOR U177 ( .A(n247), .B(n250), .Z(n249) );
  XOR U178 ( .A(n251), .B(n252), .Z(n235) );
  AND U179 ( .A(o[4]), .B(n253), .Z(n252) );
  XNOR U180 ( .A(n251), .B(n254), .Z(n253) );
  XNOR U181 ( .A(n255), .B(n256), .Z(n254) );
  AND U182 ( .A(o[5]), .B(n257), .Z(n255) );
  XOR U183 ( .A(n256), .B(n258), .Z(n257) );
  XOR U184 ( .A(n259), .B(n260), .Z(n251) );
  AND U185 ( .A(o[5]), .B(n261), .Z(n260) );
  XOR U186 ( .A(n259), .B(n262), .Z(n261) );
  XOR U187 ( .A(n263), .B(n264), .Z(n203) );
  AND U188 ( .A(o[3]), .B(n265), .Z(n264) );
  XNOR U189 ( .A(n266), .B(n267), .Z(n265) );
  XNOR U190 ( .A(n268), .B(n263), .Z(n267) );
  AND U191 ( .A(o[4]), .B(n269), .Z(n268) );
  XNOR U192 ( .A(n266), .B(n270), .Z(n269) );
  XNOR U193 ( .A(n271), .B(n272), .Z(n270) );
  AND U194 ( .A(o[5]), .B(n273), .Z(n271) );
  XOR U195 ( .A(n272), .B(n274), .Z(n273) );
  XOR U196 ( .A(n275), .B(n276), .Z(n266) );
  AND U197 ( .A(o[5]), .B(n277), .Z(n276) );
  XOR U198 ( .A(n275), .B(n278), .Z(n277) );
  XOR U199 ( .A(n279), .B(n280), .Z(o[3]) );
  AND U200 ( .A(o[4]), .B(n281), .Z(n280) );
  XNOR U201 ( .A(n279), .B(n282), .Z(n281) );
  XNOR U202 ( .A(n283), .B(n284), .Z(n282) );
  AND U203 ( .A(o[5]), .B(n285), .Z(n283) );
  XOR U204 ( .A(n284), .B(n286), .Z(n285) );
  XOR U205 ( .A(n287), .B(n288), .Z(n279) );
  AND U206 ( .A(o[5]), .B(n289), .Z(n288) );
  XOR U207 ( .A(n287), .B(n290), .Z(n289) );
  XOR U208 ( .A(n291), .B(n292), .Z(n263) );
  AND U209 ( .A(o[4]), .B(n293), .Z(n292) );
  XNOR U210 ( .A(n291), .B(n294), .Z(n293) );
  XNOR U211 ( .A(n295), .B(n296), .Z(n294) );
  AND U212 ( .A(o[5]), .B(n297), .Z(n295) );
  XOR U213 ( .A(n296), .B(n298), .Z(n297) );
  XOR U214 ( .A(n299), .B(n300), .Z(o[4]) );
  AND U215 ( .A(o[5]), .B(n301), .Z(n300) );
  XOR U216 ( .A(n299), .B(n302), .Z(n301) );
  XOR U217 ( .A(n303), .B(n304), .Z(n291) );
  AND U218 ( .A(o[5]), .B(n305), .Z(n304) );
  XOR U219 ( .A(n303), .B(n306), .Z(n305) );
  XOR U220 ( .A(n307), .B(n308), .Z(o[5]) );
  AND U221 ( .A(n309), .B(n310), .Z(n308) );
  XOR U222 ( .A(n307), .B(n22), .Z(n310) );
  XOR U223 ( .A(n311), .B(n312), .Z(n22) );
  AND U224 ( .A(n302), .B(n313), .Z(n312) );
  XOR U225 ( .A(n314), .B(n311), .Z(n313) );
  XNOR U226 ( .A(n23), .B(n307), .Z(n309) );
  IV U227 ( .A(n20), .Z(n23) );
  XNOR U228 ( .A(n315), .B(n316), .Z(n20) );
  AND U229 ( .A(n299), .B(n317), .Z(n316) );
  XOR U230 ( .A(n318), .B(n315), .Z(n317) );
  XOR U231 ( .A(n319), .B(n320), .Z(n307) );
  AND U232 ( .A(n321), .B(n322), .Z(n320) );
  XOR U233 ( .A(n319), .B(n27), .Z(n322) );
  XOR U234 ( .A(n323), .B(n324), .Z(n27) );
  AND U235 ( .A(n302), .B(n325), .Z(n324) );
  XOR U236 ( .A(n326), .B(n323), .Z(n325) );
  XNOR U237 ( .A(n28), .B(n319), .Z(n321) );
  IV U238 ( .A(n25), .Z(n28) );
  XNOR U239 ( .A(n327), .B(n328), .Z(n25) );
  AND U240 ( .A(n299), .B(n329), .Z(n328) );
  XOR U241 ( .A(n330), .B(n327), .Z(n329) );
  XOR U242 ( .A(n331), .B(n332), .Z(n319) );
  AND U243 ( .A(n333), .B(n334), .Z(n332) );
  XOR U244 ( .A(n331), .B(n32), .Z(n334) );
  XOR U245 ( .A(n335), .B(n336), .Z(n32) );
  AND U246 ( .A(n302), .B(n337), .Z(n336) );
  XOR U247 ( .A(n338), .B(n335), .Z(n337) );
  XNOR U248 ( .A(n33), .B(n331), .Z(n333) );
  IV U249 ( .A(n30), .Z(n33) );
  XNOR U250 ( .A(n339), .B(n340), .Z(n30) );
  AND U251 ( .A(n299), .B(n341), .Z(n340) );
  XOR U252 ( .A(n342), .B(n339), .Z(n341) );
  XOR U253 ( .A(n343), .B(n344), .Z(n331) );
  AND U254 ( .A(n345), .B(n346), .Z(n344) );
  XOR U255 ( .A(n343), .B(n37), .Z(n346) );
  XOR U256 ( .A(n347), .B(n348), .Z(n37) );
  AND U257 ( .A(n302), .B(n349), .Z(n348) );
  XOR U258 ( .A(n350), .B(n347), .Z(n349) );
  XNOR U259 ( .A(n38), .B(n343), .Z(n345) );
  IV U260 ( .A(n35), .Z(n38) );
  XNOR U261 ( .A(n351), .B(n352), .Z(n35) );
  AND U262 ( .A(n299), .B(n353), .Z(n352) );
  XOR U263 ( .A(n354), .B(n351), .Z(n353) );
  XOR U264 ( .A(n355), .B(n356), .Z(n343) );
  AND U265 ( .A(n357), .B(n358), .Z(n356) );
  XOR U266 ( .A(n355), .B(n42), .Z(n358) );
  XOR U267 ( .A(n359), .B(n360), .Z(n42) );
  AND U268 ( .A(n302), .B(n361), .Z(n360) );
  XOR U269 ( .A(n362), .B(n359), .Z(n361) );
  XNOR U270 ( .A(n43), .B(n355), .Z(n357) );
  IV U271 ( .A(n40), .Z(n43) );
  XNOR U272 ( .A(n363), .B(n364), .Z(n40) );
  AND U273 ( .A(n299), .B(n365), .Z(n364) );
  XOR U274 ( .A(n366), .B(n363), .Z(n365) );
  XOR U275 ( .A(n367), .B(n368), .Z(n355) );
  AND U276 ( .A(n369), .B(n370), .Z(n368) );
  XOR U277 ( .A(n367), .B(n47), .Z(n370) );
  XOR U278 ( .A(n371), .B(n372), .Z(n47) );
  AND U279 ( .A(n302), .B(n373), .Z(n372) );
  XOR U280 ( .A(n374), .B(n371), .Z(n373) );
  XNOR U281 ( .A(n48), .B(n367), .Z(n369) );
  IV U282 ( .A(n45), .Z(n48) );
  XNOR U283 ( .A(n375), .B(n376), .Z(n45) );
  AND U284 ( .A(n299), .B(n377), .Z(n376) );
  XOR U285 ( .A(n378), .B(n375), .Z(n377) );
  XOR U286 ( .A(n379), .B(n380), .Z(n367) );
  AND U287 ( .A(n381), .B(n382), .Z(n380) );
  XOR U288 ( .A(n379), .B(n52), .Z(n382) );
  XOR U289 ( .A(n383), .B(n384), .Z(n52) );
  AND U290 ( .A(n302), .B(n385), .Z(n384) );
  XOR U291 ( .A(n386), .B(n383), .Z(n385) );
  XNOR U292 ( .A(n53), .B(n379), .Z(n381) );
  IV U293 ( .A(n50), .Z(n53) );
  XNOR U294 ( .A(n387), .B(n388), .Z(n50) );
  AND U295 ( .A(n299), .B(n389), .Z(n388) );
  XOR U296 ( .A(n390), .B(n387), .Z(n389) );
  XOR U297 ( .A(n391), .B(n392), .Z(n379) );
  AND U298 ( .A(n393), .B(n394), .Z(n392) );
  XOR U299 ( .A(n391), .B(n57), .Z(n394) );
  XOR U300 ( .A(n395), .B(n396), .Z(n57) );
  AND U301 ( .A(n302), .B(n397), .Z(n396) );
  XOR U302 ( .A(n398), .B(n395), .Z(n397) );
  XNOR U303 ( .A(n58), .B(n391), .Z(n393) );
  IV U304 ( .A(n55), .Z(n58) );
  XNOR U305 ( .A(n399), .B(n400), .Z(n55) );
  AND U306 ( .A(n299), .B(n401), .Z(n400) );
  XOR U307 ( .A(n402), .B(n399), .Z(n401) );
  XOR U308 ( .A(n403), .B(n404), .Z(n391) );
  AND U309 ( .A(n405), .B(n406), .Z(n404) );
  XOR U310 ( .A(n403), .B(n62), .Z(n406) );
  XOR U311 ( .A(n407), .B(n408), .Z(n62) );
  AND U312 ( .A(n302), .B(n409), .Z(n408) );
  XOR U313 ( .A(n410), .B(n407), .Z(n409) );
  XNOR U314 ( .A(n63), .B(n403), .Z(n405) );
  IV U315 ( .A(n60), .Z(n63) );
  XNOR U316 ( .A(n411), .B(n412), .Z(n60) );
  AND U317 ( .A(n299), .B(n413), .Z(n412) );
  XOR U318 ( .A(n414), .B(n411), .Z(n413) );
  XOR U319 ( .A(n415), .B(n416), .Z(n403) );
  AND U320 ( .A(n417), .B(n418), .Z(n416) );
  XOR U321 ( .A(n415), .B(n67), .Z(n418) );
  XOR U322 ( .A(n419), .B(n420), .Z(n67) );
  AND U323 ( .A(n302), .B(n421), .Z(n420) );
  XOR U324 ( .A(n422), .B(n419), .Z(n421) );
  XNOR U325 ( .A(n68), .B(n415), .Z(n417) );
  IV U326 ( .A(n65), .Z(n68) );
  XNOR U327 ( .A(n423), .B(n424), .Z(n65) );
  AND U328 ( .A(n299), .B(n425), .Z(n424) );
  XOR U329 ( .A(n426), .B(n423), .Z(n425) );
  XOR U330 ( .A(n427), .B(n428), .Z(n415) );
  AND U331 ( .A(n429), .B(n430), .Z(n428) );
  XOR U332 ( .A(n427), .B(n72), .Z(n430) );
  XOR U333 ( .A(n431), .B(n432), .Z(n72) );
  AND U334 ( .A(n302), .B(n433), .Z(n432) );
  XOR U335 ( .A(n434), .B(n431), .Z(n433) );
  XNOR U336 ( .A(n73), .B(n427), .Z(n429) );
  IV U337 ( .A(n70), .Z(n73) );
  XNOR U338 ( .A(n435), .B(n436), .Z(n70) );
  AND U339 ( .A(n299), .B(n437), .Z(n436) );
  XOR U340 ( .A(n438), .B(n435), .Z(n437) );
  XOR U341 ( .A(n439), .B(n440), .Z(n427) );
  AND U342 ( .A(n441), .B(n442), .Z(n440) );
  XOR U343 ( .A(n439), .B(n77), .Z(n442) );
  XOR U344 ( .A(n443), .B(n444), .Z(n77) );
  AND U345 ( .A(n302), .B(n445), .Z(n444) );
  XOR U346 ( .A(n446), .B(n443), .Z(n445) );
  XNOR U347 ( .A(n78), .B(n439), .Z(n441) );
  IV U348 ( .A(n75), .Z(n78) );
  XNOR U349 ( .A(n447), .B(n448), .Z(n75) );
  AND U350 ( .A(n299), .B(n449), .Z(n448) );
  XOR U351 ( .A(n450), .B(n447), .Z(n449) );
  XOR U352 ( .A(n451), .B(n452), .Z(n439) );
  AND U353 ( .A(n453), .B(n454), .Z(n452) );
  XOR U354 ( .A(n4), .B(n451), .Z(n454) );
  XOR U355 ( .A(n455), .B(n456), .Z(n4) );
  AND U356 ( .A(n302), .B(n457), .Z(n456) );
  XOR U357 ( .A(n455), .B(n458), .Z(n457) );
  XNOR U358 ( .A(n451), .B(n2), .Z(n453) );
  XOR U359 ( .A(n459), .B(n460), .Z(n2) );
  AND U360 ( .A(n299), .B(n461), .Z(n460) );
  XOR U361 ( .A(n459), .B(n462), .Z(n461) );
  XOR U362 ( .A(n463), .B(n464), .Z(n451) );
  AND U363 ( .A(n465), .B(n466), .Z(n464) );
  XOR U364 ( .A(n463), .B(n8), .Z(n466) );
  XOR U365 ( .A(n467), .B(n468), .Z(n8) );
  AND U366 ( .A(n302), .B(n469), .Z(n468) );
  XOR U367 ( .A(n470), .B(n467), .Z(n469) );
  XNOR U368 ( .A(n9), .B(n463), .Z(n465) );
  IV U369 ( .A(n6), .Z(n9) );
  XNOR U370 ( .A(n471), .B(n472), .Z(n6) );
  AND U371 ( .A(n299), .B(n473), .Z(n472) );
  XOR U372 ( .A(n474), .B(n471), .Z(n473) );
  XNOR U373 ( .A(n475), .B(n476), .Z(n463) );
  AND U374 ( .A(n477), .B(n478), .Z(n476) );
  XNOR U375 ( .A(n475), .B(n13), .Z(n478) );
  XOR U376 ( .A(n479), .B(n480), .Z(n13) );
  AND U377 ( .A(n302), .B(n481), .Z(n480) );
  XOR U378 ( .A(n482), .B(n479), .Z(n481) );
  XOR U379 ( .A(n14), .B(n475), .Z(n477) );
  IV U380 ( .A(n11), .Z(n14) );
  XNOR U381 ( .A(n483), .B(n484), .Z(n11) );
  AND U382 ( .A(n299), .B(n485), .Z(n484) );
  XOR U383 ( .A(n486), .B(n483), .Z(n485) );
  AND U384 ( .A(n16), .B(n18), .Z(n475) );
  XNOR U385 ( .A(n487), .B(n488), .Z(n18) );
  AND U386 ( .A(n302), .B(n489), .Z(n488) );
  XNOR U387 ( .A(n490), .B(n487), .Z(n489) );
  XOR U388 ( .A(n491), .B(n492), .Z(n302) );
  AND U389 ( .A(n493), .B(n494), .Z(n492) );
  XOR U390 ( .A(n491), .B(n314), .Z(n494) );
  XNOR U391 ( .A(n495), .B(n496), .Z(n314) );
  AND U392 ( .A(n497), .B(n286), .Z(n496) );
  AND U393 ( .A(n495), .B(n498), .Z(n497) );
  XNOR U394 ( .A(n311), .B(n491), .Z(n493) );
  XOR U395 ( .A(n499), .B(n500), .Z(n311) );
  AND U396 ( .A(n501), .B(n284), .Z(n500) );
  NOR U397 ( .A(n499), .B(n502), .Z(n501) );
  XOR U398 ( .A(n503), .B(n504), .Z(n491) );
  AND U399 ( .A(n505), .B(n506), .Z(n504) );
  XOR U400 ( .A(n503), .B(n326), .Z(n506) );
  XOR U401 ( .A(n507), .B(n508), .Z(n326) );
  AND U402 ( .A(n286), .B(n509), .Z(n508) );
  XOR U403 ( .A(n510), .B(n507), .Z(n509) );
  XNOR U404 ( .A(n323), .B(n503), .Z(n505) );
  XOR U405 ( .A(n511), .B(n512), .Z(n323) );
  AND U406 ( .A(n284), .B(n513), .Z(n512) );
  XOR U407 ( .A(n514), .B(n511), .Z(n513) );
  XOR U408 ( .A(n515), .B(n516), .Z(n503) );
  AND U409 ( .A(n517), .B(n518), .Z(n516) );
  XOR U410 ( .A(n515), .B(n338), .Z(n518) );
  XOR U411 ( .A(n519), .B(n520), .Z(n338) );
  AND U412 ( .A(n286), .B(n521), .Z(n520) );
  XOR U413 ( .A(n522), .B(n519), .Z(n521) );
  XNOR U414 ( .A(n335), .B(n515), .Z(n517) );
  XOR U415 ( .A(n523), .B(n524), .Z(n335) );
  AND U416 ( .A(n284), .B(n525), .Z(n524) );
  XOR U417 ( .A(n526), .B(n523), .Z(n525) );
  XOR U418 ( .A(n527), .B(n528), .Z(n515) );
  AND U419 ( .A(n529), .B(n530), .Z(n528) );
  XOR U420 ( .A(n527), .B(n350), .Z(n530) );
  XOR U421 ( .A(n531), .B(n532), .Z(n350) );
  AND U422 ( .A(n286), .B(n533), .Z(n532) );
  XOR U423 ( .A(n534), .B(n531), .Z(n533) );
  XNOR U424 ( .A(n347), .B(n527), .Z(n529) );
  XOR U425 ( .A(n535), .B(n536), .Z(n347) );
  AND U426 ( .A(n284), .B(n537), .Z(n536) );
  XOR U427 ( .A(n538), .B(n535), .Z(n537) );
  XOR U428 ( .A(n539), .B(n540), .Z(n527) );
  AND U429 ( .A(n541), .B(n542), .Z(n540) );
  XOR U430 ( .A(n539), .B(n362), .Z(n542) );
  XOR U431 ( .A(n543), .B(n544), .Z(n362) );
  AND U432 ( .A(n286), .B(n545), .Z(n544) );
  XOR U433 ( .A(n546), .B(n543), .Z(n545) );
  XNOR U434 ( .A(n359), .B(n539), .Z(n541) );
  XOR U435 ( .A(n547), .B(n548), .Z(n359) );
  AND U436 ( .A(n284), .B(n549), .Z(n548) );
  XOR U437 ( .A(n550), .B(n547), .Z(n549) );
  XOR U438 ( .A(n551), .B(n552), .Z(n539) );
  AND U439 ( .A(n553), .B(n554), .Z(n552) );
  XOR U440 ( .A(n551), .B(n374), .Z(n554) );
  XOR U441 ( .A(n555), .B(n556), .Z(n374) );
  AND U442 ( .A(n286), .B(n557), .Z(n556) );
  XOR U443 ( .A(n558), .B(n555), .Z(n557) );
  XNOR U444 ( .A(n371), .B(n551), .Z(n553) );
  XOR U445 ( .A(n559), .B(n560), .Z(n371) );
  AND U446 ( .A(n284), .B(n561), .Z(n560) );
  XOR U447 ( .A(n562), .B(n559), .Z(n561) );
  XOR U448 ( .A(n563), .B(n564), .Z(n551) );
  AND U449 ( .A(n565), .B(n566), .Z(n564) );
  XOR U450 ( .A(n563), .B(n386), .Z(n566) );
  XOR U451 ( .A(n567), .B(n568), .Z(n386) );
  AND U452 ( .A(n286), .B(n569), .Z(n568) );
  XOR U453 ( .A(n570), .B(n567), .Z(n569) );
  XNOR U454 ( .A(n383), .B(n563), .Z(n565) );
  XOR U455 ( .A(n571), .B(n572), .Z(n383) );
  AND U456 ( .A(n284), .B(n573), .Z(n572) );
  XOR U457 ( .A(n574), .B(n571), .Z(n573) );
  XOR U458 ( .A(n575), .B(n576), .Z(n563) );
  AND U459 ( .A(n577), .B(n578), .Z(n576) );
  XOR U460 ( .A(n575), .B(n398), .Z(n578) );
  XOR U461 ( .A(n579), .B(n580), .Z(n398) );
  AND U462 ( .A(n286), .B(n581), .Z(n580) );
  XOR U463 ( .A(n582), .B(n579), .Z(n581) );
  XNOR U464 ( .A(n395), .B(n575), .Z(n577) );
  XOR U465 ( .A(n583), .B(n584), .Z(n395) );
  AND U466 ( .A(n284), .B(n585), .Z(n584) );
  XOR U467 ( .A(n586), .B(n583), .Z(n585) );
  XOR U468 ( .A(n587), .B(n588), .Z(n575) );
  AND U469 ( .A(n589), .B(n590), .Z(n588) );
  XOR U470 ( .A(n587), .B(n410), .Z(n590) );
  XOR U471 ( .A(n591), .B(n592), .Z(n410) );
  AND U472 ( .A(n286), .B(n593), .Z(n592) );
  XOR U473 ( .A(n594), .B(n591), .Z(n593) );
  XNOR U474 ( .A(n407), .B(n587), .Z(n589) );
  XOR U475 ( .A(n595), .B(n596), .Z(n407) );
  AND U476 ( .A(n284), .B(n597), .Z(n596) );
  XOR U477 ( .A(n598), .B(n595), .Z(n597) );
  XOR U478 ( .A(n599), .B(n600), .Z(n587) );
  AND U479 ( .A(n601), .B(n602), .Z(n600) );
  XOR U480 ( .A(n599), .B(n422), .Z(n602) );
  XOR U481 ( .A(n603), .B(n604), .Z(n422) );
  AND U482 ( .A(n286), .B(n605), .Z(n604) );
  XOR U483 ( .A(n606), .B(n603), .Z(n605) );
  XNOR U484 ( .A(n419), .B(n599), .Z(n601) );
  XOR U485 ( .A(n607), .B(n608), .Z(n419) );
  AND U486 ( .A(n284), .B(n609), .Z(n608) );
  XOR U487 ( .A(n610), .B(n607), .Z(n609) );
  XOR U488 ( .A(n611), .B(n612), .Z(n599) );
  AND U489 ( .A(n613), .B(n614), .Z(n612) );
  XOR U490 ( .A(n611), .B(n434), .Z(n614) );
  XOR U491 ( .A(n615), .B(n616), .Z(n434) );
  AND U492 ( .A(n286), .B(n617), .Z(n616) );
  XOR U493 ( .A(n618), .B(n615), .Z(n617) );
  XNOR U494 ( .A(n431), .B(n611), .Z(n613) );
  XOR U495 ( .A(n619), .B(n620), .Z(n431) );
  AND U496 ( .A(n284), .B(n621), .Z(n620) );
  XOR U497 ( .A(n622), .B(n619), .Z(n621) );
  XOR U498 ( .A(n623), .B(n624), .Z(n611) );
  AND U499 ( .A(n625), .B(n626), .Z(n624) );
  XOR U500 ( .A(n623), .B(n446), .Z(n626) );
  XOR U501 ( .A(n627), .B(n628), .Z(n446) );
  AND U502 ( .A(n286), .B(n629), .Z(n628) );
  XOR U503 ( .A(n630), .B(n627), .Z(n629) );
  XNOR U504 ( .A(n443), .B(n623), .Z(n625) );
  XOR U505 ( .A(n631), .B(n632), .Z(n443) );
  AND U506 ( .A(n284), .B(n633), .Z(n632) );
  XOR U507 ( .A(n634), .B(n631), .Z(n633) );
  XOR U508 ( .A(n635), .B(n636), .Z(n623) );
  AND U509 ( .A(n637), .B(n638), .Z(n636) );
  XOR U510 ( .A(n458), .B(n635), .Z(n638) );
  XOR U511 ( .A(n639), .B(n640), .Z(n458) );
  AND U512 ( .A(n286), .B(n641), .Z(n640) );
  XOR U513 ( .A(n639), .B(n642), .Z(n641) );
  XNOR U514 ( .A(n635), .B(n455), .Z(n637) );
  XOR U515 ( .A(n643), .B(n644), .Z(n455) );
  AND U516 ( .A(n284), .B(n645), .Z(n644) );
  XOR U517 ( .A(n643), .B(n646), .Z(n645) );
  XOR U518 ( .A(n647), .B(n648), .Z(n635) );
  AND U519 ( .A(n649), .B(n650), .Z(n648) );
  XOR U520 ( .A(n647), .B(n470), .Z(n650) );
  XOR U521 ( .A(n651), .B(n652), .Z(n470) );
  AND U522 ( .A(n286), .B(n653), .Z(n652) );
  XOR U523 ( .A(n654), .B(n651), .Z(n653) );
  XNOR U524 ( .A(n467), .B(n647), .Z(n649) );
  XOR U525 ( .A(n655), .B(n656), .Z(n467) );
  AND U526 ( .A(n284), .B(n657), .Z(n656) );
  XOR U527 ( .A(n658), .B(n655), .Z(n657) );
  XOR U528 ( .A(n659), .B(n660), .Z(n647) );
  AND U529 ( .A(n661), .B(n662), .Z(n660) );
  XNOR U530 ( .A(n663), .B(n482), .Z(n662) );
  XOR U531 ( .A(n664), .B(n665), .Z(n482) );
  AND U532 ( .A(n286), .B(n666), .Z(n665) );
  XOR U533 ( .A(n667), .B(n664), .Z(n666) );
  XNOR U534 ( .A(n479), .B(n659), .Z(n661) );
  XOR U535 ( .A(n668), .B(n669), .Z(n479) );
  AND U536 ( .A(n284), .B(n670), .Z(n669) );
  XOR U537 ( .A(n671), .B(n668), .Z(n670) );
  IV U538 ( .A(n663), .Z(n659) );
  AND U539 ( .A(n487), .B(n490), .Z(n663) );
  XNOR U540 ( .A(n672), .B(n673), .Z(n490) );
  AND U541 ( .A(n286), .B(n674), .Z(n673) );
  XNOR U542 ( .A(n675), .B(n672), .Z(n674) );
  XOR U543 ( .A(n676), .B(n677), .Z(n286) );
  AND U544 ( .A(n678), .B(n679), .Z(n677) );
  XOR U545 ( .A(n498), .B(n676), .Z(n679) );
  IV U546 ( .A(n680), .Z(n498) );
  AND U547 ( .A(n681), .B(n682), .Z(n680) );
  XOR U548 ( .A(n676), .B(n495), .Z(n678) );
  AND U549 ( .A(n683), .B(n684), .Z(n495) );
  XOR U550 ( .A(n685), .B(n686), .Z(n676) );
  AND U551 ( .A(n687), .B(n688), .Z(n686) );
  XOR U552 ( .A(n685), .B(n510), .Z(n688) );
  XOR U553 ( .A(n689), .B(n690), .Z(n510) );
  AND U554 ( .A(n246), .B(n691), .Z(n690) );
  XOR U555 ( .A(n692), .B(n689), .Z(n691) );
  XNOR U556 ( .A(n507), .B(n685), .Z(n687) );
  XOR U557 ( .A(n693), .B(n694), .Z(n507) );
  AND U558 ( .A(n244), .B(n695), .Z(n694) );
  XOR U559 ( .A(n696), .B(n693), .Z(n695) );
  XOR U560 ( .A(n697), .B(n698), .Z(n685) );
  AND U561 ( .A(n699), .B(n700), .Z(n698) );
  XOR U562 ( .A(n697), .B(n522), .Z(n700) );
  XOR U563 ( .A(n701), .B(n702), .Z(n522) );
  AND U564 ( .A(n246), .B(n703), .Z(n702) );
  XOR U565 ( .A(n704), .B(n701), .Z(n703) );
  XNOR U566 ( .A(n519), .B(n697), .Z(n699) );
  XOR U567 ( .A(n705), .B(n706), .Z(n519) );
  AND U568 ( .A(n244), .B(n707), .Z(n706) );
  XOR U569 ( .A(n708), .B(n705), .Z(n707) );
  XOR U570 ( .A(n709), .B(n710), .Z(n697) );
  AND U571 ( .A(n711), .B(n712), .Z(n710) );
  XOR U572 ( .A(n709), .B(n534), .Z(n712) );
  XOR U573 ( .A(n713), .B(n714), .Z(n534) );
  AND U574 ( .A(n246), .B(n715), .Z(n714) );
  XOR U575 ( .A(n716), .B(n713), .Z(n715) );
  XNOR U576 ( .A(n531), .B(n709), .Z(n711) );
  XOR U577 ( .A(n717), .B(n718), .Z(n531) );
  AND U578 ( .A(n244), .B(n719), .Z(n718) );
  XOR U579 ( .A(n720), .B(n717), .Z(n719) );
  XOR U580 ( .A(n721), .B(n722), .Z(n709) );
  AND U581 ( .A(n723), .B(n724), .Z(n722) );
  XOR U582 ( .A(n721), .B(n546), .Z(n724) );
  XOR U583 ( .A(n725), .B(n726), .Z(n546) );
  AND U584 ( .A(n246), .B(n727), .Z(n726) );
  XOR U585 ( .A(n728), .B(n725), .Z(n727) );
  XNOR U586 ( .A(n543), .B(n721), .Z(n723) );
  XOR U587 ( .A(n729), .B(n730), .Z(n543) );
  AND U588 ( .A(n244), .B(n731), .Z(n730) );
  XOR U589 ( .A(n732), .B(n729), .Z(n731) );
  XOR U590 ( .A(n733), .B(n734), .Z(n721) );
  AND U591 ( .A(n735), .B(n736), .Z(n734) );
  XOR U592 ( .A(n733), .B(n558), .Z(n736) );
  XOR U593 ( .A(n737), .B(n738), .Z(n558) );
  AND U594 ( .A(n246), .B(n739), .Z(n738) );
  XOR U595 ( .A(n740), .B(n737), .Z(n739) );
  XNOR U596 ( .A(n555), .B(n733), .Z(n735) );
  XOR U597 ( .A(n741), .B(n742), .Z(n555) );
  AND U598 ( .A(n244), .B(n743), .Z(n742) );
  XOR U599 ( .A(n744), .B(n741), .Z(n743) );
  XOR U600 ( .A(n745), .B(n746), .Z(n733) );
  AND U601 ( .A(n747), .B(n748), .Z(n746) );
  XOR U602 ( .A(n745), .B(n570), .Z(n748) );
  XOR U603 ( .A(n749), .B(n750), .Z(n570) );
  AND U604 ( .A(n246), .B(n751), .Z(n750) );
  XOR U605 ( .A(n752), .B(n749), .Z(n751) );
  XNOR U606 ( .A(n567), .B(n745), .Z(n747) );
  XOR U607 ( .A(n753), .B(n754), .Z(n567) );
  AND U608 ( .A(n244), .B(n755), .Z(n754) );
  XOR U609 ( .A(n756), .B(n753), .Z(n755) );
  XOR U610 ( .A(n757), .B(n758), .Z(n745) );
  AND U611 ( .A(n759), .B(n760), .Z(n758) );
  XOR U612 ( .A(n757), .B(n582), .Z(n760) );
  XOR U613 ( .A(n761), .B(n762), .Z(n582) );
  AND U614 ( .A(n246), .B(n763), .Z(n762) );
  XOR U615 ( .A(n764), .B(n761), .Z(n763) );
  XNOR U616 ( .A(n579), .B(n757), .Z(n759) );
  XOR U617 ( .A(n765), .B(n766), .Z(n579) );
  AND U618 ( .A(n244), .B(n767), .Z(n766) );
  XOR U619 ( .A(n768), .B(n765), .Z(n767) );
  XOR U620 ( .A(n769), .B(n770), .Z(n757) );
  AND U621 ( .A(n771), .B(n772), .Z(n770) );
  XOR U622 ( .A(n769), .B(n594), .Z(n772) );
  XOR U623 ( .A(n773), .B(n774), .Z(n594) );
  AND U624 ( .A(n246), .B(n775), .Z(n774) );
  XOR U625 ( .A(n776), .B(n773), .Z(n775) );
  XNOR U626 ( .A(n591), .B(n769), .Z(n771) );
  XOR U627 ( .A(n777), .B(n778), .Z(n591) );
  AND U628 ( .A(n244), .B(n779), .Z(n778) );
  XOR U629 ( .A(n780), .B(n777), .Z(n779) );
  XOR U630 ( .A(n781), .B(n782), .Z(n769) );
  AND U631 ( .A(n783), .B(n784), .Z(n782) );
  XOR U632 ( .A(n781), .B(n606), .Z(n784) );
  XOR U633 ( .A(n785), .B(n786), .Z(n606) );
  AND U634 ( .A(n246), .B(n787), .Z(n786) );
  XOR U635 ( .A(n788), .B(n785), .Z(n787) );
  XNOR U636 ( .A(n603), .B(n781), .Z(n783) );
  XOR U637 ( .A(n789), .B(n790), .Z(n603) );
  AND U638 ( .A(n244), .B(n791), .Z(n790) );
  XOR U639 ( .A(n792), .B(n789), .Z(n791) );
  XOR U640 ( .A(n793), .B(n794), .Z(n781) );
  AND U641 ( .A(n795), .B(n796), .Z(n794) );
  XOR U642 ( .A(n793), .B(n618), .Z(n796) );
  XOR U643 ( .A(n797), .B(n798), .Z(n618) );
  AND U644 ( .A(n246), .B(n799), .Z(n798) );
  XOR U645 ( .A(n800), .B(n797), .Z(n799) );
  XNOR U646 ( .A(n615), .B(n793), .Z(n795) );
  XOR U647 ( .A(n801), .B(n802), .Z(n615) );
  AND U648 ( .A(n244), .B(n803), .Z(n802) );
  XOR U649 ( .A(n804), .B(n801), .Z(n803) );
  XOR U650 ( .A(n805), .B(n806), .Z(n793) );
  AND U651 ( .A(n807), .B(n808), .Z(n806) );
  XOR U652 ( .A(n805), .B(n630), .Z(n808) );
  XOR U653 ( .A(n809), .B(n810), .Z(n630) );
  AND U654 ( .A(n246), .B(n811), .Z(n810) );
  XOR U655 ( .A(n812), .B(n809), .Z(n811) );
  XNOR U656 ( .A(n627), .B(n805), .Z(n807) );
  XOR U657 ( .A(n813), .B(n814), .Z(n627) );
  AND U658 ( .A(n244), .B(n815), .Z(n814) );
  XOR U659 ( .A(n816), .B(n813), .Z(n815) );
  XOR U660 ( .A(n817), .B(n818), .Z(n805) );
  AND U661 ( .A(n819), .B(n820), .Z(n818) );
  XOR U662 ( .A(n642), .B(n817), .Z(n820) );
  XOR U663 ( .A(n821), .B(n822), .Z(n642) );
  AND U664 ( .A(n246), .B(n823), .Z(n822) );
  XOR U665 ( .A(n821), .B(n824), .Z(n823) );
  XNOR U666 ( .A(n817), .B(n639), .Z(n819) );
  XOR U667 ( .A(n825), .B(n826), .Z(n639) );
  AND U668 ( .A(n244), .B(n827), .Z(n826) );
  XOR U669 ( .A(n825), .B(n828), .Z(n827) );
  XOR U670 ( .A(n829), .B(n830), .Z(n817) );
  AND U671 ( .A(n831), .B(n832), .Z(n830) );
  XOR U672 ( .A(n829), .B(n654), .Z(n832) );
  XOR U673 ( .A(n833), .B(n834), .Z(n654) );
  AND U674 ( .A(n246), .B(n835), .Z(n834) );
  XOR U675 ( .A(n836), .B(n833), .Z(n835) );
  XNOR U676 ( .A(n651), .B(n829), .Z(n831) );
  XOR U677 ( .A(n837), .B(n838), .Z(n651) );
  AND U678 ( .A(n244), .B(n839), .Z(n838) );
  XOR U679 ( .A(n840), .B(n837), .Z(n839) );
  XOR U680 ( .A(n841), .B(n842), .Z(n829) );
  AND U681 ( .A(n843), .B(n844), .Z(n842) );
  XNOR U682 ( .A(n845), .B(n667), .Z(n844) );
  XOR U683 ( .A(n846), .B(n847), .Z(n667) );
  AND U684 ( .A(n246), .B(n848), .Z(n847) );
  XOR U685 ( .A(n849), .B(n846), .Z(n848) );
  XNOR U686 ( .A(n664), .B(n841), .Z(n843) );
  XOR U687 ( .A(n850), .B(n851), .Z(n664) );
  AND U688 ( .A(n244), .B(n852), .Z(n851) );
  XOR U689 ( .A(n853), .B(n850), .Z(n852) );
  IV U690 ( .A(n845), .Z(n841) );
  AND U691 ( .A(n672), .B(n675), .Z(n845) );
  XNOR U692 ( .A(n854), .B(n855), .Z(n675) );
  AND U693 ( .A(n246), .B(n856), .Z(n855) );
  XNOR U694 ( .A(n857), .B(n854), .Z(n856) );
  XOR U695 ( .A(n858), .B(n859), .Z(n246) );
  AND U696 ( .A(n860), .B(n861), .Z(n859) );
  XNOR U697 ( .A(n681), .B(n858), .Z(n861) );
  AND U698 ( .A(n862), .B(n863), .Z(n681) );
  XOR U699 ( .A(n858), .B(n682), .Z(n860) );
  AND U700 ( .A(n864), .B(n865), .Z(n682) );
  XOR U701 ( .A(n866), .B(n867), .Z(n858) );
  AND U702 ( .A(n868), .B(n869), .Z(n867) );
  XOR U703 ( .A(n866), .B(n692), .Z(n869) );
  XOR U704 ( .A(n870), .B(n871), .Z(n692) );
  AND U705 ( .A(n158), .B(n872), .Z(n871) );
  XOR U706 ( .A(n873), .B(n870), .Z(n872) );
  XNOR U707 ( .A(n689), .B(n866), .Z(n868) );
  XOR U708 ( .A(n874), .B(n875), .Z(n689) );
  AND U709 ( .A(n156), .B(n876), .Z(n875) );
  XOR U710 ( .A(n877), .B(n874), .Z(n876) );
  XOR U711 ( .A(n878), .B(n879), .Z(n866) );
  AND U712 ( .A(n880), .B(n881), .Z(n879) );
  XOR U713 ( .A(n878), .B(n704), .Z(n881) );
  XOR U714 ( .A(n882), .B(n883), .Z(n704) );
  AND U715 ( .A(n158), .B(n884), .Z(n883) );
  XOR U716 ( .A(n885), .B(n882), .Z(n884) );
  XNOR U717 ( .A(n701), .B(n878), .Z(n880) );
  XOR U718 ( .A(n886), .B(n887), .Z(n701) );
  AND U719 ( .A(n156), .B(n888), .Z(n887) );
  XOR U720 ( .A(n889), .B(n886), .Z(n888) );
  XOR U721 ( .A(n890), .B(n891), .Z(n878) );
  AND U722 ( .A(n892), .B(n893), .Z(n891) );
  XOR U723 ( .A(n890), .B(n716), .Z(n893) );
  XOR U724 ( .A(n894), .B(n895), .Z(n716) );
  AND U725 ( .A(n158), .B(n896), .Z(n895) );
  XOR U726 ( .A(n897), .B(n894), .Z(n896) );
  XNOR U727 ( .A(n713), .B(n890), .Z(n892) );
  XOR U728 ( .A(n898), .B(n899), .Z(n713) );
  AND U729 ( .A(n156), .B(n900), .Z(n899) );
  XOR U730 ( .A(n901), .B(n898), .Z(n900) );
  XOR U731 ( .A(n902), .B(n903), .Z(n890) );
  AND U732 ( .A(n904), .B(n905), .Z(n903) );
  XOR U733 ( .A(n902), .B(n728), .Z(n905) );
  XOR U734 ( .A(n906), .B(n907), .Z(n728) );
  AND U735 ( .A(n158), .B(n908), .Z(n907) );
  XOR U736 ( .A(n909), .B(n906), .Z(n908) );
  XNOR U737 ( .A(n725), .B(n902), .Z(n904) );
  XOR U738 ( .A(n910), .B(n911), .Z(n725) );
  AND U739 ( .A(n156), .B(n912), .Z(n911) );
  XOR U740 ( .A(n913), .B(n910), .Z(n912) );
  XOR U741 ( .A(n914), .B(n915), .Z(n902) );
  AND U742 ( .A(n916), .B(n917), .Z(n915) );
  XOR U743 ( .A(n914), .B(n740), .Z(n917) );
  XOR U744 ( .A(n918), .B(n919), .Z(n740) );
  AND U745 ( .A(n158), .B(n920), .Z(n919) );
  XOR U746 ( .A(n921), .B(n918), .Z(n920) );
  XNOR U747 ( .A(n737), .B(n914), .Z(n916) );
  XOR U748 ( .A(n922), .B(n923), .Z(n737) );
  AND U749 ( .A(n156), .B(n924), .Z(n923) );
  XOR U750 ( .A(n925), .B(n922), .Z(n924) );
  XOR U751 ( .A(n926), .B(n927), .Z(n914) );
  AND U752 ( .A(n928), .B(n929), .Z(n927) );
  XOR U753 ( .A(n926), .B(n752), .Z(n929) );
  XOR U754 ( .A(n930), .B(n931), .Z(n752) );
  AND U755 ( .A(n158), .B(n932), .Z(n931) );
  XOR U756 ( .A(n933), .B(n930), .Z(n932) );
  XNOR U757 ( .A(n749), .B(n926), .Z(n928) );
  XOR U758 ( .A(n934), .B(n935), .Z(n749) );
  AND U759 ( .A(n156), .B(n936), .Z(n935) );
  XOR U760 ( .A(n937), .B(n934), .Z(n936) );
  XOR U761 ( .A(n938), .B(n939), .Z(n926) );
  AND U762 ( .A(n940), .B(n941), .Z(n939) );
  XOR U763 ( .A(n938), .B(n764), .Z(n941) );
  XOR U764 ( .A(n942), .B(n943), .Z(n764) );
  AND U765 ( .A(n158), .B(n944), .Z(n943) );
  XOR U766 ( .A(n945), .B(n942), .Z(n944) );
  XNOR U767 ( .A(n761), .B(n938), .Z(n940) );
  XOR U768 ( .A(n946), .B(n947), .Z(n761) );
  AND U769 ( .A(n156), .B(n948), .Z(n947) );
  XOR U770 ( .A(n949), .B(n946), .Z(n948) );
  XOR U771 ( .A(n950), .B(n951), .Z(n938) );
  AND U772 ( .A(n952), .B(n953), .Z(n951) );
  XOR U773 ( .A(n950), .B(n776), .Z(n953) );
  XOR U774 ( .A(n954), .B(n955), .Z(n776) );
  AND U775 ( .A(n158), .B(n956), .Z(n955) );
  XOR U776 ( .A(n957), .B(n954), .Z(n956) );
  XNOR U777 ( .A(n773), .B(n950), .Z(n952) );
  XOR U778 ( .A(n958), .B(n959), .Z(n773) );
  AND U779 ( .A(n156), .B(n960), .Z(n959) );
  XOR U780 ( .A(n961), .B(n958), .Z(n960) );
  XOR U781 ( .A(n962), .B(n963), .Z(n950) );
  AND U782 ( .A(n964), .B(n965), .Z(n963) );
  XOR U783 ( .A(n962), .B(n788), .Z(n965) );
  XOR U784 ( .A(n966), .B(n967), .Z(n788) );
  AND U785 ( .A(n158), .B(n968), .Z(n967) );
  XOR U786 ( .A(n969), .B(n966), .Z(n968) );
  XNOR U787 ( .A(n785), .B(n962), .Z(n964) );
  XOR U788 ( .A(n970), .B(n971), .Z(n785) );
  AND U789 ( .A(n156), .B(n972), .Z(n971) );
  XOR U790 ( .A(n973), .B(n970), .Z(n972) );
  XOR U791 ( .A(n974), .B(n975), .Z(n962) );
  AND U792 ( .A(n976), .B(n977), .Z(n975) );
  XOR U793 ( .A(n974), .B(n800), .Z(n977) );
  XOR U794 ( .A(n978), .B(n979), .Z(n800) );
  AND U795 ( .A(n158), .B(n980), .Z(n979) );
  XOR U796 ( .A(n981), .B(n978), .Z(n980) );
  XNOR U797 ( .A(n797), .B(n974), .Z(n976) );
  XOR U798 ( .A(n982), .B(n983), .Z(n797) );
  AND U799 ( .A(n156), .B(n984), .Z(n983) );
  XOR U800 ( .A(n985), .B(n982), .Z(n984) );
  XOR U801 ( .A(n986), .B(n987), .Z(n974) );
  AND U802 ( .A(n988), .B(n989), .Z(n987) );
  XOR U803 ( .A(n986), .B(n812), .Z(n989) );
  XOR U804 ( .A(n990), .B(n991), .Z(n812) );
  AND U805 ( .A(n158), .B(n992), .Z(n991) );
  XOR U806 ( .A(n993), .B(n990), .Z(n992) );
  XNOR U807 ( .A(n809), .B(n986), .Z(n988) );
  XOR U808 ( .A(n994), .B(n995), .Z(n809) );
  AND U809 ( .A(n156), .B(n996), .Z(n995) );
  XOR U810 ( .A(n997), .B(n994), .Z(n996) );
  XOR U811 ( .A(n998), .B(n999), .Z(n986) );
  AND U812 ( .A(n1000), .B(n1001), .Z(n999) );
  XOR U813 ( .A(n824), .B(n998), .Z(n1001) );
  XOR U814 ( .A(n1002), .B(n1003), .Z(n824) );
  AND U815 ( .A(n158), .B(n1004), .Z(n1003) );
  XOR U816 ( .A(n1002), .B(n1005), .Z(n1004) );
  XNOR U817 ( .A(n998), .B(n821), .Z(n1000) );
  XOR U818 ( .A(n1006), .B(n1007), .Z(n821) );
  AND U819 ( .A(n156), .B(n1008), .Z(n1007) );
  XOR U820 ( .A(n1006), .B(n1009), .Z(n1008) );
  XOR U821 ( .A(n1010), .B(n1011), .Z(n998) );
  AND U822 ( .A(n1012), .B(n1013), .Z(n1011) );
  XOR U823 ( .A(n1010), .B(n836), .Z(n1013) );
  XOR U824 ( .A(n1014), .B(n1015), .Z(n836) );
  AND U825 ( .A(n158), .B(n1016), .Z(n1015) );
  XOR U826 ( .A(n1017), .B(n1014), .Z(n1016) );
  XNOR U827 ( .A(n833), .B(n1010), .Z(n1012) );
  XOR U828 ( .A(n1018), .B(n1019), .Z(n833) );
  AND U829 ( .A(n156), .B(n1020), .Z(n1019) );
  XOR U830 ( .A(n1021), .B(n1018), .Z(n1020) );
  XOR U831 ( .A(n1022), .B(n1023), .Z(n1010) );
  AND U832 ( .A(n1024), .B(n1025), .Z(n1023) );
  XNOR U833 ( .A(n1026), .B(n849), .Z(n1025) );
  XOR U834 ( .A(n1027), .B(n1028), .Z(n849) );
  AND U835 ( .A(n158), .B(n1029), .Z(n1028) );
  XOR U836 ( .A(n1030), .B(n1027), .Z(n1029) );
  XNOR U837 ( .A(n846), .B(n1022), .Z(n1024) );
  XOR U838 ( .A(n1031), .B(n1032), .Z(n846) );
  AND U839 ( .A(n156), .B(n1033), .Z(n1032) );
  XOR U840 ( .A(n1034), .B(n1031), .Z(n1033) );
  IV U841 ( .A(n1026), .Z(n1022) );
  AND U842 ( .A(n854), .B(n857), .Z(n1026) );
  XNOR U843 ( .A(n1035), .B(n1036), .Z(n857) );
  AND U844 ( .A(n158), .B(n1037), .Z(n1036) );
  XNOR U845 ( .A(n1038), .B(n1035), .Z(n1037) );
  XOR U846 ( .A(n1039), .B(n1040), .Z(n158) );
  AND U847 ( .A(n1041), .B(n1042), .Z(n1040) );
  XNOR U848 ( .A(n862), .B(n1039), .Z(n1042) );
  AND U849 ( .A(p_input[1023]), .B(p_input[1007]), .Z(n862) );
  XOR U850 ( .A(n1039), .B(n863), .Z(n1041) );
  AND U851 ( .A(p_input[991]), .B(p_input[975]), .Z(n863) );
  XOR U852 ( .A(n1043), .B(n1044), .Z(n1039) );
  AND U853 ( .A(n1045), .B(n1046), .Z(n1044) );
  XOR U854 ( .A(n1043), .B(n873), .Z(n1046) );
  XNOR U855 ( .A(p_input[1006]), .B(n1047), .Z(n873) );
  AND U856 ( .A(n98), .B(n1048), .Z(n1047) );
  XOR U857 ( .A(p_input[1022]), .B(p_input[1006]), .Z(n1048) );
  XNOR U858 ( .A(n870), .B(n1043), .Z(n1045) );
  XOR U859 ( .A(n1049), .B(n1050), .Z(n870) );
  AND U860 ( .A(n96), .B(n1051), .Z(n1050) );
  XOR U861 ( .A(p_input[990]), .B(p_input[974]), .Z(n1051) );
  XOR U862 ( .A(n1052), .B(n1053), .Z(n1043) );
  AND U863 ( .A(n1054), .B(n1055), .Z(n1053) );
  XOR U864 ( .A(n1052), .B(n885), .Z(n1055) );
  XNOR U865 ( .A(p_input[1005]), .B(n1056), .Z(n885) );
  AND U866 ( .A(n98), .B(n1057), .Z(n1056) );
  XOR U867 ( .A(p_input[1021]), .B(p_input[1005]), .Z(n1057) );
  XNOR U868 ( .A(n882), .B(n1052), .Z(n1054) );
  XOR U869 ( .A(n1058), .B(n1059), .Z(n882) );
  AND U870 ( .A(n96), .B(n1060), .Z(n1059) );
  XOR U871 ( .A(p_input[989]), .B(p_input[973]), .Z(n1060) );
  XOR U872 ( .A(n1061), .B(n1062), .Z(n1052) );
  AND U873 ( .A(n1063), .B(n1064), .Z(n1062) );
  XOR U874 ( .A(n1061), .B(n897), .Z(n1064) );
  XNOR U875 ( .A(p_input[1004]), .B(n1065), .Z(n897) );
  AND U876 ( .A(n98), .B(n1066), .Z(n1065) );
  XOR U877 ( .A(p_input[1020]), .B(p_input[1004]), .Z(n1066) );
  XNOR U878 ( .A(n894), .B(n1061), .Z(n1063) );
  XOR U879 ( .A(n1067), .B(n1068), .Z(n894) );
  AND U880 ( .A(n96), .B(n1069), .Z(n1068) );
  XOR U881 ( .A(p_input[988]), .B(p_input[972]), .Z(n1069) );
  XOR U882 ( .A(n1070), .B(n1071), .Z(n1061) );
  AND U883 ( .A(n1072), .B(n1073), .Z(n1071) );
  XOR U884 ( .A(n1070), .B(n909), .Z(n1073) );
  XNOR U885 ( .A(p_input[1003]), .B(n1074), .Z(n909) );
  AND U886 ( .A(n98), .B(n1075), .Z(n1074) );
  XOR U887 ( .A(p_input[1019]), .B(p_input[1003]), .Z(n1075) );
  XNOR U888 ( .A(n906), .B(n1070), .Z(n1072) );
  XOR U889 ( .A(n1076), .B(n1077), .Z(n906) );
  AND U890 ( .A(n96), .B(n1078), .Z(n1077) );
  XOR U891 ( .A(p_input[987]), .B(p_input[971]), .Z(n1078) );
  XOR U892 ( .A(n1079), .B(n1080), .Z(n1070) );
  AND U893 ( .A(n1081), .B(n1082), .Z(n1080) );
  XOR U894 ( .A(n1079), .B(n921), .Z(n1082) );
  XNOR U895 ( .A(p_input[1002]), .B(n1083), .Z(n921) );
  AND U896 ( .A(n98), .B(n1084), .Z(n1083) );
  XOR U897 ( .A(p_input[1018]), .B(p_input[1002]), .Z(n1084) );
  XNOR U898 ( .A(n918), .B(n1079), .Z(n1081) );
  XOR U899 ( .A(n1085), .B(n1086), .Z(n918) );
  AND U900 ( .A(n96), .B(n1087), .Z(n1086) );
  XOR U901 ( .A(p_input[986]), .B(p_input[970]), .Z(n1087) );
  XOR U902 ( .A(n1088), .B(n1089), .Z(n1079) );
  AND U903 ( .A(n1090), .B(n1091), .Z(n1089) );
  XOR U904 ( .A(n1088), .B(n933), .Z(n1091) );
  XNOR U905 ( .A(p_input[1001]), .B(n1092), .Z(n933) );
  AND U906 ( .A(n98), .B(n1093), .Z(n1092) );
  XOR U907 ( .A(p_input[1017]), .B(p_input[1001]), .Z(n1093) );
  XNOR U908 ( .A(n930), .B(n1088), .Z(n1090) );
  XOR U909 ( .A(n1094), .B(n1095), .Z(n930) );
  AND U910 ( .A(n96), .B(n1096), .Z(n1095) );
  XOR U911 ( .A(p_input[985]), .B(p_input[969]), .Z(n1096) );
  XOR U912 ( .A(n1097), .B(n1098), .Z(n1088) );
  AND U913 ( .A(n1099), .B(n1100), .Z(n1098) );
  XOR U914 ( .A(n1097), .B(n945), .Z(n1100) );
  XNOR U915 ( .A(p_input[1000]), .B(n1101), .Z(n945) );
  AND U916 ( .A(n98), .B(n1102), .Z(n1101) );
  XOR U917 ( .A(p_input[1016]), .B(p_input[1000]), .Z(n1102) );
  XNOR U918 ( .A(n942), .B(n1097), .Z(n1099) );
  XOR U919 ( .A(n1103), .B(n1104), .Z(n942) );
  AND U920 ( .A(n96), .B(n1105), .Z(n1104) );
  XOR U921 ( .A(p_input[984]), .B(p_input[968]), .Z(n1105) );
  XOR U922 ( .A(n1106), .B(n1107), .Z(n1097) );
  AND U923 ( .A(n1108), .B(n1109), .Z(n1107) );
  XOR U924 ( .A(n1106), .B(n957), .Z(n1109) );
  XNOR U925 ( .A(p_input[999]), .B(n1110), .Z(n957) );
  AND U926 ( .A(n98), .B(n1111), .Z(n1110) );
  XOR U927 ( .A(p_input[999]), .B(p_input[1015]), .Z(n1111) );
  XNOR U928 ( .A(n954), .B(n1106), .Z(n1108) );
  XOR U929 ( .A(n1112), .B(n1113), .Z(n954) );
  AND U930 ( .A(n96), .B(n1114), .Z(n1113) );
  XOR U931 ( .A(p_input[983]), .B(p_input[967]), .Z(n1114) );
  XOR U932 ( .A(n1115), .B(n1116), .Z(n1106) );
  AND U933 ( .A(n1117), .B(n1118), .Z(n1116) );
  XOR U934 ( .A(n1115), .B(n969), .Z(n1118) );
  XNOR U935 ( .A(p_input[998]), .B(n1119), .Z(n969) );
  AND U936 ( .A(n98), .B(n1120), .Z(n1119) );
  XOR U937 ( .A(p_input[998]), .B(p_input[1014]), .Z(n1120) );
  XNOR U938 ( .A(n966), .B(n1115), .Z(n1117) );
  XOR U939 ( .A(n1121), .B(n1122), .Z(n966) );
  AND U940 ( .A(n96), .B(n1123), .Z(n1122) );
  XOR U941 ( .A(p_input[982]), .B(p_input[966]), .Z(n1123) );
  XOR U942 ( .A(n1124), .B(n1125), .Z(n1115) );
  AND U943 ( .A(n1126), .B(n1127), .Z(n1125) );
  XOR U944 ( .A(n1124), .B(n981), .Z(n1127) );
  XNOR U945 ( .A(p_input[997]), .B(n1128), .Z(n981) );
  AND U946 ( .A(n98), .B(n1129), .Z(n1128) );
  XOR U947 ( .A(p_input[997]), .B(p_input[1013]), .Z(n1129) );
  XNOR U948 ( .A(n978), .B(n1124), .Z(n1126) );
  XOR U949 ( .A(n1130), .B(n1131), .Z(n978) );
  AND U950 ( .A(n96), .B(n1132), .Z(n1131) );
  XOR U951 ( .A(p_input[981]), .B(p_input[965]), .Z(n1132) );
  XOR U952 ( .A(n1133), .B(n1134), .Z(n1124) );
  AND U953 ( .A(n1135), .B(n1136), .Z(n1134) );
  XOR U954 ( .A(n1133), .B(n993), .Z(n1136) );
  XNOR U955 ( .A(p_input[996]), .B(n1137), .Z(n993) );
  AND U956 ( .A(n98), .B(n1138), .Z(n1137) );
  XOR U957 ( .A(p_input[996]), .B(p_input[1012]), .Z(n1138) );
  XNOR U958 ( .A(n990), .B(n1133), .Z(n1135) );
  XOR U959 ( .A(n1139), .B(n1140), .Z(n990) );
  AND U960 ( .A(n96), .B(n1141), .Z(n1140) );
  XOR U961 ( .A(p_input[980]), .B(p_input[964]), .Z(n1141) );
  XOR U962 ( .A(n1142), .B(n1143), .Z(n1133) );
  AND U963 ( .A(n1144), .B(n1145), .Z(n1143) );
  XOR U964 ( .A(n1005), .B(n1142), .Z(n1145) );
  XNOR U965 ( .A(p_input[995]), .B(n1146), .Z(n1005) );
  AND U966 ( .A(n98), .B(n1147), .Z(n1146) );
  XOR U967 ( .A(p_input[995]), .B(p_input[1011]), .Z(n1147) );
  XNOR U968 ( .A(n1142), .B(n1002), .Z(n1144) );
  XOR U969 ( .A(n1148), .B(n1149), .Z(n1002) );
  AND U970 ( .A(n96), .B(n1150), .Z(n1149) );
  XOR U971 ( .A(p_input[979]), .B(p_input[963]), .Z(n1150) );
  XOR U972 ( .A(n1151), .B(n1152), .Z(n1142) );
  AND U973 ( .A(n1153), .B(n1154), .Z(n1152) );
  XOR U974 ( .A(n1151), .B(n1017), .Z(n1154) );
  XNOR U975 ( .A(p_input[994]), .B(n1155), .Z(n1017) );
  AND U976 ( .A(n98), .B(n1156), .Z(n1155) );
  XOR U977 ( .A(p_input[994]), .B(p_input[1010]), .Z(n1156) );
  XNOR U978 ( .A(n1014), .B(n1151), .Z(n1153) );
  XOR U979 ( .A(n1157), .B(n1158), .Z(n1014) );
  AND U980 ( .A(n96), .B(n1159), .Z(n1158) );
  XOR U981 ( .A(p_input[978]), .B(p_input[962]), .Z(n1159) );
  XOR U982 ( .A(n1160), .B(n1161), .Z(n1151) );
  AND U983 ( .A(n1162), .B(n1163), .Z(n1161) );
  XNOR U984 ( .A(n1164), .B(n1030), .Z(n1163) );
  XNOR U985 ( .A(p_input[993]), .B(n1165), .Z(n1030) );
  AND U986 ( .A(n98), .B(n1166), .Z(n1165) );
  XNOR U987 ( .A(n1167), .B(p_input[1009]), .Z(n1166) );
  IV U988 ( .A(p_input[993]), .Z(n1167) );
  XNOR U989 ( .A(n1027), .B(n1160), .Z(n1162) );
  XNOR U990 ( .A(p_input[961]), .B(n1168), .Z(n1027) );
  AND U991 ( .A(n96), .B(n1169), .Z(n1168) );
  XOR U992 ( .A(p_input[977]), .B(p_input[961]), .Z(n1169) );
  IV U993 ( .A(n1164), .Z(n1160) );
  AND U994 ( .A(n1035), .B(n1038), .Z(n1164) );
  XOR U995 ( .A(p_input[992]), .B(n1170), .Z(n1038) );
  AND U996 ( .A(n98), .B(n1171), .Z(n1170) );
  XOR U997 ( .A(p_input[992]), .B(p_input[1008]), .Z(n1171) );
  XOR U998 ( .A(n1172), .B(n1173), .Z(n98) );
  AND U999 ( .A(n1174), .B(n1175), .Z(n1173) );
  XNOR U1000 ( .A(p_input[1023]), .B(n1172), .Z(n1175) );
  XOR U1001 ( .A(n1172), .B(p_input[1007]), .Z(n1174) );
  XOR U1002 ( .A(n1176), .B(n1177), .Z(n1172) );
  AND U1003 ( .A(n1178), .B(n1179), .Z(n1177) );
  XNOR U1004 ( .A(p_input[1022]), .B(n1176), .Z(n1179) );
  XOR U1005 ( .A(n1176), .B(p_input[1006]), .Z(n1178) );
  XOR U1006 ( .A(n1180), .B(n1181), .Z(n1176) );
  AND U1007 ( .A(n1182), .B(n1183), .Z(n1181) );
  XNOR U1008 ( .A(p_input[1021]), .B(n1180), .Z(n1183) );
  XOR U1009 ( .A(n1180), .B(p_input[1005]), .Z(n1182) );
  XOR U1010 ( .A(n1184), .B(n1185), .Z(n1180) );
  AND U1011 ( .A(n1186), .B(n1187), .Z(n1185) );
  XNOR U1012 ( .A(p_input[1020]), .B(n1184), .Z(n1187) );
  XOR U1013 ( .A(n1184), .B(p_input[1004]), .Z(n1186) );
  XOR U1014 ( .A(n1188), .B(n1189), .Z(n1184) );
  AND U1015 ( .A(n1190), .B(n1191), .Z(n1189) );
  XNOR U1016 ( .A(p_input[1019]), .B(n1188), .Z(n1191) );
  XOR U1017 ( .A(n1188), .B(p_input[1003]), .Z(n1190) );
  XOR U1018 ( .A(n1192), .B(n1193), .Z(n1188) );
  AND U1019 ( .A(n1194), .B(n1195), .Z(n1193) );
  XNOR U1020 ( .A(p_input[1018]), .B(n1192), .Z(n1195) );
  XOR U1021 ( .A(n1192), .B(p_input[1002]), .Z(n1194) );
  XOR U1022 ( .A(n1196), .B(n1197), .Z(n1192) );
  AND U1023 ( .A(n1198), .B(n1199), .Z(n1197) );
  XNOR U1024 ( .A(p_input[1017]), .B(n1196), .Z(n1199) );
  XOR U1025 ( .A(n1196), .B(p_input[1001]), .Z(n1198) );
  XOR U1026 ( .A(n1200), .B(n1201), .Z(n1196) );
  AND U1027 ( .A(n1202), .B(n1203), .Z(n1201) );
  XNOR U1028 ( .A(p_input[1016]), .B(n1200), .Z(n1203) );
  XOR U1029 ( .A(n1200), .B(p_input[1000]), .Z(n1202) );
  XOR U1030 ( .A(n1204), .B(n1205), .Z(n1200) );
  AND U1031 ( .A(n1206), .B(n1207), .Z(n1205) );
  XNOR U1032 ( .A(p_input[1015]), .B(n1204), .Z(n1207) );
  XOR U1033 ( .A(n1204), .B(p_input[999]), .Z(n1206) );
  XOR U1034 ( .A(n1208), .B(n1209), .Z(n1204) );
  AND U1035 ( .A(n1210), .B(n1211), .Z(n1209) );
  XNOR U1036 ( .A(p_input[1014]), .B(n1208), .Z(n1211) );
  XOR U1037 ( .A(n1208), .B(p_input[998]), .Z(n1210) );
  XOR U1038 ( .A(n1212), .B(n1213), .Z(n1208) );
  AND U1039 ( .A(n1214), .B(n1215), .Z(n1213) );
  XNOR U1040 ( .A(p_input[1013]), .B(n1212), .Z(n1215) );
  XOR U1041 ( .A(n1212), .B(p_input[997]), .Z(n1214) );
  XOR U1042 ( .A(n1216), .B(n1217), .Z(n1212) );
  AND U1043 ( .A(n1218), .B(n1219), .Z(n1217) );
  XNOR U1044 ( .A(p_input[1012]), .B(n1216), .Z(n1219) );
  XOR U1045 ( .A(n1216), .B(p_input[996]), .Z(n1218) );
  XOR U1046 ( .A(n1220), .B(n1221), .Z(n1216) );
  AND U1047 ( .A(n1222), .B(n1223), .Z(n1221) );
  XNOR U1048 ( .A(p_input[1011]), .B(n1220), .Z(n1223) );
  XOR U1049 ( .A(n1220), .B(p_input[995]), .Z(n1222) );
  XOR U1050 ( .A(n1224), .B(n1225), .Z(n1220) );
  AND U1051 ( .A(n1226), .B(n1227), .Z(n1225) );
  XNOR U1052 ( .A(p_input[1010]), .B(n1224), .Z(n1227) );
  XOR U1053 ( .A(n1224), .B(p_input[994]), .Z(n1226) );
  XNOR U1054 ( .A(n1228), .B(n1229), .Z(n1224) );
  AND U1055 ( .A(n1230), .B(n1231), .Z(n1229) );
  XOR U1056 ( .A(p_input[1009]), .B(n1228), .Z(n1231) );
  XNOR U1057 ( .A(p_input[993]), .B(n1228), .Z(n1230) );
  AND U1058 ( .A(p_input[1008]), .B(n1232), .Z(n1228) );
  IV U1059 ( .A(p_input[992]), .Z(n1232) );
  XNOR U1060 ( .A(p_input[960]), .B(n1233), .Z(n1035) );
  AND U1061 ( .A(n96), .B(n1234), .Z(n1233) );
  XOR U1062 ( .A(p_input[976]), .B(p_input[960]), .Z(n1234) );
  XOR U1063 ( .A(n1235), .B(n1236), .Z(n96) );
  AND U1064 ( .A(n1237), .B(n1238), .Z(n1236) );
  XNOR U1065 ( .A(p_input[991]), .B(n1235), .Z(n1238) );
  XOR U1066 ( .A(n1235), .B(p_input[975]), .Z(n1237) );
  XOR U1067 ( .A(n1239), .B(n1240), .Z(n1235) );
  AND U1068 ( .A(n1241), .B(n1242), .Z(n1240) );
  XNOR U1069 ( .A(p_input[990]), .B(n1239), .Z(n1242) );
  XNOR U1070 ( .A(n1239), .B(n1049), .Z(n1241) );
  IV U1071 ( .A(p_input[974]), .Z(n1049) );
  XOR U1072 ( .A(n1243), .B(n1244), .Z(n1239) );
  AND U1073 ( .A(n1245), .B(n1246), .Z(n1244) );
  XNOR U1074 ( .A(p_input[989]), .B(n1243), .Z(n1246) );
  XNOR U1075 ( .A(n1243), .B(n1058), .Z(n1245) );
  IV U1076 ( .A(p_input[973]), .Z(n1058) );
  XOR U1077 ( .A(n1247), .B(n1248), .Z(n1243) );
  AND U1078 ( .A(n1249), .B(n1250), .Z(n1248) );
  XNOR U1079 ( .A(p_input[988]), .B(n1247), .Z(n1250) );
  XNOR U1080 ( .A(n1247), .B(n1067), .Z(n1249) );
  IV U1081 ( .A(p_input[972]), .Z(n1067) );
  XOR U1082 ( .A(n1251), .B(n1252), .Z(n1247) );
  AND U1083 ( .A(n1253), .B(n1254), .Z(n1252) );
  XNOR U1084 ( .A(p_input[987]), .B(n1251), .Z(n1254) );
  XNOR U1085 ( .A(n1251), .B(n1076), .Z(n1253) );
  IV U1086 ( .A(p_input[971]), .Z(n1076) );
  XOR U1087 ( .A(n1255), .B(n1256), .Z(n1251) );
  AND U1088 ( .A(n1257), .B(n1258), .Z(n1256) );
  XNOR U1089 ( .A(p_input[986]), .B(n1255), .Z(n1258) );
  XNOR U1090 ( .A(n1255), .B(n1085), .Z(n1257) );
  IV U1091 ( .A(p_input[970]), .Z(n1085) );
  XOR U1092 ( .A(n1259), .B(n1260), .Z(n1255) );
  AND U1093 ( .A(n1261), .B(n1262), .Z(n1260) );
  XNOR U1094 ( .A(p_input[985]), .B(n1259), .Z(n1262) );
  XNOR U1095 ( .A(n1259), .B(n1094), .Z(n1261) );
  IV U1096 ( .A(p_input[969]), .Z(n1094) );
  XOR U1097 ( .A(n1263), .B(n1264), .Z(n1259) );
  AND U1098 ( .A(n1265), .B(n1266), .Z(n1264) );
  XNOR U1099 ( .A(p_input[984]), .B(n1263), .Z(n1266) );
  XNOR U1100 ( .A(n1263), .B(n1103), .Z(n1265) );
  IV U1101 ( .A(p_input[968]), .Z(n1103) );
  XOR U1102 ( .A(n1267), .B(n1268), .Z(n1263) );
  AND U1103 ( .A(n1269), .B(n1270), .Z(n1268) );
  XNOR U1104 ( .A(p_input[983]), .B(n1267), .Z(n1270) );
  XNOR U1105 ( .A(n1267), .B(n1112), .Z(n1269) );
  IV U1106 ( .A(p_input[967]), .Z(n1112) );
  XOR U1107 ( .A(n1271), .B(n1272), .Z(n1267) );
  AND U1108 ( .A(n1273), .B(n1274), .Z(n1272) );
  XNOR U1109 ( .A(p_input[982]), .B(n1271), .Z(n1274) );
  XNOR U1110 ( .A(n1271), .B(n1121), .Z(n1273) );
  IV U1111 ( .A(p_input[966]), .Z(n1121) );
  XOR U1112 ( .A(n1275), .B(n1276), .Z(n1271) );
  AND U1113 ( .A(n1277), .B(n1278), .Z(n1276) );
  XNOR U1114 ( .A(p_input[981]), .B(n1275), .Z(n1278) );
  XNOR U1115 ( .A(n1275), .B(n1130), .Z(n1277) );
  IV U1116 ( .A(p_input[965]), .Z(n1130) );
  XOR U1117 ( .A(n1279), .B(n1280), .Z(n1275) );
  AND U1118 ( .A(n1281), .B(n1282), .Z(n1280) );
  XNOR U1119 ( .A(p_input[980]), .B(n1279), .Z(n1282) );
  XNOR U1120 ( .A(n1279), .B(n1139), .Z(n1281) );
  IV U1121 ( .A(p_input[964]), .Z(n1139) );
  XOR U1122 ( .A(n1283), .B(n1284), .Z(n1279) );
  AND U1123 ( .A(n1285), .B(n1286), .Z(n1284) );
  XNOR U1124 ( .A(p_input[979]), .B(n1283), .Z(n1286) );
  XNOR U1125 ( .A(n1283), .B(n1148), .Z(n1285) );
  IV U1126 ( .A(p_input[963]), .Z(n1148) );
  XOR U1127 ( .A(n1287), .B(n1288), .Z(n1283) );
  AND U1128 ( .A(n1289), .B(n1290), .Z(n1288) );
  XNOR U1129 ( .A(p_input[978]), .B(n1287), .Z(n1290) );
  XNOR U1130 ( .A(n1287), .B(n1157), .Z(n1289) );
  IV U1131 ( .A(p_input[962]), .Z(n1157) );
  XNOR U1132 ( .A(n1291), .B(n1292), .Z(n1287) );
  AND U1133 ( .A(n1293), .B(n1294), .Z(n1292) );
  XOR U1134 ( .A(p_input[977]), .B(n1291), .Z(n1294) );
  XNOR U1135 ( .A(p_input[961]), .B(n1291), .Z(n1293) );
  AND U1136 ( .A(p_input[976]), .B(n1295), .Z(n1291) );
  IV U1137 ( .A(p_input[960]), .Z(n1295) );
  XOR U1138 ( .A(n1296), .B(n1297), .Z(n854) );
  AND U1139 ( .A(n156), .B(n1298), .Z(n1297) );
  XNOR U1140 ( .A(n1299), .B(n1296), .Z(n1298) );
  XOR U1141 ( .A(n1300), .B(n1301), .Z(n156) );
  AND U1142 ( .A(n1302), .B(n1303), .Z(n1301) );
  XNOR U1143 ( .A(n864), .B(n1300), .Z(n1303) );
  AND U1144 ( .A(p_input[959]), .B(p_input[943]), .Z(n864) );
  XOR U1145 ( .A(n1300), .B(n865), .Z(n1302) );
  AND U1146 ( .A(p_input[927]), .B(p_input[911]), .Z(n865) );
  XOR U1147 ( .A(n1304), .B(n1305), .Z(n1300) );
  AND U1148 ( .A(n1306), .B(n1307), .Z(n1305) );
  XOR U1149 ( .A(n1304), .B(n877), .Z(n1307) );
  XNOR U1150 ( .A(p_input[942]), .B(n1308), .Z(n877) );
  AND U1151 ( .A(n102), .B(n1309), .Z(n1308) );
  XOR U1152 ( .A(p_input[958]), .B(p_input[942]), .Z(n1309) );
  XNOR U1153 ( .A(n874), .B(n1304), .Z(n1306) );
  XOR U1154 ( .A(n1310), .B(n1311), .Z(n874) );
  AND U1155 ( .A(n99), .B(n1312), .Z(n1311) );
  XOR U1156 ( .A(p_input[926]), .B(p_input[910]), .Z(n1312) );
  XOR U1157 ( .A(n1313), .B(n1314), .Z(n1304) );
  AND U1158 ( .A(n1315), .B(n1316), .Z(n1314) );
  XOR U1159 ( .A(n1313), .B(n889), .Z(n1316) );
  XNOR U1160 ( .A(p_input[941]), .B(n1317), .Z(n889) );
  AND U1161 ( .A(n102), .B(n1318), .Z(n1317) );
  XOR U1162 ( .A(p_input[957]), .B(p_input[941]), .Z(n1318) );
  XNOR U1163 ( .A(n886), .B(n1313), .Z(n1315) );
  XOR U1164 ( .A(n1319), .B(n1320), .Z(n886) );
  AND U1165 ( .A(n99), .B(n1321), .Z(n1320) );
  XOR U1166 ( .A(p_input[925]), .B(p_input[909]), .Z(n1321) );
  XOR U1167 ( .A(n1322), .B(n1323), .Z(n1313) );
  AND U1168 ( .A(n1324), .B(n1325), .Z(n1323) );
  XOR U1169 ( .A(n1322), .B(n901), .Z(n1325) );
  XNOR U1170 ( .A(p_input[940]), .B(n1326), .Z(n901) );
  AND U1171 ( .A(n102), .B(n1327), .Z(n1326) );
  XOR U1172 ( .A(p_input[956]), .B(p_input[940]), .Z(n1327) );
  XNOR U1173 ( .A(n898), .B(n1322), .Z(n1324) );
  XOR U1174 ( .A(n1328), .B(n1329), .Z(n898) );
  AND U1175 ( .A(n99), .B(n1330), .Z(n1329) );
  XOR U1176 ( .A(p_input[924]), .B(p_input[908]), .Z(n1330) );
  XOR U1177 ( .A(n1331), .B(n1332), .Z(n1322) );
  AND U1178 ( .A(n1333), .B(n1334), .Z(n1332) );
  XOR U1179 ( .A(n1331), .B(n913), .Z(n1334) );
  XNOR U1180 ( .A(p_input[939]), .B(n1335), .Z(n913) );
  AND U1181 ( .A(n102), .B(n1336), .Z(n1335) );
  XOR U1182 ( .A(p_input[955]), .B(p_input[939]), .Z(n1336) );
  XNOR U1183 ( .A(n910), .B(n1331), .Z(n1333) );
  XOR U1184 ( .A(n1337), .B(n1338), .Z(n910) );
  AND U1185 ( .A(n99), .B(n1339), .Z(n1338) );
  XOR U1186 ( .A(p_input[923]), .B(p_input[907]), .Z(n1339) );
  XOR U1187 ( .A(n1340), .B(n1341), .Z(n1331) );
  AND U1188 ( .A(n1342), .B(n1343), .Z(n1341) );
  XOR U1189 ( .A(n1340), .B(n925), .Z(n1343) );
  XNOR U1190 ( .A(p_input[938]), .B(n1344), .Z(n925) );
  AND U1191 ( .A(n102), .B(n1345), .Z(n1344) );
  XOR U1192 ( .A(p_input[954]), .B(p_input[938]), .Z(n1345) );
  XNOR U1193 ( .A(n922), .B(n1340), .Z(n1342) );
  XOR U1194 ( .A(n1346), .B(n1347), .Z(n922) );
  AND U1195 ( .A(n99), .B(n1348), .Z(n1347) );
  XOR U1196 ( .A(p_input[922]), .B(p_input[906]), .Z(n1348) );
  XOR U1197 ( .A(n1349), .B(n1350), .Z(n1340) );
  AND U1198 ( .A(n1351), .B(n1352), .Z(n1350) );
  XOR U1199 ( .A(n1349), .B(n937), .Z(n1352) );
  XNOR U1200 ( .A(p_input[937]), .B(n1353), .Z(n937) );
  AND U1201 ( .A(n102), .B(n1354), .Z(n1353) );
  XOR U1202 ( .A(p_input[953]), .B(p_input[937]), .Z(n1354) );
  XNOR U1203 ( .A(n934), .B(n1349), .Z(n1351) );
  XOR U1204 ( .A(n1355), .B(n1356), .Z(n934) );
  AND U1205 ( .A(n99), .B(n1357), .Z(n1356) );
  XOR U1206 ( .A(p_input[921]), .B(p_input[905]), .Z(n1357) );
  XOR U1207 ( .A(n1358), .B(n1359), .Z(n1349) );
  AND U1208 ( .A(n1360), .B(n1361), .Z(n1359) );
  XOR U1209 ( .A(n1358), .B(n949), .Z(n1361) );
  XNOR U1210 ( .A(p_input[936]), .B(n1362), .Z(n949) );
  AND U1211 ( .A(n102), .B(n1363), .Z(n1362) );
  XOR U1212 ( .A(p_input[952]), .B(p_input[936]), .Z(n1363) );
  XNOR U1213 ( .A(n946), .B(n1358), .Z(n1360) );
  XOR U1214 ( .A(n1364), .B(n1365), .Z(n946) );
  AND U1215 ( .A(n99), .B(n1366), .Z(n1365) );
  XOR U1216 ( .A(p_input[920]), .B(p_input[904]), .Z(n1366) );
  XOR U1217 ( .A(n1367), .B(n1368), .Z(n1358) );
  AND U1218 ( .A(n1369), .B(n1370), .Z(n1368) );
  XOR U1219 ( .A(n1367), .B(n961), .Z(n1370) );
  XNOR U1220 ( .A(p_input[935]), .B(n1371), .Z(n961) );
  AND U1221 ( .A(n102), .B(n1372), .Z(n1371) );
  XOR U1222 ( .A(p_input[951]), .B(p_input[935]), .Z(n1372) );
  XNOR U1223 ( .A(n958), .B(n1367), .Z(n1369) );
  XOR U1224 ( .A(n1373), .B(n1374), .Z(n958) );
  AND U1225 ( .A(n99), .B(n1375), .Z(n1374) );
  XOR U1226 ( .A(p_input[919]), .B(p_input[903]), .Z(n1375) );
  XOR U1227 ( .A(n1376), .B(n1377), .Z(n1367) );
  AND U1228 ( .A(n1378), .B(n1379), .Z(n1377) );
  XOR U1229 ( .A(n1376), .B(n973), .Z(n1379) );
  XNOR U1230 ( .A(p_input[934]), .B(n1380), .Z(n973) );
  AND U1231 ( .A(n102), .B(n1381), .Z(n1380) );
  XOR U1232 ( .A(p_input[950]), .B(p_input[934]), .Z(n1381) );
  XNOR U1233 ( .A(n970), .B(n1376), .Z(n1378) );
  XOR U1234 ( .A(n1382), .B(n1383), .Z(n970) );
  AND U1235 ( .A(n99), .B(n1384), .Z(n1383) );
  XOR U1236 ( .A(p_input[918]), .B(p_input[902]), .Z(n1384) );
  XOR U1237 ( .A(n1385), .B(n1386), .Z(n1376) );
  AND U1238 ( .A(n1387), .B(n1388), .Z(n1386) );
  XOR U1239 ( .A(n1385), .B(n985), .Z(n1388) );
  XNOR U1240 ( .A(p_input[933]), .B(n1389), .Z(n985) );
  AND U1241 ( .A(n102), .B(n1390), .Z(n1389) );
  XOR U1242 ( .A(p_input[949]), .B(p_input[933]), .Z(n1390) );
  XNOR U1243 ( .A(n982), .B(n1385), .Z(n1387) );
  XOR U1244 ( .A(n1391), .B(n1392), .Z(n982) );
  AND U1245 ( .A(n99), .B(n1393), .Z(n1392) );
  XOR U1246 ( .A(p_input[917]), .B(p_input[901]), .Z(n1393) );
  XOR U1247 ( .A(n1394), .B(n1395), .Z(n1385) );
  AND U1248 ( .A(n1396), .B(n1397), .Z(n1395) );
  XOR U1249 ( .A(n1394), .B(n997), .Z(n1397) );
  XNOR U1250 ( .A(p_input[932]), .B(n1398), .Z(n997) );
  AND U1251 ( .A(n102), .B(n1399), .Z(n1398) );
  XOR U1252 ( .A(p_input[948]), .B(p_input[932]), .Z(n1399) );
  XNOR U1253 ( .A(n994), .B(n1394), .Z(n1396) );
  XOR U1254 ( .A(n1400), .B(n1401), .Z(n994) );
  AND U1255 ( .A(n99), .B(n1402), .Z(n1401) );
  XOR U1256 ( .A(p_input[916]), .B(p_input[900]), .Z(n1402) );
  XOR U1257 ( .A(n1403), .B(n1404), .Z(n1394) );
  AND U1258 ( .A(n1405), .B(n1406), .Z(n1404) );
  XOR U1259 ( .A(n1009), .B(n1403), .Z(n1406) );
  XNOR U1260 ( .A(p_input[931]), .B(n1407), .Z(n1009) );
  AND U1261 ( .A(n102), .B(n1408), .Z(n1407) );
  XOR U1262 ( .A(p_input[947]), .B(p_input[931]), .Z(n1408) );
  XNOR U1263 ( .A(n1403), .B(n1006), .Z(n1405) );
  XOR U1264 ( .A(n1409), .B(n1410), .Z(n1006) );
  AND U1265 ( .A(n99), .B(n1411), .Z(n1410) );
  XOR U1266 ( .A(p_input[915]), .B(p_input[899]), .Z(n1411) );
  XOR U1267 ( .A(n1412), .B(n1413), .Z(n1403) );
  AND U1268 ( .A(n1414), .B(n1415), .Z(n1413) );
  XOR U1269 ( .A(n1412), .B(n1021), .Z(n1415) );
  XNOR U1270 ( .A(p_input[930]), .B(n1416), .Z(n1021) );
  AND U1271 ( .A(n102), .B(n1417), .Z(n1416) );
  XOR U1272 ( .A(p_input[946]), .B(p_input[930]), .Z(n1417) );
  XNOR U1273 ( .A(n1018), .B(n1412), .Z(n1414) );
  XOR U1274 ( .A(n1418), .B(n1419), .Z(n1018) );
  AND U1275 ( .A(n99), .B(n1420), .Z(n1419) );
  XOR U1276 ( .A(p_input[914]), .B(p_input[898]), .Z(n1420) );
  XOR U1277 ( .A(n1421), .B(n1422), .Z(n1412) );
  AND U1278 ( .A(n1423), .B(n1424), .Z(n1422) );
  XNOR U1279 ( .A(n1425), .B(n1034), .Z(n1424) );
  XNOR U1280 ( .A(p_input[929]), .B(n1426), .Z(n1034) );
  AND U1281 ( .A(n102), .B(n1427), .Z(n1426) );
  XNOR U1282 ( .A(p_input[945]), .B(n1428), .Z(n1427) );
  IV U1283 ( .A(p_input[929]), .Z(n1428) );
  XNOR U1284 ( .A(n1031), .B(n1421), .Z(n1423) );
  XNOR U1285 ( .A(p_input[897]), .B(n1429), .Z(n1031) );
  AND U1286 ( .A(n99), .B(n1430), .Z(n1429) );
  XOR U1287 ( .A(p_input[913]), .B(p_input[897]), .Z(n1430) );
  IV U1288 ( .A(n1425), .Z(n1421) );
  AND U1289 ( .A(n1296), .B(n1299), .Z(n1425) );
  XOR U1290 ( .A(p_input[928]), .B(n1431), .Z(n1299) );
  AND U1291 ( .A(n102), .B(n1432), .Z(n1431) );
  XOR U1292 ( .A(p_input[944]), .B(p_input[928]), .Z(n1432) );
  XOR U1293 ( .A(n1433), .B(n1434), .Z(n102) );
  AND U1294 ( .A(n1435), .B(n1436), .Z(n1434) );
  XNOR U1295 ( .A(p_input[959]), .B(n1433), .Z(n1436) );
  XOR U1296 ( .A(n1433), .B(p_input[943]), .Z(n1435) );
  XOR U1297 ( .A(n1437), .B(n1438), .Z(n1433) );
  AND U1298 ( .A(n1439), .B(n1440), .Z(n1438) );
  XNOR U1299 ( .A(p_input[958]), .B(n1437), .Z(n1440) );
  XOR U1300 ( .A(n1437), .B(p_input[942]), .Z(n1439) );
  XOR U1301 ( .A(n1441), .B(n1442), .Z(n1437) );
  AND U1302 ( .A(n1443), .B(n1444), .Z(n1442) );
  XNOR U1303 ( .A(p_input[957]), .B(n1441), .Z(n1444) );
  XOR U1304 ( .A(n1441), .B(p_input[941]), .Z(n1443) );
  XOR U1305 ( .A(n1445), .B(n1446), .Z(n1441) );
  AND U1306 ( .A(n1447), .B(n1448), .Z(n1446) );
  XNOR U1307 ( .A(p_input[956]), .B(n1445), .Z(n1448) );
  XOR U1308 ( .A(n1445), .B(p_input[940]), .Z(n1447) );
  XOR U1309 ( .A(n1449), .B(n1450), .Z(n1445) );
  AND U1310 ( .A(n1451), .B(n1452), .Z(n1450) );
  XNOR U1311 ( .A(p_input[955]), .B(n1449), .Z(n1452) );
  XOR U1312 ( .A(n1449), .B(p_input[939]), .Z(n1451) );
  XOR U1313 ( .A(n1453), .B(n1454), .Z(n1449) );
  AND U1314 ( .A(n1455), .B(n1456), .Z(n1454) );
  XNOR U1315 ( .A(p_input[954]), .B(n1453), .Z(n1456) );
  XOR U1316 ( .A(n1453), .B(p_input[938]), .Z(n1455) );
  XOR U1317 ( .A(n1457), .B(n1458), .Z(n1453) );
  AND U1318 ( .A(n1459), .B(n1460), .Z(n1458) );
  XNOR U1319 ( .A(p_input[953]), .B(n1457), .Z(n1460) );
  XOR U1320 ( .A(n1457), .B(p_input[937]), .Z(n1459) );
  XOR U1321 ( .A(n1461), .B(n1462), .Z(n1457) );
  AND U1322 ( .A(n1463), .B(n1464), .Z(n1462) );
  XNOR U1323 ( .A(p_input[952]), .B(n1461), .Z(n1464) );
  XOR U1324 ( .A(n1461), .B(p_input[936]), .Z(n1463) );
  XOR U1325 ( .A(n1465), .B(n1466), .Z(n1461) );
  AND U1326 ( .A(n1467), .B(n1468), .Z(n1466) );
  XNOR U1327 ( .A(p_input[951]), .B(n1465), .Z(n1468) );
  XOR U1328 ( .A(n1465), .B(p_input[935]), .Z(n1467) );
  XOR U1329 ( .A(n1469), .B(n1470), .Z(n1465) );
  AND U1330 ( .A(n1471), .B(n1472), .Z(n1470) );
  XNOR U1331 ( .A(p_input[950]), .B(n1469), .Z(n1472) );
  XOR U1332 ( .A(n1469), .B(p_input[934]), .Z(n1471) );
  XOR U1333 ( .A(n1473), .B(n1474), .Z(n1469) );
  AND U1334 ( .A(n1475), .B(n1476), .Z(n1474) );
  XNOR U1335 ( .A(p_input[949]), .B(n1473), .Z(n1476) );
  XOR U1336 ( .A(n1473), .B(p_input[933]), .Z(n1475) );
  XOR U1337 ( .A(n1477), .B(n1478), .Z(n1473) );
  AND U1338 ( .A(n1479), .B(n1480), .Z(n1478) );
  XNOR U1339 ( .A(p_input[948]), .B(n1477), .Z(n1480) );
  XOR U1340 ( .A(n1477), .B(p_input[932]), .Z(n1479) );
  XOR U1341 ( .A(n1481), .B(n1482), .Z(n1477) );
  AND U1342 ( .A(n1483), .B(n1484), .Z(n1482) );
  XNOR U1343 ( .A(p_input[947]), .B(n1481), .Z(n1484) );
  XOR U1344 ( .A(n1481), .B(p_input[931]), .Z(n1483) );
  XOR U1345 ( .A(n1485), .B(n1486), .Z(n1481) );
  AND U1346 ( .A(n1487), .B(n1488), .Z(n1486) );
  XNOR U1347 ( .A(p_input[946]), .B(n1485), .Z(n1488) );
  XOR U1348 ( .A(n1485), .B(p_input[930]), .Z(n1487) );
  XNOR U1349 ( .A(n1489), .B(n1490), .Z(n1485) );
  AND U1350 ( .A(n1491), .B(n1492), .Z(n1490) );
  XOR U1351 ( .A(p_input[945]), .B(n1489), .Z(n1492) );
  XNOR U1352 ( .A(p_input[929]), .B(n1489), .Z(n1491) );
  AND U1353 ( .A(p_input[944]), .B(n1493), .Z(n1489) );
  IV U1354 ( .A(p_input[928]), .Z(n1493) );
  XNOR U1355 ( .A(p_input[896]), .B(n1494), .Z(n1296) );
  AND U1356 ( .A(n99), .B(n1495), .Z(n1494) );
  XOR U1357 ( .A(p_input[912]), .B(p_input[896]), .Z(n1495) );
  XOR U1358 ( .A(n1496), .B(n1497), .Z(n99) );
  AND U1359 ( .A(n1498), .B(n1499), .Z(n1497) );
  XNOR U1360 ( .A(p_input[927]), .B(n1496), .Z(n1499) );
  XOR U1361 ( .A(n1496), .B(p_input[911]), .Z(n1498) );
  XOR U1362 ( .A(n1500), .B(n1501), .Z(n1496) );
  AND U1363 ( .A(n1502), .B(n1503), .Z(n1501) );
  XNOR U1364 ( .A(p_input[926]), .B(n1500), .Z(n1503) );
  XNOR U1365 ( .A(n1500), .B(n1310), .Z(n1502) );
  IV U1366 ( .A(p_input[910]), .Z(n1310) );
  XOR U1367 ( .A(n1504), .B(n1505), .Z(n1500) );
  AND U1368 ( .A(n1506), .B(n1507), .Z(n1505) );
  XNOR U1369 ( .A(p_input[925]), .B(n1504), .Z(n1507) );
  XNOR U1370 ( .A(n1504), .B(n1319), .Z(n1506) );
  IV U1371 ( .A(p_input[909]), .Z(n1319) );
  XOR U1372 ( .A(n1508), .B(n1509), .Z(n1504) );
  AND U1373 ( .A(n1510), .B(n1511), .Z(n1509) );
  XNOR U1374 ( .A(p_input[924]), .B(n1508), .Z(n1511) );
  XNOR U1375 ( .A(n1508), .B(n1328), .Z(n1510) );
  IV U1376 ( .A(p_input[908]), .Z(n1328) );
  XOR U1377 ( .A(n1512), .B(n1513), .Z(n1508) );
  AND U1378 ( .A(n1514), .B(n1515), .Z(n1513) );
  XNOR U1379 ( .A(p_input[923]), .B(n1512), .Z(n1515) );
  XNOR U1380 ( .A(n1512), .B(n1337), .Z(n1514) );
  IV U1381 ( .A(p_input[907]), .Z(n1337) );
  XOR U1382 ( .A(n1516), .B(n1517), .Z(n1512) );
  AND U1383 ( .A(n1518), .B(n1519), .Z(n1517) );
  XNOR U1384 ( .A(p_input[922]), .B(n1516), .Z(n1519) );
  XNOR U1385 ( .A(n1516), .B(n1346), .Z(n1518) );
  IV U1386 ( .A(p_input[906]), .Z(n1346) );
  XOR U1387 ( .A(n1520), .B(n1521), .Z(n1516) );
  AND U1388 ( .A(n1522), .B(n1523), .Z(n1521) );
  XNOR U1389 ( .A(p_input[921]), .B(n1520), .Z(n1523) );
  XNOR U1390 ( .A(n1520), .B(n1355), .Z(n1522) );
  IV U1391 ( .A(p_input[905]), .Z(n1355) );
  XOR U1392 ( .A(n1524), .B(n1525), .Z(n1520) );
  AND U1393 ( .A(n1526), .B(n1527), .Z(n1525) );
  XNOR U1394 ( .A(p_input[920]), .B(n1524), .Z(n1527) );
  XNOR U1395 ( .A(n1524), .B(n1364), .Z(n1526) );
  IV U1396 ( .A(p_input[904]), .Z(n1364) );
  XOR U1397 ( .A(n1528), .B(n1529), .Z(n1524) );
  AND U1398 ( .A(n1530), .B(n1531), .Z(n1529) );
  XNOR U1399 ( .A(p_input[919]), .B(n1528), .Z(n1531) );
  XNOR U1400 ( .A(n1528), .B(n1373), .Z(n1530) );
  IV U1401 ( .A(p_input[903]), .Z(n1373) );
  XOR U1402 ( .A(n1532), .B(n1533), .Z(n1528) );
  AND U1403 ( .A(n1534), .B(n1535), .Z(n1533) );
  XNOR U1404 ( .A(p_input[918]), .B(n1532), .Z(n1535) );
  XNOR U1405 ( .A(n1532), .B(n1382), .Z(n1534) );
  IV U1406 ( .A(p_input[902]), .Z(n1382) );
  XOR U1407 ( .A(n1536), .B(n1537), .Z(n1532) );
  AND U1408 ( .A(n1538), .B(n1539), .Z(n1537) );
  XNOR U1409 ( .A(p_input[917]), .B(n1536), .Z(n1539) );
  XNOR U1410 ( .A(n1536), .B(n1391), .Z(n1538) );
  IV U1411 ( .A(p_input[901]), .Z(n1391) );
  XOR U1412 ( .A(n1540), .B(n1541), .Z(n1536) );
  AND U1413 ( .A(n1542), .B(n1543), .Z(n1541) );
  XNOR U1414 ( .A(p_input[916]), .B(n1540), .Z(n1543) );
  XNOR U1415 ( .A(n1540), .B(n1400), .Z(n1542) );
  IV U1416 ( .A(p_input[900]), .Z(n1400) );
  XOR U1417 ( .A(n1544), .B(n1545), .Z(n1540) );
  AND U1418 ( .A(n1546), .B(n1547), .Z(n1545) );
  XNOR U1419 ( .A(p_input[915]), .B(n1544), .Z(n1547) );
  XNOR U1420 ( .A(n1544), .B(n1409), .Z(n1546) );
  IV U1421 ( .A(p_input[899]), .Z(n1409) );
  XOR U1422 ( .A(n1548), .B(n1549), .Z(n1544) );
  AND U1423 ( .A(n1550), .B(n1551), .Z(n1549) );
  XNOR U1424 ( .A(p_input[914]), .B(n1548), .Z(n1551) );
  XNOR U1425 ( .A(n1548), .B(n1418), .Z(n1550) );
  IV U1426 ( .A(p_input[898]), .Z(n1418) );
  XNOR U1427 ( .A(n1552), .B(n1553), .Z(n1548) );
  AND U1428 ( .A(n1554), .B(n1555), .Z(n1553) );
  XOR U1429 ( .A(p_input[913]), .B(n1552), .Z(n1555) );
  XNOR U1430 ( .A(p_input[897]), .B(n1552), .Z(n1554) );
  AND U1431 ( .A(p_input[912]), .B(n1556), .Z(n1552) );
  IV U1432 ( .A(p_input[896]), .Z(n1556) );
  XOR U1433 ( .A(n1557), .B(n1558), .Z(n672) );
  AND U1434 ( .A(n244), .B(n1559), .Z(n1558) );
  XNOR U1435 ( .A(n1560), .B(n1557), .Z(n1559) );
  XOR U1436 ( .A(n1561), .B(n1562), .Z(n244) );
  AND U1437 ( .A(n1563), .B(n1564), .Z(n1562) );
  XNOR U1438 ( .A(n684), .B(n1561), .Z(n1564) );
  AND U1439 ( .A(n1565), .B(n1566), .Z(n684) );
  XOR U1440 ( .A(n1561), .B(n683), .Z(n1563) );
  AND U1441 ( .A(n1567), .B(n1568), .Z(n683) );
  XOR U1442 ( .A(n1569), .B(n1570), .Z(n1561) );
  AND U1443 ( .A(n1571), .B(n1572), .Z(n1570) );
  XOR U1444 ( .A(n1569), .B(n696), .Z(n1572) );
  XOR U1445 ( .A(n1573), .B(n1574), .Z(n696) );
  AND U1446 ( .A(n162), .B(n1575), .Z(n1574) );
  XOR U1447 ( .A(n1576), .B(n1573), .Z(n1575) );
  XNOR U1448 ( .A(n693), .B(n1569), .Z(n1571) );
  XOR U1449 ( .A(n1577), .B(n1578), .Z(n693) );
  AND U1450 ( .A(n159), .B(n1579), .Z(n1578) );
  XOR U1451 ( .A(n1580), .B(n1577), .Z(n1579) );
  XOR U1452 ( .A(n1581), .B(n1582), .Z(n1569) );
  AND U1453 ( .A(n1583), .B(n1584), .Z(n1582) );
  XOR U1454 ( .A(n1581), .B(n708), .Z(n1584) );
  XOR U1455 ( .A(n1585), .B(n1586), .Z(n708) );
  AND U1456 ( .A(n162), .B(n1587), .Z(n1586) );
  XOR U1457 ( .A(n1588), .B(n1585), .Z(n1587) );
  XNOR U1458 ( .A(n705), .B(n1581), .Z(n1583) );
  XOR U1459 ( .A(n1589), .B(n1590), .Z(n705) );
  AND U1460 ( .A(n159), .B(n1591), .Z(n1590) );
  XOR U1461 ( .A(n1592), .B(n1589), .Z(n1591) );
  XOR U1462 ( .A(n1593), .B(n1594), .Z(n1581) );
  AND U1463 ( .A(n1595), .B(n1596), .Z(n1594) );
  XOR U1464 ( .A(n1593), .B(n720), .Z(n1596) );
  XOR U1465 ( .A(n1597), .B(n1598), .Z(n720) );
  AND U1466 ( .A(n162), .B(n1599), .Z(n1598) );
  XOR U1467 ( .A(n1600), .B(n1597), .Z(n1599) );
  XNOR U1468 ( .A(n717), .B(n1593), .Z(n1595) );
  XOR U1469 ( .A(n1601), .B(n1602), .Z(n717) );
  AND U1470 ( .A(n159), .B(n1603), .Z(n1602) );
  XOR U1471 ( .A(n1604), .B(n1601), .Z(n1603) );
  XOR U1472 ( .A(n1605), .B(n1606), .Z(n1593) );
  AND U1473 ( .A(n1607), .B(n1608), .Z(n1606) );
  XOR U1474 ( .A(n1605), .B(n732), .Z(n1608) );
  XOR U1475 ( .A(n1609), .B(n1610), .Z(n732) );
  AND U1476 ( .A(n162), .B(n1611), .Z(n1610) );
  XOR U1477 ( .A(n1612), .B(n1609), .Z(n1611) );
  XNOR U1478 ( .A(n729), .B(n1605), .Z(n1607) );
  XOR U1479 ( .A(n1613), .B(n1614), .Z(n729) );
  AND U1480 ( .A(n159), .B(n1615), .Z(n1614) );
  XOR U1481 ( .A(n1616), .B(n1613), .Z(n1615) );
  XOR U1482 ( .A(n1617), .B(n1618), .Z(n1605) );
  AND U1483 ( .A(n1619), .B(n1620), .Z(n1618) );
  XOR U1484 ( .A(n1617), .B(n744), .Z(n1620) );
  XOR U1485 ( .A(n1621), .B(n1622), .Z(n744) );
  AND U1486 ( .A(n162), .B(n1623), .Z(n1622) );
  XOR U1487 ( .A(n1624), .B(n1621), .Z(n1623) );
  XNOR U1488 ( .A(n741), .B(n1617), .Z(n1619) );
  XOR U1489 ( .A(n1625), .B(n1626), .Z(n741) );
  AND U1490 ( .A(n159), .B(n1627), .Z(n1626) );
  XOR U1491 ( .A(n1628), .B(n1625), .Z(n1627) );
  XOR U1492 ( .A(n1629), .B(n1630), .Z(n1617) );
  AND U1493 ( .A(n1631), .B(n1632), .Z(n1630) );
  XOR U1494 ( .A(n1629), .B(n756), .Z(n1632) );
  XOR U1495 ( .A(n1633), .B(n1634), .Z(n756) );
  AND U1496 ( .A(n162), .B(n1635), .Z(n1634) );
  XOR U1497 ( .A(n1636), .B(n1633), .Z(n1635) );
  XNOR U1498 ( .A(n753), .B(n1629), .Z(n1631) );
  XOR U1499 ( .A(n1637), .B(n1638), .Z(n753) );
  AND U1500 ( .A(n159), .B(n1639), .Z(n1638) );
  XOR U1501 ( .A(n1640), .B(n1637), .Z(n1639) );
  XOR U1502 ( .A(n1641), .B(n1642), .Z(n1629) );
  AND U1503 ( .A(n1643), .B(n1644), .Z(n1642) );
  XOR U1504 ( .A(n1641), .B(n768), .Z(n1644) );
  XOR U1505 ( .A(n1645), .B(n1646), .Z(n768) );
  AND U1506 ( .A(n162), .B(n1647), .Z(n1646) );
  XOR U1507 ( .A(n1648), .B(n1645), .Z(n1647) );
  XNOR U1508 ( .A(n765), .B(n1641), .Z(n1643) );
  XOR U1509 ( .A(n1649), .B(n1650), .Z(n765) );
  AND U1510 ( .A(n159), .B(n1651), .Z(n1650) );
  XOR U1511 ( .A(n1652), .B(n1649), .Z(n1651) );
  XOR U1512 ( .A(n1653), .B(n1654), .Z(n1641) );
  AND U1513 ( .A(n1655), .B(n1656), .Z(n1654) );
  XOR U1514 ( .A(n1653), .B(n780), .Z(n1656) );
  XOR U1515 ( .A(n1657), .B(n1658), .Z(n780) );
  AND U1516 ( .A(n162), .B(n1659), .Z(n1658) );
  XOR U1517 ( .A(n1660), .B(n1657), .Z(n1659) );
  XNOR U1518 ( .A(n777), .B(n1653), .Z(n1655) );
  XOR U1519 ( .A(n1661), .B(n1662), .Z(n777) );
  AND U1520 ( .A(n159), .B(n1663), .Z(n1662) );
  XOR U1521 ( .A(n1664), .B(n1661), .Z(n1663) );
  XOR U1522 ( .A(n1665), .B(n1666), .Z(n1653) );
  AND U1523 ( .A(n1667), .B(n1668), .Z(n1666) );
  XOR U1524 ( .A(n1665), .B(n792), .Z(n1668) );
  XOR U1525 ( .A(n1669), .B(n1670), .Z(n792) );
  AND U1526 ( .A(n162), .B(n1671), .Z(n1670) );
  XOR U1527 ( .A(n1672), .B(n1669), .Z(n1671) );
  XNOR U1528 ( .A(n789), .B(n1665), .Z(n1667) );
  XOR U1529 ( .A(n1673), .B(n1674), .Z(n789) );
  AND U1530 ( .A(n159), .B(n1675), .Z(n1674) );
  XOR U1531 ( .A(n1676), .B(n1673), .Z(n1675) );
  XOR U1532 ( .A(n1677), .B(n1678), .Z(n1665) );
  AND U1533 ( .A(n1679), .B(n1680), .Z(n1678) );
  XOR U1534 ( .A(n1677), .B(n804), .Z(n1680) );
  XOR U1535 ( .A(n1681), .B(n1682), .Z(n804) );
  AND U1536 ( .A(n162), .B(n1683), .Z(n1682) );
  XOR U1537 ( .A(n1684), .B(n1681), .Z(n1683) );
  XNOR U1538 ( .A(n801), .B(n1677), .Z(n1679) );
  XOR U1539 ( .A(n1685), .B(n1686), .Z(n801) );
  AND U1540 ( .A(n159), .B(n1687), .Z(n1686) );
  XOR U1541 ( .A(n1688), .B(n1685), .Z(n1687) );
  XOR U1542 ( .A(n1689), .B(n1690), .Z(n1677) );
  AND U1543 ( .A(n1691), .B(n1692), .Z(n1690) );
  XOR U1544 ( .A(n1689), .B(n816), .Z(n1692) );
  XOR U1545 ( .A(n1693), .B(n1694), .Z(n816) );
  AND U1546 ( .A(n162), .B(n1695), .Z(n1694) );
  XOR U1547 ( .A(n1696), .B(n1693), .Z(n1695) );
  XNOR U1548 ( .A(n813), .B(n1689), .Z(n1691) );
  XOR U1549 ( .A(n1697), .B(n1698), .Z(n813) );
  AND U1550 ( .A(n159), .B(n1699), .Z(n1698) );
  XOR U1551 ( .A(n1700), .B(n1697), .Z(n1699) );
  XOR U1552 ( .A(n1701), .B(n1702), .Z(n1689) );
  AND U1553 ( .A(n1703), .B(n1704), .Z(n1702) );
  XOR U1554 ( .A(n828), .B(n1701), .Z(n1704) );
  XOR U1555 ( .A(n1705), .B(n1706), .Z(n828) );
  AND U1556 ( .A(n162), .B(n1707), .Z(n1706) );
  XOR U1557 ( .A(n1705), .B(n1708), .Z(n1707) );
  XNOR U1558 ( .A(n1701), .B(n825), .Z(n1703) );
  XOR U1559 ( .A(n1709), .B(n1710), .Z(n825) );
  AND U1560 ( .A(n159), .B(n1711), .Z(n1710) );
  XOR U1561 ( .A(n1709), .B(n1712), .Z(n1711) );
  XOR U1562 ( .A(n1713), .B(n1714), .Z(n1701) );
  AND U1563 ( .A(n1715), .B(n1716), .Z(n1714) );
  XOR U1564 ( .A(n1713), .B(n840), .Z(n1716) );
  XOR U1565 ( .A(n1717), .B(n1718), .Z(n840) );
  AND U1566 ( .A(n162), .B(n1719), .Z(n1718) );
  XOR U1567 ( .A(n1720), .B(n1717), .Z(n1719) );
  XNOR U1568 ( .A(n837), .B(n1713), .Z(n1715) );
  XOR U1569 ( .A(n1721), .B(n1722), .Z(n837) );
  AND U1570 ( .A(n159), .B(n1723), .Z(n1722) );
  XOR U1571 ( .A(n1724), .B(n1721), .Z(n1723) );
  XOR U1572 ( .A(n1725), .B(n1726), .Z(n1713) );
  AND U1573 ( .A(n1727), .B(n1728), .Z(n1726) );
  XNOR U1574 ( .A(n1729), .B(n853), .Z(n1728) );
  XOR U1575 ( .A(n1730), .B(n1731), .Z(n853) );
  AND U1576 ( .A(n162), .B(n1732), .Z(n1731) );
  XOR U1577 ( .A(n1733), .B(n1730), .Z(n1732) );
  XNOR U1578 ( .A(n850), .B(n1725), .Z(n1727) );
  XOR U1579 ( .A(n1734), .B(n1735), .Z(n850) );
  AND U1580 ( .A(n159), .B(n1736), .Z(n1735) );
  XOR U1581 ( .A(n1737), .B(n1734), .Z(n1736) );
  IV U1582 ( .A(n1729), .Z(n1725) );
  AND U1583 ( .A(n1557), .B(n1560), .Z(n1729) );
  XNOR U1584 ( .A(n1738), .B(n1739), .Z(n1560) );
  AND U1585 ( .A(n162), .B(n1740), .Z(n1739) );
  XNOR U1586 ( .A(n1741), .B(n1738), .Z(n1740) );
  XOR U1587 ( .A(n1742), .B(n1743), .Z(n162) );
  AND U1588 ( .A(n1744), .B(n1745), .Z(n1743) );
  XNOR U1589 ( .A(n1565), .B(n1742), .Z(n1745) );
  AND U1590 ( .A(p_input[895]), .B(p_input[879]), .Z(n1565) );
  XOR U1591 ( .A(n1742), .B(n1566), .Z(n1744) );
  AND U1592 ( .A(p_input[863]), .B(p_input[847]), .Z(n1566) );
  XOR U1593 ( .A(n1746), .B(n1747), .Z(n1742) );
  AND U1594 ( .A(n1748), .B(n1749), .Z(n1747) );
  XOR U1595 ( .A(n1746), .B(n1576), .Z(n1749) );
  XNOR U1596 ( .A(p_input[878]), .B(n1750), .Z(n1576) );
  AND U1597 ( .A(n110), .B(n1751), .Z(n1750) );
  XOR U1598 ( .A(p_input[894]), .B(p_input[878]), .Z(n1751) );
  XNOR U1599 ( .A(n1573), .B(n1746), .Z(n1748) );
  XOR U1600 ( .A(n1752), .B(n1753), .Z(n1573) );
  AND U1601 ( .A(n108), .B(n1754), .Z(n1753) );
  XOR U1602 ( .A(p_input[862]), .B(p_input[846]), .Z(n1754) );
  XOR U1603 ( .A(n1755), .B(n1756), .Z(n1746) );
  AND U1604 ( .A(n1757), .B(n1758), .Z(n1756) );
  XOR U1605 ( .A(n1755), .B(n1588), .Z(n1758) );
  XNOR U1606 ( .A(p_input[877]), .B(n1759), .Z(n1588) );
  AND U1607 ( .A(n110), .B(n1760), .Z(n1759) );
  XOR U1608 ( .A(p_input[893]), .B(p_input[877]), .Z(n1760) );
  XNOR U1609 ( .A(n1585), .B(n1755), .Z(n1757) );
  XOR U1610 ( .A(n1761), .B(n1762), .Z(n1585) );
  AND U1611 ( .A(n108), .B(n1763), .Z(n1762) );
  XOR U1612 ( .A(p_input[861]), .B(p_input[845]), .Z(n1763) );
  XOR U1613 ( .A(n1764), .B(n1765), .Z(n1755) );
  AND U1614 ( .A(n1766), .B(n1767), .Z(n1765) );
  XOR U1615 ( .A(n1764), .B(n1600), .Z(n1767) );
  XNOR U1616 ( .A(p_input[876]), .B(n1768), .Z(n1600) );
  AND U1617 ( .A(n110), .B(n1769), .Z(n1768) );
  XOR U1618 ( .A(p_input[892]), .B(p_input[876]), .Z(n1769) );
  XNOR U1619 ( .A(n1597), .B(n1764), .Z(n1766) );
  XOR U1620 ( .A(n1770), .B(n1771), .Z(n1597) );
  AND U1621 ( .A(n108), .B(n1772), .Z(n1771) );
  XOR U1622 ( .A(p_input[860]), .B(p_input[844]), .Z(n1772) );
  XOR U1623 ( .A(n1773), .B(n1774), .Z(n1764) );
  AND U1624 ( .A(n1775), .B(n1776), .Z(n1774) );
  XOR U1625 ( .A(n1773), .B(n1612), .Z(n1776) );
  XNOR U1626 ( .A(p_input[875]), .B(n1777), .Z(n1612) );
  AND U1627 ( .A(n110), .B(n1778), .Z(n1777) );
  XOR U1628 ( .A(p_input[891]), .B(p_input[875]), .Z(n1778) );
  XNOR U1629 ( .A(n1609), .B(n1773), .Z(n1775) );
  XOR U1630 ( .A(n1779), .B(n1780), .Z(n1609) );
  AND U1631 ( .A(n108), .B(n1781), .Z(n1780) );
  XOR U1632 ( .A(p_input[859]), .B(p_input[843]), .Z(n1781) );
  XOR U1633 ( .A(n1782), .B(n1783), .Z(n1773) );
  AND U1634 ( .A(n1784), .B(n1785), .Z(n1783) );
  XOR U1635 ( .A(n1782), .B(n1624), .Z(n1785) );
  XNOR U1636 ( .A(p_input[874]), .B(n1786), .Z(n1624) );
  AND U1637 ( .A(n110), .B(n1787), .Z(n1786) );
  XOR U1638 ( .A(p_input[890]), .B(p_input[874]), .Z(n1787) );
  XNOR U1639 ( .A(n1621), .B(n1782), .Z(n1784) );
  XOR U1640 ( .A(n1788), .B(n1789), .Z(n1621) );
  AND U1641 ( .A(n108), .B(n1790), .Z(n1789) );
  XOR U1642 ( .A(p_input[858]), .B(p_input[842]), .Z(n1790) );
  XOR U1643 ( .A(n1791), .B(n1792), .Z(n1782) );
  AND U1644 ( .A(n1793), .B(n1794), .Z(n1792) );
  XOR U1645 ( .A(n1791), .B(n1636), .Z(n1794) );
  XNOR U1646 ( .A(p_input[873]), .B(n1795), .Z(n1636) );
  AND U1647 ( .A(n110), .B(n1796), .Z(n1795) );
  XOR U1648 ( .A(p_input[889]), .B(p_input[873]), .Z(n1796) );
  XNOR U1649 ( .A(n1633), .B(n1791), .Z(n1793) );
  XOR U1650 ( .A(n1797), .B(n1798), .Z(n1633) );
  AND U1651 ( .A(n108), .B(n1799), .Z(n1798) );
  XOR U1652 ( .A(p_input[857]), .B(p_input[841]), .Z(n1799) );
  XOR U1653 ( .A(n1800), .B(n1801), .Z(n1791) );
  AND U1654 ( .A(n1802), .B(n1803), .Z(n1801) );
  XOR U1655 ( .A(n1800), .B(n1648), .Z(n1803) );
  XNOR U1656 ( .A(p_input[872]), .B(n1804), .Z(n1648) );
  AND U1657 ( .A(n110), .B(n1805), .Z(n1804) );
  XOR U1658 ( .A(p_input[888]), .B(p_input[872]), .Z(n1805) );
  XNOR U1659 ( .A(n1645), .B(n1800), .Z(n1802) );
  XOR U1660 ( .A(n1806), .B(n1807), .Z(n1645) );
  AND U1661 ( .A(n108), .B(n1808), .Z(n1807) );
  XOR U1662 ( .A(p_input[856]), .B(p_input[840]), .Z(n1808) );
  XOR U1663 ( .A(n1809), .B(n1810), .Z(n1800) );
  AND U1664 ( .A(n1811), .B(n1812), .Z(n1810) );
  XOR U1665 ( .A(n1809), .B(n1660), .Z(n1812) );
  XNOR U1666 ( .A(p_input[871]), .B(n1813), .Z(n1660) );
  AND U1667 ( .A(n110), .B(n1814), .Z(n1813) );
  XOR U1668 ( .A(p_input[887]), .B(p_input[871]), .Z(n1814) );
  XNOR U1669 ( .A(n1657), .B(n1809), .Z(n1811) );
  XOR U1670 ( .A(n1815), .B(n1816), .Z(n1657) );
  AND U1671 ( .A(n108), .B(n1817), .Z(n1816) );
  XOR U1672 ( .A(p_input[855]), .B(p_input[839]), .Z(n1817) );
  XOR U1673 ( .A(n1818), .B(n1819), .Z(n1809) );
  AND U1674 ( .A(n1820), .B(n1821), .Z(n1819) );
  XOR U1675 ( .A(n1818), .B(n1672), .Z(n1821) );
  XNOR U1676 ( .A(p_input[870]), .B(n1822), .Z(n1672) );
  AND U1677 ( .A(n110), .B(n1823), .Z(n1822) );
  XOR U1678 ( .A(p_input[886]), .B(p_input[870]), .Z(n1823) );
  XNOR U1679 ( .A(n1669), .B(n1818), .Z(n1820) );
  XOR U1680 ( .A(n1824), .B(n1825), .Z(n1669) );
  AND U1681 ( .A(n108), .B(n1826), .Z(n1825) );
  XOR U1682 ( .A(p_input[854]), .B(p_input[838]), .Z(n1826) );
  XOR U1683 ( .A(n1827), .B(n1828), .Z(n1818) );
  AND U1684 ( .A(n1829), .B(n1830), .Z(n1828) );
  XOR U1685 ( .A(n1827), .B(n1684), .Z(n1830) );
  XNOR U1686 ( .A(p_input[869]), .B(n1831), .Z(n1684) );
  AND U1687 ( .A(n110), .B(n1832), .Z(n1831) );
  XOR U1688 ( .A(p_input[885]), .B(p_input[869]), .Z(n1832) );
  XNOR U1689 ( .A(n1681), .B(n1827), .Z(n1829) );
  XOR U1690 ( .A(n1833), .B(n1834), .Z(n1681) );
  AND U1691 ( .A(n108), .B(n1835), .Z(n1834) );
  XOR U1692 ( .A(p_input[853]), .B(p_input[837]), .Z(n1835) );
  XOR U1693 ( .A(n1836), .B(n1837), .Z(n1827) );
  AND U1694 ( .A(n1838), .B(n1839), .Z(n1837) );
  XOR U1695 ( .A(n1836), .B(n1696), .Z(n1839) );
  XNOR U1696 ( .A(p_input[868]), .B(n1840), .Z(n1696) );
  AND U1697 ( .A(n110), .B(n1841), .Z(n1840) );
  XOR U1698 ( .A(p_input[884]), .B(p_input[868]), .Z(n1841) );
  XNOR U1699 ( .A(n1693), .B(n1836), .Z(n1838) );
  XOR U1700 ( .A(n1842), .B(n1843), .Z(n1693) );
  AND U1701 ( .A(n108), .B(n1844), .Z(n1843) );
  XOR U1702 ( .A(p_input[852]), .B(p_input[836]), .Z(n1844) );
  XOR U1703 ( .A(n1845), .B(n1846), .Z(n1836) );
  AND U1704 ( .A(n1847), .B(n1848), .Z(n1846) );
  XOR U1705 ( .A(n1708), .B(n1845), .Z(n1848) );
  XNOR U1706 ( .A(p_input[867]), .B(n1849), .Z(n1708) );
  AND U1707 ( .A(n110), .B(n1850), .Z(n1849) );
  XOR U1708 ( .A(p_input[883]), .B(p_input[867]), .Z(n1850) );
  XNOR U1709 ( .A(n1845), .B(n1705), .Z(n1847) );
  XOR U1710 ( .A(n1851), .B(n1852), .Z(n1705) );
  AND U1711 ( .A(n108), .B(n1853), .Z(n1852) );
  XOR U1712 ( .A(p_input[851]), .B(p_input[835]), .Z(n1853) );
  XOR U1713 ( .A(n1854), .B(n1855), .Z(n1845) );
  AND U1714 ( .A(n1856), .B(n1857), .Z(n1855) );
  XOR U1715 ( .A(n1854), .B(n1720), .Z(n1857) );
  XNOR U1716 ( .A(p_input[866]), .B(n1858), .Z(n1720) );
  AND U1717 ( .A(n110), .B(n1859), .Z(n1858) );
  XOR U1718 ( .A(p_input[882]), .B(p_input[866]), .Z(n1859) );
  XNOR U1719 ( .A(n1717), .B(n1854), .Z(n1856) );
  XOR U1720 ( .A(n1860), .B(n1861), .Z(n1717) );
  AND U1721 ( .A(n108), .B(n1862), .Z(n1861) );
  XOR U1722 ( .A(p_input[850]), .B(p_input[834]), .Z(n1862) );
  XOR U1723 ( .A(n1863), .B(n1864), .Z(n1854) );
  AND U1724 ( .A(n1865), .B(n1866), .Z(n1864) );
  XNOR U1725 ( .A(n1867), .B(n1733), .Z(n1866) );
  XNOR U1726 ( .A(p_input[865]), .B(n1868), .Z(n1733) );
  AND U1727 ( .A(n110), .B(n1869), .Z(n1868) );
  XNOR U1728 ( .A(p_input[881]), .B(n1870), .Z(n1869) );
  IV U1729 ( .A(p_input[865]), .Z(n1870) );
  XNOR U1730 ( .A(n1730), .B(n1863), .Z(n1865) );
  XNOR U1731 ( .A(p_input[833]), .B(n1871), .Z(n1730) );
  AND U1732 ( .A(n108), .B(n1872), .Z(n1871) );
  XOR U1733 ( .A(p_input[849]), .B(p_input[833]), .Z(n1872) );
  IV U1734 ( .A(n1867), .Z(n1863) );
  AND U1735 ( .A(n1738), .B(n1741), .Z(n1867) );
  XOR U1736 ( .A(p_input[864]), .B(n1873), .Z(n1741) );
  AND U1737 ( .A(n110), .B(n1874), .Z(n1873) );
  XOR U1738 ( .A(p_input[880]), .B(p_input[864]), .Z(n1874) );
  XOR U1739 ( .A(n1875), .B(n1876), .Z(n110) );
  AND U1740 ( .A(n1877), .B(n1878), .Z(n1876) );
  XNOR U1741 ( .A(p_input[895]), .B(n1875), .Z(n1878) );
  XOR U1742 ( .A(n1875), .B(p_input[879]), .Z(n1877) );
  XOR U1743 ( .A(n1879), .B(n1880), .Z(n1875) );
  AND U1744 ( .A(n1881), .B(n1882), .Z(n1880) );
  XNOR U1745 ( .A(p_input[894]), .B(n1879), .Z(n1882) );
  XOR U1746 ( .A(n1879), .B(p_input[878]), .Z(n1881) );
  XOR U1747 ( .A(n1883), .B(n1884), .Z(n1879) );
  AND U1748 ( .A(n1885), .B(n1886), .Z(n1884) );
  XNOR U1749 ( .A(p_input[893]), .B(n1883), .Z(n1886) );
  XOR U1750 ( .A(n1883), .B(p_input[877]), .Z(n1885) );
  XOR U1751 ( .A(n1887), .B(n1888), .Z(n1883) );
  AND U1752 ( .A(n1889), .B(n1890), .Z(n1888) );
  XNOR U1753 ( .A(p_input[892]), .B(n1887), .Z(n1890) );
  XOR U1754 ( .A(n1887), .B(p_input[876]), .Z(n1889) );
  XOR U1755 ( .A(n1891), .B(n1892), .Z(n1887) );
  AND U1756 ( .A(n1893), .B(n1894), .Z(n1892) );
  XNOR U1757 ( .A(p_input[891]), .B(n1891), .Z(n1894) );
  XOR U1758 ( .A(n1891), .B(p_input[875]), .Z(n1893) );
  XOR U1759 ( .A(n1895), .B(n1896), .Z(n1891) );
  AND U1760 ( .A(n1897), .B(n1898), .Z(n1896) );
  XNOR U1761 ( .A(p_input[890]), .B(n1895), .Z(n1898) );
  XOR U1762 ( .A(n1895), .B(p_input[874]), .Z(n1897) );
  XOR U1763 ( .A(n1899), .B(n1900), .Z(n1895) );
  AND U1764 ( .A(n1901), .B(n1902), .Z(n1900) );
  XNOR U1765 ( .A(p_input[889]), .B(n1899), .Z(n1902) );
  XOR U1766 ( .A(n1899), .B(p_input[873]), .Z(n1901) );
  XOR U1767 ( .A(n1903), .B(n1904), .Z(n1899) );
  AND U1768 ( .A(n1905), .B(n1906), .Z(n1904) );
  XNOR U1769 ( .A(p_input[888]), .B(n1903), .Z(n1906) );
  XOR U1770 ( .A(n1903), .B(p_input[872]), .Z(n1905) );
  XOR U1771 ( .A(n1907), .B(n1908), .Z(n1903) );
  AND U1772 ( .A(n1909), .B(n1910), .Z(n1908) );
  XNOR U1773 ( .A(p_input[887]), .B(n1907), .Z(n1910) );
  XOR U1774 ( .A(n1907), .B(p_input[871]), .Z(n1909) );
  XOR U1775 ( .A(n1911), .B(n1912), .Z(n1907) );
  AND U1776 ( .A(n1913), .B(n1914), .Z(n1912) );
  XNOR U1777 ( .A(p_input[886]), .B(n1911), .Z(n1914) );
  XOR U1778 ( .A(n1911), .B(p_input[870]), .Z(n1913) );
  XOR U1779 ( .A(n1915), .B(n1916), .Z(n1911) );
  AND U1780 ( .A(n1917), .B(n1918), .Z(n1916) );
  XNOR U1781 ( .A(p_input[885]), .B(n1915), .Z(n1918) );
  XOR U1782 ( .A(n1915), .B(p_input[869]), .Z(n1917) );
  XOR U1783 ( .A(n1919), .B(n1920), .Z(n1915) );
  AND U1784 ( .A(n1921), .B(n1922), .Z(n1920) );
  XNOR U1785 ( .A(p_input[884]), .B(n1919), .Z(n1922) );
  XOR U1786 ( .A(n1919), .B(p_input[868]), .Z(n1921) );
  XOR U1787 ( .A(n1923), .B(n1924), .Z(n1919) );
  AND U1788 ( .A(n1925), .B(n1926), .Z(n1924) );
  XNOR U1789 ( .A(p_input[883]), .B(n1923), .Z(n1926) );
  XOR U1790 ( .A(n1923), .B(p_input[867]), .Z(n1925) );
  XOR U1791 ( .A(n1927), .B(n1928), .Z(n1923) );
  AND U1792 ( .A(n1929), .B(n1930), .Z(n1928) );
  XNOR U1793 ( .A(p_input[882]), .B(n1927), .Z(n1930) );
  XOR U1794 ( .A(n1927), .B(p_input[866]), .Z(n1929) );
  XNOR U1795 ( .A(n1931), .B(n1932), .Z(n1927) );
  AND U1796 ( .A(n1933), .B(n1934), .Z(n1932) );
  XOR U1797 ( .A(p_input[881]), .B(n1931), .Z(n1934) );
  XNOR U1798 ( .A(p_input[865]), .B(n1931), .Z(n1933) );
  AND U1799 ( .A(p_input[880]), .B(n1935), .Z(n1931) );
  IV U1800 ( .A(p_input[864]), .Z(n1935) );
  XNOR U1801 ( .A(p_input[832]), .B(n1936), .Z(n1738) );
  AND U1802 ( .A(n108), .B(n1937), .Z(n1936) );
  XOR U1803 ( .A(p_input[848]), .B(p_input[832]), .Z(n1937) );
  XOR U1804 ( .A(n1938), .B(n1939), .Z(n108) );
  AND U1805 ( .A(n1940), .B(n1941), .Z(n1939) );
  XNOR U1806 ( .A(p_input[863]), .B(n1938), .Z(n1941) );
  XOR U1807 ( .A(n1938), .B(p_input[847]), .Z(n1940) );
  XOR U1808 ( .A(n1942), .B(n1943), .Z(n1938) );
  AND U1809 ( .A(n1944), .B(n1945), .Z(n1943) );
  XNOR U1810 ( .A(p_input[862]), .B(n1942), .Z(n1945) );
  XNOR U1811 ( .A(n1942), .B(n1752), .Z(n1944) );
  IV U1812 ( .A(p_input[846]), .Z(n1752) );
  XOR U1813 ( .A(n1946), .B(n1947), .Z(n1942) );
  AND U1814 ( .A(n1948), .B(n1949), .Z(n1947) );
  XNOR U1815 ( .A(p_input[861]), .B(n1946), .Z(n1949) );
  XNOR U1816 ( .A(n1946), .B(n1761), .Z(n1948) );
  IV U1817 ( .A(p_input[845]), .Z(n1761) );
  XOR U1818 ( .A(n1950), .B(n1951), .Z(n1946) );
  AND U1819 ( .A(n1952), .B(n1953), .Z(n1951) );
  XNOR U1820 ( .A(p_input[860]), .B(n1950), .Z(n1953) );
  XNOR U1821 ( .A(n1950), .B(n1770), .Z(n1952) );
  IV U1822 ( .A(p_input[844]), .Z(n1770) );
  XOR U1823 ( .A(n1954), .B(n1955), .Z(n1950) );
  AND U1824 ( .A(n1956), .B(n1957), .Z(n1955) );
  XNOR U1825 ( .A(p_input[859]), .B(n1954), .Z(n1957) );
  XNOR U1826 ( .A(n1954), .B(n1779), .Z(n1956) );
  IV U1827 ( .A(p_input[843]), .Z(n1779) );
  XOR U1828 ( .A(n1958), .B(n1959), .Z(n1954) );
  AND U1829 ( .A(n1960), .B(n1961), .Z(n1959) );
  XNOR U1830 ( .A(p_input[858]), .B(n1958), .Z(n1961) );
  XNOR U1831 ( .A(n1958), .B(n1788), .Z(n1960) );
  IV U1832 ( .A(p_input[842]), .Z(n1788) );
  XOR U1833 ( .A(n1962), .B(n1963), .Z(n1958) );
  AND U1834 ( .A(n1964), .B(n1965), .Z(n1963) );
  XNOR U1835 ( .A(p_input[857]), .B(n1962), .Z(n1965) );
  XNOR U1836 ( .A(n1962), .B(n1797), .Z(n1964) );
  IV U1837 ( .A(p_input[841]), .Z(n1797) );
  XOR U1838 ( .A(n1966), .B(n1967), .Z(n1962) );
  AND U1839 ( .A(n1968), .B(n1969), .Z(n1967) );
  XNOR U1840 ( .A(p_input[856]), .B(n1966), .Z(n1969) );
  XNOR U1841 ( .A(n1966), .B(n1806), .Z(n1968) );
  IV U1842 ( .A(p_input[840]), .Z(n1806) );
  XOR U1843 ( .A(n1970), .B(n1971), .Z(n1966) );
  AND U1844 ( .A(n1972), .B(n1973), .Z(n1971) );
  XNOR U1845 ( .A(p_input[855]), .B(n1970), .Z(n1973) );
  XNOR U1846 ( .A(n1970), .B(n1815), .Z(n1972) );
  IV U1847 ( .A(p_input[839]), .Z(n1815) );
  XOR U1848 ( .A(n1974), .B(n1975), .Z(n1970) );
  AND U1849 ( .A(n1976), .B(n1977), .Z(n1975) );
  XNOR U1850 ( .A(p_input[854]), .B(n1974), .Z(n1977) );
  XNOR U1851 ( .A(n1974), .B(n1824), .Z(n1976) );
  IV U1852 ( .A(p_input[838]), .Z(n1824) );
  XOR U1853 ( .A(n1978), .B(n1979), .Z(n1974) );
  AND U1854 ( .A(n1980), .B(n1981), .Z(n1979) );
  XNOR U1855 ( .A(p_input[853]), .B(n1978), .Z(n1981) );
  XNOR U1856 ( .A(n1978), .B(n1833), .Z(n1980) );
  IV U1857 ( .A(p_input[837]), .Z(n1833) );
  XOR U1858 ( .A(n1982), .B(n1983), .Z(n1978) );
  AND U1859 ( .A(n1984), .B(n1985), .Z(n1983) );
  XNOR U1860 ( .A(p_input[852]), .B(n1982), .Z(n1985) );
  XNOR U1861 ( .A(n1982), .B(n1842), .Z(n1984) );
  IV U1862 ( .A(p_input[836]), .Z(n1842) );
  XOR U1863 ( .A(n1986), .B(n1987), .Z(n1982) );
  AND U1864 ( .A(n1988), .B(n1989), .Z(n1987) );
  XNOR U1865 ( .A(p_input[851]), .B(n1986), .Z(n1989) );
  XNOR U1866 ( .A(n1986), .B(n1851), .Z(n1988) );
  IV U1867 ( .A(p_input[835]), .Z(n1851) );
  XOR U1868 ( .A(n1990), .B(n1991), .Z(n1986) );
  AND U1869 ( .A(n1992), .B(n1993), .Z(n1991) );
  XNOR U1870 ( .A(p_input[850]), .B(n1990), .Z(n1993) );
  XNOR U1871 ( .A(n1990), .B(n1860), .Z(n1992) );
  IV U1872 ( .A(p_input[834]), .Z(n1860) );
  XNOR U1873 ( .A(n1994), .B(n1995), .Z(n1990) );
  AND U1874 ( .A(n1996), .B(n1997), .Z(n1995) );
  XOR U1875 ( .A(p_input[849]), .B(n1994), .Z(n1997) );
  XNOR U1876 ( .A(p_input[833]), .B(n1994), .Z(n1996) );
  AND U1877 ( .A(p_input[848]), .B(n1998), .Z(n1994) );
  IV U1878 ( .A(p_input[832]), .Z(n1998) );
  XOR U1879 ( .A(n1999), .B(n2000), .Z(n1557) );
  AND U1880 ( .A(n159), .B(n2001), .Z(n2000) );
  XNOR U1881 ( .A(n2002), .B(n1999), .Z(n2001) );
  XOR U1882 ( .A(n2003), .B(n2004), .Z(n159) );
  AND U1883 ( .A(n2005), .B(n2006), .Z(n2004) );
  XNOR U1884 ( .A(n1568), .B(n2003), .Z(n2006) );
  AND U1885 ( .A(p_input[831]), .B(p_input[815]), .Z(n1568) );
  XOR U1886 ( .A(n2003), .B(n1567), .Z(n2005) );
  AND U1887 ( .A(p_input[783]), .B(p_input[799]), .Z(n1567) );
  XOR U1888 ( .A(n2007), .B(n2008), .Z(n2003) );
  AND U1889 ( .A(n2009), .B(n2010), .Z(n2008) );
  XOR U1890 ( .A(n2007), .B(n1580), .Z(n2010) );
  XNOR U1891 ( .A(p_input[814]), .B(n2011), .Z(n1580) );
  AND U1892 ( .A(n114), .B(n2012), .Z(n2011) );
  XOR U1893 ( .A(p_input[830]), .B(p_input[814]), .Z(n2012) );
  XNOR U1894 ( .A(n1577), .B(n2007), .Z(n2009) );
  XOR U1895 ( .A(n2013), .B(n2014), .Z(n1577) );
  AND U1896 ( .A(n111), .B(n2015), .Z(n2014) );
  XOR U1897 ( .A(p_input[798]), .B(p_input[782]), .Z(n2015) );
  XOR U1898 ( .A(n2016), .B(n2017), .Z(n2007) );
  AND U1899 ( .A(n2018), .B(n2019), .Z(n2017) );
  XOR U1900 ( .A(n2016), .B(n1592), .Z(n2019) );
  XNOR U1901 ( .A(p_input[813]), .B(n2020), .Z(n1592) );
  AND U1902 ( .A(n114), .B(n2021), .Z(n2020) );
  XOR U1903 ( .A(p_input[829]), .B(p_input[813]), .Z(n2021) );
  XNOR U1904 ( .A(n1589), .B(n2016), .Z(n2018) );
  XOR U1905 ( .A(n2022), .B(n2023), .Z(n1589) );
  AND U1906 ( .A(n111), .B(n2024), .Z(n2023) );
  XOR U1907 ( .A(p_input[797]), .B(p_input[781]), .Z(n2024) );
  XOR U1908 ( .A(n2025), .B(n2026), .Z(n2016) );
  AND U1909 ( .A(n2027), .B(n2028), .Z(n2026) );
  XOR U1910 ( .A(n2025), .B(n1604), .Z(n2028) );
  XNOR U1911 ( .A(p_input[812]), .B(n2029), .Z(n1604) );
  AND U1912 ( .A(n114), .B(n2030), .Z(n2029) );
  XOR U1913 ( .A(p_input[828]), .B(p_input[812]), .Z(n2030) );
  XNOR U1914 ( .A(n1601), .B(n2025), .Z(n2027) );
  XOR U1915 ( .A(n2031), .B(n2032), .Z(n1601) );
  AND U1916 ( .A(n111), .B(n2033), .Z(n2032) );
  XOR U1917 ( .A(p_input[796]), .B(p_input[780]), .Z(n2033) );
  XOR U1918 ( .A(n2034), .B(n2035), .Z(n2025) );
  AND U1919 ( .A(n2036), .B(n2037), .Z(n2035) );
  XOR U1920 ( .A(n2034), .B(n1616), .Z(n2037) );
  XNOR U1921 ( .A(p_input[811]), .B(n2038), .Z(n1616) );
  AND U1922 ( .A(n114), .B(n2039), .Z(n2038) );
  XOR U1923 ( .A(p_input[827]), .B(p_input[811]), .Z(n2039) );
  XNOR U1924 ( .A(n1613), .B(n2034), .Z(n2036) );
  XOR U1925 ( .A(n2040), .B(n2041), .Z(n1613) );
  AND U1926 ( .A(n111), .B(n2042), .Z(n2041) );
  XOR U1927 ( .A(p_input[795]), .B(p_input[779]), .Z(n2042) );
  XOR U1928 ( .A(n2043), .B(n2044), .Z(n2034) );
  AND U1929 ( .A(n2045), .B(n2046), .Z(n2044) );
  XOR U1930 ( .A(n2043), .B(n1628), .Z(n2046) );
  XNOR U1931 ( .A(p_input[810]), .B(n2047), .Z(n1628) );
  AND U1932 ( .A(n114), .B(n2048), .Z(n2047) );
  XOR U1933 ( .A(p_input[826]), .B(p_input[810]), .Z(n2048) );
  XNOR U1934 ( .A(n1625), .B(n2043), .Z(n2045) );
  XOR U1935 ( .A(n2049), .B(n2050), .Z(n1625) );
  AND U1936 ( .A(n111), .B(n2051), .Z(n2050) );
  XOR U1937 ( .A(p_input[794]), .B(p_input[778]), .Z(n2051) );
  XOR U1938 ( .A(n2052), .B(n2053), .Z(n2043) );
  AND U1939 ( .A(n2054), .B(n2055), .Z(n2053) );
  XOR U1940 ( .A(n2052), .B(n1640), .Z(n2055) );
  XNOR U1941 ( .A(p_input[809]), .B(n2056), .Z(n1640) );
  AND U1942 ( .A(n114), .B(n2057), .Z(n2056) );
  XOR U1943 ( .A(p_input[825]), .B(p_input[809]), .Z(n2057) );
  XNOR U1944 ( .A(n1637), .B(n2052), .Z(n2054) );
  XOR U1945 ( .A(n2058), .B(n2059), .Z(n1637) );
  AND U1946 ( .A(n111), .B(n2060), .Z(n2059) );
  XOR U1947 ( .A(p_input[793]), .B(p_input[777]), .Z(n2060) );
  XOR U1948 ( .A(n2061), .B(n2062), .Z(n2052) );
  AND U1949 ( .A(n2063), .B(n2064), .Z(n2062) );
  XOR U1950 ( .A(n2061), .B(n1652), .Z(n2064) );
  XNOR U1951 ( .A(p_input[808]), .B(n2065), .Z(n1652) );
  AND U1952 ( .A(n114), .B(n2066), .Z(n2065) );
  XOR U1953 ( .A(p_input[824]), .B(p_input[808]), .Z(n2066) );
  XNOR U1954 ( .A(n1649), .B(n2061), .Z(n2063) );
  XOR U1955 ( .A(n2067), .B(n2068), .Z(n1649) );
  AND U1956 ( .A(n111), .B(n2069), .Z(n2068) );
  XOR U1957 ( .A(p_input[792]), .B(p_input[776]), .Z(n2069) );
  XOR U1958 ( .A(n2070), .B(n2071), .Z(n2061) );
  AND U1959 ( .A(n2072), .B(n2073), .Z(n2071) );
  XOR U1960 ( .A(n2070), .B(n1664), .Z(n2073) );
  XNOR U1961 ( .A(p_input[807]), .B(n2074), .Z(n1664) );
  AND U1962 ( .A(n114), .B(n2075), .Z(n2074) );
  XOR U1963 ( .A(p_input[823]), .B(p_input[807]), .Z(n2075) );
  XNOR U1964 ( .A(n1661), .B(n2070), .Z(n2072) );
  XOR U1965 ( .A(n2076), .B(n2077), .Z(n1661) );
  AND U1966 ( .A(n111), .B(n2078), .Z(n2077) );
  XOR U1967 ( .A(p_input[791]), .B(p_input[775]), .Z(n2078) );
  XOR U1968 ( .A(n2079), .B(n2080), .Z(n2070) );
  AND U1969 ( .A(n2081), .B(n2082), .Z(n2080) );
  XOR U1970 ( .A(n2079), .B(n1676), .Z(n2082) );
  XNOR U1971 ( .A(p_input[806]), .B(n2083), .Z(n1676) );
  AND U1972 ( .A(n114), .B(n2084), .Z(n2083) );
  XOR U1973 ( .A(p_input[822]), .B(p_input[806]), .Z(n2084) );
  XNOR U1974 ( .A(n1673), .B(n2079), .Z(n2081) );
  XOR U1975 ( .A(n2085), .B(n2086), .Z(n1673) );
  AND U1976 ( .A(n111), .B(n2087), .Z(n2086) );
  XOR U1977 ( .A(p_input[790]), .B(p_input[774]), .Z(n2087) );
  XOR U1978 ( .A(n2088), .B(n2089), .Z(n2079) );
  AND U1979 ( .A(n2090), .B(n2091), .Z(n2089) );
  XOR U1980 ( .A(n2088), .B(n1688), .Z(n2091) );
  XNOR U1981 ( .A(p_input[805]), .B(n2092), .Z(n1688) );
  AND U1982 ( .A(n114), .B(n2093), .Z(n2092) );
  XOR U1983 ( .A(p_input[821]), .B(p_input[805]), .Z(n2093) );
  XNOR U1984 ( .A(n1685), .B(n2088), .Z(n2090) );
  XOR U1985 ( .A(n2094), .B(n2095), .Z(n1685) );
  AND U1986 ( .A(n111), .B(n2096), .Z(n2095) );
  XOR U1987 ( .A(p_input[789]), .B(p_input[773]), .Z(n2096) );
  XOR U1988 ( .A(n2097), .B(n2098), .Z(n2088) );
  AND U1989 ( .A(n2099), .B(n2100), .Z(n2098) );
  XOR U1990 ( .A(n2097), .B(n1700), .Z(n2100) );
  XNOR U1991 ( .A(p_input[804]), .B(n2101), .Z(n1700) );
  AND U1992 ( .A(n114), .B(n2102), .Z(n2101) );
  XOR U1993 ( .A(p_input[820]), .B(p_input[804]), .Z(n2102) );
  XNOR U1994 ( .A(n1697), .B(n2097), .Z(n2099) );
  XOR U1995 ( .A(n2103), .B(n2104), .Z(n1697) );
  AND U1996 ( .A(n111), .B(n2105), .Z(n2104) );
  XOR U1997 ( .A(p_input[788]), .B(p_input[772]), .Z(n2105) );
  XOR U1998 ( .A(n2106), .B(n2107), .Z(n2097) );
  AND U1999 ( .A(n2108), .B(n2109), .Z(n2107) );
  XOR U2000 ( .A(n1712), .B(n2106), .Z(n2109) );
  XNOR U2001 ( .A(p_input[803]), .B(n2110), .Z(n1712) );
  AND U2002 ( .A(n114), .B(n2111), .Z(n2110) );
  XOR U2003 ( .A(p_input[819]), .B(p_input[803]), .Z(n2111) );
  XNOR U2004 ( .A(n2106), .B(n1709), .Z(n2108) );
  XOR U2005 ( .A(n2112), .B(n2113), .Z(n1709) );
  AND U2006 ( .A(n111), .B(n2114), .Z(n2113) );
  XOR U2007 ( .A(p_input[787]), .B(p_input[771]), .Z(n2114) );
  XOR U2008 ( .A(n2115), .B(n2116), .Z(n2106) );
  AND U2009 ( .A(n2117), .B(n2118), .Z(n2116) );
  XOR U2010 ( .A(n2115), .B(n1724), .Z(n2118) );
  XNOR U2011 ( .A(p_input[802]), .B(n2119), .Z(n1724) );
  AND U2012 ( .A(n114), .B(n2120), .Z(n2119) );
  XOR U2013 ( .A(p_input[818]), .B(p_input[802]), .Z(n2120) );
  XNOR U2014 ( .A(n1721), .B(n2115), .Z(n2117) );
  XOR U2015 ( .A(n2121), .B(n2122), .Z(n1721) );
  AND U2016 ( .A(n111), .B(n2123), .Z(n2122) );
  XOR U2017 ( .A(p_input[786]), .B(p_input[770]), .Z(n2123) );
  XOR U2018 ( .A(n2124), .B(n2125), .Z(n2115) );
  AND U2019 ( .A(n2126), .B(n2127), .Z(n2125) );
  XNOR U2020 ( .A(n2128), .B(n1737), .Z(n2127) );
  XNOR U2021 ( .A(p_input[801]), .B(n2129), .Z(n1737) );
  AND U2022 ( .A(n114), .B(n2130), .Z(n2129) );
  XNOR U2023 ( .A(p_input[817]), .B(n2131), .Z(n2130) );
  IV U2024 ( .A(p_input[801]), .Z(n2131) );
  XNOR U2025 ( .A(n1734), .B(n2124), .Z(n2126) );
  XNOR U2026 ( .A(p_input[769]), .B(n2132), .Z(n1734) );
  AND U2027 ( .A(n111), .B(n2133), .Z(n2132) );
  XOR U2028 ( .A(p_input[785]), .B(p_input[769]), .Z(n2133) );
  IV U2029 ( .A(n2128), .Z(n2124) );
  AND U2030 ( .A(n1999), .B(n2002), .Z(n2128) );
  XOR U2031 ( .A(p_input[800]), .B(n2134), .Z(n2002) );
  AND U2032 ( .A(n114), .B(n2135), .Z(n2134) );
  XOR U2033 ( .A(p_input[816]), .B(p_input[800]), .Z(n2135) );
  XOR U2034 ( .A(n2136), .B(n2137), .Z(n114) );
  AND U2035 ( .A(n2138), .B(n2139), .Z(n2137) );
  XNOR U2036 ( .A(p_input[831]), .B(n2136), .Z(n2139) );
  XOR U2037 ( .A(n2136), .B(p_input[815]), .Z(n2138) );
  XOR U2038 ( .A(n2140), .B(n2141), .Z(n2136) );
  AND U2039 ( .A(n2142), .B(n2143), .Z(n2141) );
  XNOR U2040 ( .A(p_input[830]), .B(n2140), .Z(n2143) );
  XOR U2041 ( .A(n2140), .B(p_input[814]), .Z(n2142) );
  XOR U2042 ( .A(n2144), .B(n2145), .Z(n2140) );
  AND U2043 ( .A(n2146), .B(n2147), .Z(n2145) );
  XNOR U2044 ( .A(p_input[829]), .B(n2144), .Z(n2147) );
  XOR U2045 ( .A(n2144), .B(p_input[813]), .Z(n2146) );
  XOR U2046 ( .A(n2148), .B(n2149), .Z(n2144) );
  AND U2047 ( .A(n2150), .B(n2151), .Z(n2149) );
  XNOR U2048 ( .A(p_input[828]), .B(n2148), .Z(n2151) );
  XOR U2049 ( .A(n2148), .B(p_input[812]), .Z(n2150) );
  XOR U2050 ( .A(n2152), .B(n2153), .Z(n2148) );
  AND U2051 ( .A(n2154), .B(n2155), .Z(n2153) );
  XNOR U2052 ( .A(p_input[827]), .B(n2152), .Z(n2155) );
  XOR U2053 ( .A(n2152), .B(p_input[811]), .Z(n2154) );
  XOR U2054 ( .A(n2156), .B(n2157), .Z(n2152) );
  AND U2055 ( .A(n2158), .B(n2159), .Z(n2157) );
  XNOR U2056 ( .A(p_input[826]), .B(n2156), .Z(n2159) );
  XOR U2057 ( .A(n2156), .B(p_input[810]), .Z(n2158) );
  XOR U2058 ( .A(n2160), .B(n2161), .Z(n2156) );
  AND U2059 ( .A(n2162), .B(n2163), .Z(n2161) );
  XNOR U2060 ( .A(p_input[825]), .B(n2160), .Z(n2163) );
  XOR U2061 ( .A(n2160), .B(p_input[809]), .Z(n2162) );
  XOR U2062 ( .A(n2164), .B(n2165), .Z(n2160) );
  AND U2063 ( .A(n2166), .B(n2167), .Z(n2165) );
  XNOR U2064 ( .A(p_input[824]), .B(n2164), .Z(n2167) );
  XOR U2065 ( .A(n2164), .B(p_input[808]), .Z(n2166) );
  XOR U2066 ( .A(n2168), .B(n2169), .Z(n2164) );
  AND U2067 ( .A(n2170), .B(n2171), .Z(n2169) );
  XNOR U2068 ( .A(p_input[823]), .B(n2168), .Z(n2171) );
  XOR U2069 ( .A(n2168), .B(p_input[807]), .Z(n2170) );
  XOR U2070 ( .A(n2172), .B(n2173), .Z(n2168) );
  AND U2071 ( .A(n2174), .B(n2175), .Z(n2173) );
  XNOR U2072 ( .A(p_input[822]), .B(n2172), .Z(n2175) );
  XOR U2073 ( .A(n2172), .B(p_input[806]), .Z(n2174) );
  XOR U2074 ( .A(n2176), .B(n2177), .Z(n2172) );
  AND U2075 ( .A(n2178), .B(n2179), .Z(n2177) );
  XNOR U2076 ( .A(p_input[821]), .B(n2176), .Z(n2179) );
  XOR U2077 ( .A(n2176), .B(p_input[805]), .Z(n2178) );
  XOR U2078 ( .A(n2180), .B(n2181), .Z(n2176) );
  AND U2079 ( .A(n2182), .B(n2183), .Z(n2181) );
  XNOR U2080 ( .A(p_input[820]), .B(n2180), .Z(n2183) );
  XOR U2081 ( .A(n2180), .B(p_input[804]), .Z(n2182) );
  XOR U2082 ( .A(n2184), .B(n2185), .Z(n2180) );
  AND U2083 ( .A(n2186), .B(n2187), .Z(n2185) );
  XNOR U2084 ( .A(p_input[819]), .B(n2184), .Z(n2187) );
  XOR U2085 ( .A(n2184), .B(p_input[803]), .Z(n2186) );
  XOR U2086 ( .A(n2188), .B(n2189), .Z(n2184) );
  AND U2087 ( .A(n2190), .B(n2191), .Z(n2189) );
  XNOR U2088 ( .A(p_input[818]), .B(n2188), .Z(n2191) );
  XOR U2089 ( .A(n2188), .B(p_input[802]), .Z(n2190) );
  XNOR U2090 ( .A(n2192), .B(n2193), .Z(n2188) );
  AND U2091 ( .A(n2194), .B(n2195), .Z(n2193) );
  XOR U2092 ( .A(p_input[817]), .B(n2192), .Z(n2195) );
  XNOR U2093 ( .A(p_input[801]), .B(n2192), .Z(n2194) );
  AND U2094 ( .A(p_input[816]), .B(n2196), .Z(n2192) );
  IV U2095 ( .A(p_input[800]), .Z(n2196) );
  XNOR U2096 ( .A(p_input[768]), .B(n2197), .Z(n1999) );
  AND U2097 ( .A(n111), .B(n2198), .Z(n2197) );
  XOR U2098 ( .A(p_input[784]), .B(p_input[768]), .Z(n2198) );
  XOR U2099 ( .A(n2199), .B(n2200), .Z(n111) );
  AND U2100 ( .A(n2201), .B(n2202), .Z(n2200) );
  XNOR U2101 ( .A(p_input[799]), .B(n2199), .Z(n2202) );
  XOR U2102 ( .A(n2199), .B(p_input[783]), .Z(n2201) );
  XOR U2103 ( .A(n2203), .B(n2204), .Z(n2199) );
  AND U2104 ( .A(n2205), .B(n2206), .Z(n2204) );
  XNOR U2105 ( .A(p_input[798]), .B(n2203), .Z(n2206) );
  XNOR U2106 ( .A(n2203), .B(n2013), .Z(n2205) );
  IV U2107 ( .A(p_input[782]), .Z(n2013) );
  XOR U2108 ( .A(n2207), .B(n2208), .Z(n2203) );
  AND U2109 ( .A(n2209), .B(n2210), .Z(n2208) );
  XNOR U2110 ( .A(p_input[797]), .B(n2207), .Z(n2210) );
  XNOR U2111 ( .A(n2207), .B(n2022), .Z(n2209) );
  IV U2112 ( .A(p_input[781]), .Z(n2022) );
  XOR U2113 ( .A(n2211), .B(n2212), .Z(n2207) );
  AND U2114 ( .A(n2213), .B(n2214), .Z(n2212) );
  XNOR U2115 ( .A(p_input[796]), .B(n2211), .Z(n2214) );
  XNOR U2116 ( .A(n2211), .B(n2031), .Z(n2213) );
  IV U2117 ( .A(p_input[780]), .Z(n2031) );
  XOR U2118 ( .A(n2215), .B(n2216), .Z(n2211) );
  AND U2119 ( .A(n2217), .B(n2218), .Z(n2216) );
  XNOR U2120 ( .A(p_input[795]), .B(n2215), .Z(n2218) );
  XNOR U2121 ( .A(n2215), .B(n2040), .Z(n2217) );
  IV U2122 ( .A(p_input[779]), .Z(n2040) );
  XOR U2123 ( .A(n2219), .B(n2220), .Z(n2215) );
  AND U2124 ( .A(n2221), .B(n2222), .Z(n2220) );
  XNOR U2125 ( .A(p_input[794]), .B(n2219), .Z(n2222) );
  XNOR U2126 ( .A(n2219), .B(n2049), .Z(n2221) );
  IV U2127 ( .A(p_input[778]), .Z(n2049) );
  XOR U2128 ( .A(n2223), .B(n2224), .Z(n2219) );
  AND U2129 ( .A(n2225), .B(n2226), .Z(n2224) );
  XNOR U2130 ( .A(p_input[793]), .B(n2223), .Z(n2226) );
  XNOR U2131 ( .A(n2223), .B(n2058), .Z(n2225) );
  IV U2132 ( .A(p_input[777]), .Z(n2058) );
  XOR U2133 ( .A(n2227), .B(n2228), .Z(n2223) );
  AND U2134 ( .A(n2229), .B(n2230), .Z(n2228) );
  XNOR U2135 ( .A(p_input[792]), .B(n2227), .Z(n2230) );
  XNOR U2136 ( .A(n2227), .B(n2067), .Z(n2229) );
  IV U2137 ( .A(p_input[776]), .Z(n2067) );
  XOR U2138 ( .A(n2231), .B(n2232), .Z(n2227) );
  AND U2139 ( .A(n2233), .B(n2234), .Z(n2232) );
  XNOR U2140 ( .A(p_input[791]), .B(n2231), .Z(n2234) );
  XNOR U2141 ( .A(n2231), .B(n2076), .Z(n2233) );
  IV U2142 ( .A(p_input[775]), .Z(n2076) );
  XOR U2143 ( .A(n2235), .B(n2236), .Z(n2231) );
  AND U2144 ( .A(n2237), .B(n2238), .Z(n2236) );
  XNOR U2145 ( .A(p_input[790]), .B(n2235), .Z(n2238) );
  XNOR U2146 ( .A(n2235), .B(n2085), .Z(n2237) );
  IV U2147 ( .A(p_input[774]), .Z(n2085) );
  XOR U2148 ( .A(n2239), .B(n2240), .Z(n2235) );
  AND U2149 ( .A(n2241), .B(n2242), .Z(n2240) );
  XNOR U2150 ( .A(p_input[789]), .B(n2239), .Z(n2242) );
  XNOR U2151 ( .A(n2239), .B(n2094), .Z(n2241) );
  IV U2152 ( .A(p_input[773]), .Z(n2094) );
  XOR U2153 ( .A(n2243), .B(n2244), .Z(n2239) );
  AND U2154 ( .A(n2245), .B(n2246), .Z(n2244) );
  XNOR U2155 ( .A(p_input[788]), .B(n2243), .Z(n2246) );
  XNOR U2156 ( .A(n2243), .B(n2103), .Z(n2245) );
  IV U2157 ( .A(p_input[772]), .Z(n2103) );
  XOR U2158 ( .A(n2247), .B(n2248), .Z(n2243) );
  AND U2159 ( .A(n2249), .B(n2250), .Z(n2248) );
  XNOR U2160 ( .A(p_input[787]), .B(n2247), .Z(n2250) );
  XNOR U2161 ( .A(n2247), .B(n2112), .Z(n2249) );
  IV U2162 ( .A(p_input[771]), .Z(n2112) );
  XOR U2163 ( .A(n2251), .B(n2252), .Z(n2247) );
  AND U2164 ( .A(n2253), .B(n2254), .Z(n2252) );
  XNOR U2165 ( .A(p_input[786]), .B(n2251), .Z(n2254) );
  XNOR U2166 ( .A(n2251), .B(n2121), .Z(n2253) );
  IV U2167 ( .A(p_input[770]), .Z(n2121) );
  XNOR U2168 ( .A(n2255), .B(n2256), .Z(n2251) );
  AND U2169 ( .A(n2257), .B(n2258), .Z(n2256) );
  XOR U2170 ( .A(p_input[785]), .B(n2255), .Z(n2258) );
  XNOR U2171 ( .A(p_input[769]), .B(n2255), .Z(n2257) );
  AND U2172 ( .A(p_input[784]), .B(n2259), .Z(n2255) );
  IV U2173 ( .A(p_input[768]), .Z(n2259) );
  XOR U2174 ( .A(n2260), .B(n2261), .Z(n487) );
  AND U2175 ( .A(n284), .B(n2262), .Z(n2261) );
  XNOR U2176 ( .A(n2263), .B(n2260), .Z(n2262) );
  XOR U2177 ( .A(n2264), .B(n2265), .Z(n284) );
  AND U2178 ( .A(n2266), .B(n2267), .Z(n2265) );
  XNOR U2179 ( .A(n502), .B(n2264), .Z(n2267) );
  AND U2180 ( .A(n2268), .B(n2269), .Z(n502) );
  XNOR U2181 ( .A(n2264), .B(n499), .Z(n2266) );
  IV U2182 ( .A(n2270), .Z(n499) );
  AND U2183 ( .A(n2271), .B(n2272), .Z(n2270) );
  XOR U2184 ( .A(n2273), .B(n2274), .Z(n2264) );
  AND U2185 ( .A(n2275), .B(n2276), .Z(n2274) );
  XOR U2186 ( .A(n2273), .B(n514), .Z(n2276) );
  XOR U2187 ( .A(n2277), .B(n2278), .Z(n514) );
  AND U2188 ( .A(n250), .B(n2279), .Z(n2278) );
  XOR U2189 ( .A(n2280), .B(n2277), .Z(n2279) );
  XNOR U2190 ( .A(n511), .B(n2273), .Z(n2275) );
  XOR U2191 ( .A(n2281), .B(n2282), .Z(n511) );
  AND U2192 ( .A(n247), .B(n2283), .Z(n2282) );
  XOR U2193 ( .A(n2284), .B(n2281), .Z(n2283) );
  XOR U2194 ( .A(n2285), .B(n2286), .Z(n2273) );
  AND U2195 ( .A(n2287), .B(n2288), .Z(n2286) );
  XOR U2196 ( .A(n2285), .B(n526), .Z(n2288) );
  XOR U2197 ( .A(n2289), .B(n2290), .Z(n526) );
  AND U2198 ( .A(n250), .B(n2291), .Z(n2290) );
  XOR U2199 ( .A(n2292), .B(n2289), .Z(n2291) );
  XNOR U2200 ( .A(n523), .B(n2285), .Z(n2287) );
  XOR U2201 ( .A(n2293), .B(n2294), .Z(n523) );
  AND U2202 ( .A(n247), .B(n2295), .Z(n2294) );
  XOR U2203 ( .A(n2296), .B(n2293), .Z(n2295) );
  XOR U2204 ( .A(n2297), .B(n2298), .Z(n2285) );
  AND U2205 ( .A(n2299), .B(n2300), .Z(n2298) );
  XOR U2206 ( .A(n2297), .B(n538), .Z(n2300) );
  XOR U2207 ( .A(n2301), .B(n2302), .Z(n538) );
  AND U2208 ( .A(n250), .B(n2303), .Z(n2302) );
  XOR U2209 ( .A(n2304), .B(n2301), .Z(n2303) );
  XNOR U2210 ( .A(n535), .B(n2297), .Z(n2299) );
  XOR U2211 ( .A(n2305), .B(n2306), .Z(n535) );
  AND U2212 ( .A(n247), .B(n2307), .Z(n2306) );
  XOR U2213 ( .A(n2308), .B(n2305), .Z(n2307) );
  XOR U2214 ( .A(n2309), .B(n2310), .Z(n2297) );
  AND U2215 ( .A(n2311), .B(n2312), .Z(n2310) );
  XOR U2216 ( .A(n2309), .B(n550), .Z(n2312) );
  XOR U2217 ( .A(n2313), .B(n2314), .Z(n550) );
  AND U2218 ( .A(n250), .B(n2315), .Z(n2314) );
  XOR U2219 ( .A(n2316), .B(n2313), .Z(n2315) );
  XNOR U2220 ( .A(n547), .B(n2309), .Z(n2311) );
  XOR U2221 ( .A(n2317), .B(n2318), .Z(n547) );
  AND U2222 ( .A(n247), .B(n2319), .Z(n2318) );
  XOR U2223 ( .A(n2320), .B(n2317), .Z(n2319) );
  XOR U2224 ( .A(n2321), .B(n2322), .Z(n2309) );
  AND U2225 ( .A(n2323), .B(n2324), .Z(n2322) );
  XOR U2226 ( .A(n2321), .B(n562), .Z(n2324) );
  XOR U2227 ( .A(n2325), .B(n2326), .Z(n562) );
  AND U2228 ( .A(n250), .B(n2327), .Z(n2326) );
  XOR U2229 ( .A(n2328), .B(n2325), .Z(n2327) );
  XNOR U2230 ( .A(n559), .B(n2321), .Z(n2323) );
  XOR U2231 ( .A(n2329), .B(n2330), .Z(n559) );
  AND U2232 ( .A(n247), .B(n2331), .Z(n2330) );
  XOR U2233 ( .A(n2332), .B(n2329), .Z(n2331) );
  XOR U2234 ( .A(n2333), .B(n2334), .Z(n2321) );
  AND U2235 ( .A(n2335), .B(n2336), .Z(n2334) );
  XOR U2236 ( .A(n2333), .B(n574), .Z(n2336) );
  XOR U2237 ( .A(n2337), .B(n2338), .Z(n574) );
  AND U2238 ( .A(n250), .B(n2339), .Z(n2338) );
  XOR U2239 ( .A(n2340), .B(n2337), .Z(n2339) );
  XNOR U2240 ( .A(n571), .B(n2333), .Z(n2335) );
  XOR U2241 ( .A(n2341), .B(n2342), .Z(n571) );
  AND U2242 ( .A(n247), .B(n2343), .Z(n2342) );
  XOR U2243 ( .A(n2344), .B(n2341), .Z(n2343) );
  XOR U2244 ( .A(n2345), .B(n2346), .Z(n2333) );
  AND U2245 ( .A(n2347), .B(n2348), .Z(n2346) );
  XOR U2246 ( .A(n2345), .B(n586), .Z(n2348) );
  XOR U2247 ( .A(n2349), .B(n2350), .Z(n586) );
  AND U2248 ( .A(n250), .B(n2351), .Z(n2350) );
  XOR U2249 ( .A(n2352), .B(n2349), .Z(n2351) );
  XNOR U2250 ( .A(n583), .B(n2345), .Z(n2347) );
  XOR U2251 ( .A(n2353), .B(n2354), .Z(n583) );
  AND U2252 ( .A(n247), .B(n2355), .Z(n2354) );
  XOR U2253 ( .A(n2356), .B(n2353), .Z(n2355) );
  XOR U2254 ( .A(n2357), .B(n2358), .Z(n2345) );
  AND U2255 ( .A(n2359), .B(n2360), .Z(n2358) );
  XOR U2256 ( .A(n2357), .B(n598), .Z(n2360) );
  XOR U2257 ( .A(n2361), .B(n2362), .Z(n598) );
  AND U2258 ( .A(n250), .B(n2363), .Z(n2362) );
  XOR U2259 ( .A(n2364), .B(n2361), .Z(n2363) );
  XNOR U2260 ( .A(n595), .B(n2357), .Z(n2359) );
  XOR U2261 ( .A(n2365), .B(n2366), .Z(n595) );
  AND U2262 ( .A(n247), .B(n2367), .Z(n2366) );
  XOR U2263 ( .A(n2368), .B(n2365), .Z(n2367) );
  XOR U2264 ( .A(n2369), .B(n2370), .Z(n2357) );
  AND U2265 ( .A(n2371), .B(n2372), .Z(n2370) );
  XOR U2266 ( .A(n2369), .B(n610), .Z(n2372) );
  XOR U2267 ( .A(n2373), .B(n2374), .Z(n610) );
  AND U2268 ( .A(n250), .B(n2375), .Z(n2374) );
  XOR U2269 ( .A(n2376), .B(n2373), .Z(n2375) );
  XNOR U2270 ( .A(n607), .B(n2369), .Z(n2371) );
  XOR U2271 ( .A(n2377), .B(n2378), .Z(n607) );
  AND U2272 ( .A(n247), .B(n2379), .Z(n2378) );
  XOR U2273 ( .A(n2380), .B(n2377), .Z(n2379) );
  XOR U2274 ( .A(n2381), .B(n2382), .Z(n2369) );
  AND U2275 ( .A(n2383), .B(n2384), .Z(n2382) );
  XOR U2276 ( .A(n2381), .B(n622), .Z(n2384) );
  XOR U2277 ( .A(n2385), .B(n2386), .Z(n622) );
  AND U2278 ( .A(n250), .B(n2387), .Z(n2386) );
  XOR U2279 ( .A(n2388), .B(n2385), .Z(n2387) );
  XNOR U2280 ( .A(n619), .B(n2381), .Z(n2383) );
  XOR U2281 ( .A(n2389), .B(n2390), .Z(n619) );
  AND U2282 ( .A(n247), .B(n2391), .Z(n2390) );
  XOR U2283 ( .A(n2392), .B(n2389), .Z(n2391) );
  XOR U2284 ( .A(n2393), .B(n2394), .Z(n2381) );
  AND U2285 ( .A(n2395), .B(n2396), .Z(n2394) );
  XOR U2286 ( .A(n2393), .B(n634), .Z(n2396) );
  XOR U2287 ( .A(n2397), .B(n2398), .Z(n634) );
  AND U2288 ( .A(n250), .B(n2399), .Z(n2398) );
  XOR U2289 ( .A(n2400), .B(n2397), .Z(n2399) );
  XNOR U2290 ( .A(n631), .B(n2393), .Z(n2395) );
  XOR U2291 ( .A(n2401), .B(n2402), .Z(n631) );
  AND U2292 ( .A(n247), .B(n2403), .Z(n2402) );
  XOR U2293 ( .A(n2404), .B(n2401), .Z(n2403) );
  XOR U2294 ( .A(n2405), .B(n2406), .Z(n2393) );
  AND U2295 ( .A(n2407), .B(n2408), .Z(n2406) );
  XOR U2296 ( .A(n646), .B(n2405), .Z(n2408) );
  XOR U2297 ( .A(n2409), .B(n2410), .Z(n646) );
  AND U2298 ( .A(n250), .B(n2411), .Z(n2410) );
  XOR U2299 ( .A(n2409), .B(n2412), .Z(n2411) );
  XNOR U2300 ( .A(n2405), .B(n643), .Z(n2407) );
  XOR U2301 ( .A(n2413), .B(n2414), .Z(n643) );
  AND U2302 ( .A(n247), .B(n2415), .Z(n2414) );
  XOR U2303 ( .A(n2413), .B(n2416), .Z(n2415) );
  XOR U2304 ( .A(n2417), .B(n2418), .Z(n2405) );
  AND U2305 ( .A(n2419), .B(n2420), .Z(n2418) );
  XOR U2306 ( .A(n2417), .B(n658), .Z(n2420) );
  XOR U2307 ( .A(n2421), .B(n2422), .Z(n658) );
  AND U2308 ( .A(n250), .B(n2423), .Z(n2422) );
  XOR U2309 ( .A(n2424), .B(n2421), .Z(n2423) );
  XNOR U2310 ( .A(n655), .B(n2417), .Z(n2419) );
  XOR U2311 ( .A(n2425), .B(n2426), .Z(n655) );
  AND U2312 ( .A(n247), .B(n2427), .Z(n2426) );
  XOR U2313 ( .A(n2428), .B(n2425), .Z(n2427) );
  XOR U2314 ( .A(n2429), .B(n2430), .Z(n2417) );
  AND U2315 ( .A(n2431), .B(n2432), .Z(n2430) );
  XNOR U2316 ( .A(n2433), .B(n671), .Z(n2432) );
  XOR U2317 ( .A(n2434), .B(n2435), .Z(n671) );
  AND U2318 ( .A(n250), .B(n2436), .Z(n2435) );
  XOR U2319 ( .A(n2437), .B(n2434), .Z(n2436) );
  XNOR U2320 ( .A(n668), .B(n2429), .Z(n2431) );
  XOR U2321 ( .A(n2438), .B(n2439), .Z(n668) );
  AND U2322 ( .A(n247), .B(n2440), .Z(n2439) );
  XOR U2323 ( .A(n2441), .B(n2438), .Z(n2440) );
  IV U2324 ( .A(n2433), .Z(n2429) );
  AND U2325 ( .A(n2260), .B(n2263), .Z(n2433) );
  XNOR U2326 ( .A(n2442), .B(n2443), .Z(n2263) );
  AND U2327 ( .A(n250), .B(n2444), .Z(n2443) );
  XNOR U2328 ( .A(n2445), .B(n2442), .Z(n2444) );
  XOR U2329 ( .A(n2446), .B(n2447), .Z(n250) );
  AND U2330 ( .A(n2448), .B(n2449), .Z(n2447) );
  XNOR U2331 ( .A(n2268), .B(n2446), .Z(n2449) );
  AND U2332 ( .A(n2450), .B(n2451), .Z(n2268) );
  XOR U2333 ( .A(n2446), .B(n2269), .Z(n2448) );
  AND U2334 ( .A(n2452), .B(n2453), .Z(n2269) );
  XOR U2335 ( .A(n2454), .B(n2455), .Z(n2446) );
  AND U2336 ( .A(n2456), .B(n2457), .Z(n2455) );
  XOR U2337 ( .A(n2454), .B(n2280), .Z(n2457) );
  XOR U2338 ( .A(n2458), .B(n2459), .Z(n2280) );
  AND U2339 ( .A(n170), .B(n2460), .Z(n2459) );
  XOR U2340 ( .A(n2461), .B(n2458), .Z(n2460) );
  XNOR U2341 ( .A(n2277), .B(n2454), .Z(n2456) );
  XOR U2342 ( .A(n2462), .B(n2463), .Z(n2277) );
  AND U2343 ( .A(n168), .B(n2464), .Z(n2463) );
  XOR U2344 ( .A(n2465), .B(n2462), .Z(n2464) );
  XOR U2345 ( .A(n2466), .B(n2467), .Z(n2454) );
  AND U2346 ( .A(n2468), .B(n2469), .Z(n2467) );
  XOR U2347 ( .A(n2466), .B(n2292), .Z(n2469) );
  XOR U2348 ( .A(n2470), .B(n2471), .Z(n2292) );
  AND U2349 ( .A(n170), .B(n2472), .Z(n2471) );
  XOR U2350 ( .A(n2473), .B(n2470), .Z(n2472) );
  XNOR U2351 ( .A(n2289), .B(n2466), .Z(n2468) );
  XOR U2352 ( .A(n2474), .B(n2475), .Z(n2289) );
  AND U2353 ( .A(n168), .B(n2476), .Z(n2475) );
  XOR U2354 ( .A(n2477), .B(n2474), .Z(n2476) );
  XOR U2355 ( .A(n2478), .B(n2479), .Z(n2466) );
  AND U2356 ( .A(n2480), .B(n2481), .Z(n2479) );
  XOR U2357 ( .A(n2478), .B(n2304), .Z(n2481) );
  XOR U2358 ( .A(n2482), .B(n2483), .Z(n2304) );
  AND U2359 ( .A(n170), .B(n2484), .Z(n2483) );
  XOR U2360 ( .A(n2485), .B(n2482), .Z(n2484) );
  XNOR U2361 ( .A(n2301), .B(n2478), .Z(n2480) );
  XOR U2362 ( .A(n2486), .B(n2487), .Z(n2301) );
  AND U2363 ( .A(n168), .B(n2488), .Z(n2487) );
  XOR U2364 ( .A(n2489), .B(n2486), .Z(n2488) );
  XOR U2365 ( .A(n2490), .B(n2491), .Z(n2478) );
  AND U2366 ( .A(n2492), .B(n2493), .Z(n2491) );
  XOR U2367 ( .A(n2490), .B(n2316), .Z(n2493) );
  XOR U2368 ( .A(n2494), .B(n2495), .Z(n2316) );
  AND U2369 ( .A(n170), .B(n2496), .Z(n2495) );
  XOR U2370 ( .A(n2497), .B(n2494), .Z(n2496) );
  XNOR U2371 ( .A(n2313), .B(n2490), .Z(n2492) );
  XOR U2372 ( .A(n2498), .B(n2499), .Z(n2313) );
  AND U2373 ( .A(n168), .B(n2500), .Z(n2499) );
  XOR U2374 ( .A(n2501), .B(n2498), .Z(n2500) );
  XOR U2375 ( .A(n2502), .B(n2503), .Z(n2490) );
  AND U2376 ( .A(n2504), .B(n2505), .Z(n2503) );
  XOR U2377 ( .A(n2502), .B(n2328), .Z(n2505) );
  XOR U2378 ( .A(n2506), .B(n2507), .Z(n2328) );
  AND U2379 ( .A(n170), .B(n2508), .Z(n2507) );
  XOR U2380 ( .A(n2509), .B(n2506), .Z(n2508) );
  XNOR U2381 ( .A(n2325), .B(n2502), .Z(n2504) );
  XOR U2382 ( .A(n2510), .B(n2511), .Z(n2325) );
  AND U2383 ( .A(n168), .B(n2512), .Z(n2511) );
  XOR U2384 ( .A(n2513), .B(n2510), .Z(n2512) );
  XOR U2385 ( .A(n2514), .B(n2515), .Z(n2502) );
  AND U2386 ( .A(n2516), .B(n2517), .Z(n2515) );
  XOR U2387 ( .A(n2514), .B(n2340), .Z(n2517) );
  XOR U2388 ( .A(n2518), .B(n2519), .Z(n2340) );
  AND U2389 ( .A(n170), .B(n2520), .Z(n2519) );
  XOR U2390 ( .A(n2521), .B(n2518), .Z(n2520) );
  XNOR U2391 ( .A(n2337), .B(n2514), .Z(n2516) );
  XOR U2392 ( .A(n2522), .B(n2523), .Z(n2337) );
  AND U2393 ( .A(n168), .B(n2524), .Z(n2523) );
  XOR U2394 ( .A(n2525), .B(n2522), .Z(n2524) );
  XOR U2395 ( .A(n2526), .B(n2527), .Z(n2514) );
  AND U2396 ( .A(n2528), .B(n2529), .Z(n2527) );
  XOR U2397 ( .A(n2526), .B(n2352), .Z(n2529) );
  XOR U2398 ( .A(n2530), .B(n2531), .Z(n2352) );
  AND U2399 ( .A(n170), .B(n2532), .Z(n2531) );
  XOR U2400 ( .A(n2533), .B(n2530), .Z(n2532) );
  XNOR U2401 ( .A(n2349), .B(n2526), .Z(n2528) );
  XOR U2402 ( .A(n2534), .B(n2535), .Z(n2349) );
  AND U2403 ( .A(n168), .B(n2536), .Z(n2535) );
  XOR U2404 ( .A(n2537), .B(n2534), .Z(n2536) );
  XOR U2405 ( .A(n2538), .B(n2539), .Z(n2526) );
  AND U2406 ( .A(n2540), .B(n2541), .Z(n2539) );
  XOR U2407 ( .A(n2538), .B(n2364), .Z(n2541) );
  XOR U2408 ( .A(n2542), .B(n2543), .Z(n2364) );
  AND U2409 ( .A(n170), .B(n2544), .Z(n2543) );
  XOR U2410 ( .A(n2545), .B(n2542), .Z(n2544) );
  XNOR U2411 ( .A(n2361), .B(n2538), .Z(n2540) );
  XOR U2412 ( .A(n2546), .B(n2547), .Z(n2361) );
  AND U2413 ( .A(n168), .B(n2548), .Z(n2547) );
  XOR U2414 ( .A(n2549), .B(n2546), .Z(n2548) );
  XOR U2415 ( .A(n2550), .B(n2551), .Z(n2538) );
  AND U2416 ( .A(n2552), .B(n2553), .Z(n2551) );
  XOR U2417 ( .A(n2550), .B(n2376), .Z(n2553) );
  XOR U2418 ( .A(n2554), .B(n2555), .Z(n2376) );
  AND U2419 ( .A(n170), .B(n2556), .Z(n2555) );
  XOR U2420 ( .A(n2557), .B(n2554), .Z(n2556) );
  XNOR U2421 ( .A(n2373), .B(n2550), .Z(n2552) );
  XOR U2422 ( .A(n2558), .B(n2559), .Z(n2373) );
  AND U2423 ( .A(n168), .B(n2560), .Z(n2559) );
  XOR U2424 ( .A(n2561), .B(n2558), .Z(n2560) );
  XOR U2425 ( .A(n2562), .B(n2563), .Z(n2550) );
  AND U2426 ( .A(n2564), .B(n2565), .Z(n2563) );
  XOR U2427 ( .A(n2562), .B(n2388), .Z(n2565) );
  XOR U2428 ( .A(n2566), .B(n2567), .Z(n2388) );
  AND U2429 ( .A(n170), .B(n2568), .Z(n2567) );
  XOR U2430 ( .A(n2569), .B(n2566), .Z(n2568) );
  XNOR U2431 ( .A(n2385), .B(n2562), .Z(n2564) );
  XOR U2432 ( .A(n2570), .B(n2571), .Z(n2385) );
  AND U2433 ( .A(n168), .B(n2572), .Z(n2571) );
  XOR U2434 ( .A(n2573), .B(n2570), .Z(n2572) );
  XOR U2435 ( .A(n2574), .B(n2575), .Z(n2562) );
  AND U2436 ( .A(n2576), .B(n2577), .Z(n2575) );
  XOR U2437 ( .A(n2574), .B(n2400), .Z(n2577) );
  XOR U2438 ( .A(n2578), .B(n2579), .Z(n2400) );
  AND U2439 ( .A(n170), .B(n2580), .Z(n2579) );
  XOR U2440 ( .A(n2581), .B(n2578), .Z(n2580) );
  XNOR U2441 ( .A(n2397), .B(n2574), .Z(n2576) );
  XOR U2442 ( .A(n2582), .B(n2583), .Z(n2397) );
  AND U2443 ( .A(n168), .B(n2584), .Z(n2583) );
  XOR U2444 ( .A(n2585), .B(n2582), .Z(n2584) );
  XOR U2445 ( .A(n2586), .B(n2587), .Z(n2574) );
  AND U2446 ( .A(n2588), .B(n2589), .Z(n2587) );
  XOR U2447 ( .A(n2412), .B(n2586), .Z(n2589) );
  XOR U2448 ( .A(n2590), .B(n2591), .Z(n2412) );
  AND U2449 ( .A(n170), .B(n2592), .Z(n2591) );
  XOR U2450 ( .A(n2590), .B(n2593), .Z(n2592) );
  XNOR U2451 ( .A(n2586), .B(n2409), .Z(n2588) );
  XOR U2452 ( .A(n2594), .B(n2595), .Z(n2409) );
  AND U2453 ( .A(n168), .B(n2596), .Z(n2595) );
  XOR U2454 ( .A(n2594), .B(n2597), .Z(n2596) );
  XOR U2455 ( .A(n2598), .B(n2599), .Z(n2586) );
  AND U2456 ( .A(n2600), .B(n2601), .Z(n2599) );
  XOR U2457 ( .A(n2598), .B(n2424), .Z(n2601) );
  XOR U2458 ( .A(n2602), .B(n2603), .Z(n2424) );
  AND U2459 ( .A(n170), .B(n2604), .Z(n2603) );
  XOR U2460 ( .A(n2605), .B(n2602), .Z(n2604) );
  XNOR U2461 ( .A(n2421), .B(n2598), .Z(n2600) );
  XOR U2462 ( .A(n2606), .B(n2607), .Z(n2421) );
  AND U2463 ( .A(n168), .B(n2608), .Z(n2607) );
  XOR U2464 ( .A(n2609), .B(n2606), .Z(n2608) );
  XOR U2465 ( .A(n2610), .B(n2611), .Z(n2598) );
  AND U2466 ( .A(n2612), .B(n2613), .Z(n2611) );
  XNOR U2467 ( .A(n2614), .B(n2437), .Z(n2613) );
  XOR U2468 ( .A(n2615), .B(n2616), .Z(n2437) );
  AND U2469 ( .A(n170), .B(n2617), .Z(n2616) );
  XOR U2470 ( .A(n2618), .B(n2615), .Z(n2617) );
  XNOR U2471 ( .A(n2434), .B(n2610), .Z(n2612) );
  XOR U2472 ( .A(n2619), .B(n2620), .Z(n2434) );
  AND U2473 ( .A(n168), .B(n2621), .Z(n2620) );
  XOR U2474 ( .A(n2622), .B(n2619), .Z(n2621) );
  IV U2475 ( .A(n2614), .Z(n2610) );
  AND U2476 ( .A(n2442), .B(n2445), .Z(n2614) );
  XNOR U2477 ( .A(n2623), .B(n2624), .Z(n2445) );
  AND U2478 ( .A(n170), .B(n2625), .Z(n2624) );
  XNOR U2479 ( .A(n2626), .B(n2623), .Z(n2625) );
  XOR U2480 ( .A(n2627), .B(n2628), .Z(n170) );
  AND U2481 ( .A(n2629), .B(n2630), .Z(n2628) );
  XNOR U2482 ( .A(n2450), .B(n2627), .Z(n2630) );
  AND U2483 ( .A(p_input[767]), .B(p_input[751]), .Z(n2450) );
  XOR U2484 ( .A(n2627), .B(n2451), .Z(n2629) );
  AND U2485 ( .A(p_input[735]), .B(p_input[719]), .Z(n2451) );
  XOR U2486 ( .A(n2631), .B(n2632), .Z(n2627) );
  AND U2487 ( .A(n2633), .B(n2634), .Z(n2632) );
  XOR U2488 ( .A(n2631), .B(n2461), .Z(n2634) );
  XNOR U2489 ( .A(p_input[750]), .B(n2635), .Z(n2461) );
  AND U2490 ( .A(n126), .B(n2636), .Z(n2635) );
  XOR U2491 ( .A(p_input[766]), .B(p_input[750]), .Z(n2636) );
  XNOR U2492 ( .A(n2458), .B(n2631), .Z(n2633) );
  XOR U2493 ( .A(n2637), .B(n2638), .Z(n2458) );
  AND U2494 ( .A(n124), .B(n2639), .Z(n2638) );
  XOR U2495 ( .A(p_input[734]), .B(p_input[718]), .Z(n2639) );
  XOR U2496 ( .A(n2640), .B(n2641), .Z(n2631) );
  AND U2497 ( .A(n2642), .B(n2643), .Z(n2641) );
  XOR U2498 ( .A(n2640), .B(n2473), .Z(n2643) );
  XNOR U2499 ( .A(p_input[749]), .B(n2644), .Z(n2473) );
  AND U2500 ( .A(n126), .B(n2645), .Z(n2644) );
  XOR U2501 ( .A(p_input[765]), .B(p_input[749]), .Z(n2645) );
  XNOR U2502 ( .A(n2470), .B(n2640), .Z(n2642) );
  XOR U2503 ( .A(n2646), .B(n2647), .Z(n2470) );
  AND U2504 ( .A(n124), .B(n2648), .Z(n2647) );
  XOR U2505 ( .A(p_input[733]), .B(p_input[717]), .Z(n2648) );
  XOR U2506 ( .A(n2649), .B(n2650), .Z(n2640) );
  AND U2507 ( .A(n2651), .B(n2652), .Z(n2650) );
  XOR U2508 ( .A(n2649), .B(n2485), .Z(n2652) );
  XNOR U2509 ( .A(p_input[748]), .B(n2653), .Z(n2485) );
  AND U2510 ( .A(n126), .B(n2654), .Z(n2653) );
  XOR U2511 ( .A(p_input[764]), .B(p_input[748]), .Z(n2654) );
  XNOR U2512 ( .A(n2482), .B(n2649), .Z(n2651) );
  XOR U2513 ( .A(n2655), .B(n2656), .Z(n2482) );
  AND U2514 ( .A(n124), .B(n2657), .Z(n2656) );
  XOR U2515 ( .A(p_input[732]), .B(p_input[716]), .Z(n2657) );
  XOR U2516 ( .A(n2658), .B(n2659), .Z(n2649) );
  AND U2517 ( .A(n2660), .B(n2661), .Z(n2659) );
  XOR U2518 ( .A(n2658), .B(n2497), .Z(n2661) );
  XNOR U2519 ( .A(p_input[747]), .B(n2662), .Z(n2497) );
  AND U2520 ( .A(n126), .B(n2663), .Z(n2662) );
  XOR U2521 ( .A(p_input[763]), .B(p_input[747]), .Z(n2663) );
  XNOR U2522 ( .A(n2494), .B(n2658), .Z(n2660) );
  XOR U2523 ( .A(n2664), .B(n2665), .Z(n2494) );
  AND U2524 ( .A(n124), .B(n2666), .Z(n2665) );
  XOR U2525 ( .A(p_input[731]), .B(p_input[715]), .Z(n2666) );
  XOR U2526 ( .A(n2667), .B(n2668), .Z(n2658) );
  AND U2527 ( .A(n2669), .B(n2670), .Z(n2668) );
  XOR U2528 ( .A(n2667), .B(n2509), .Z(n2670) );
  XNOR U2529 ( .A(p_input[746]), .B(n2671), .Z(n2509) );
  AND U2530 ( .A(n126), .B(n2672), .Z(n2671) );
  XOR U2531 ( .A(p_input[762]), .B(p_input[746]), .Z(n2672) );
  XNOR U2532 ( .A(n2506), .B(n2667), .Z(n2669) );
  XOR U2533 ( .A(n2673), .B(n2674), .Z(n2506) );
  AND U2534 ( .A(n124), .B(n2675), .Z(n2674) );
  XOR U2535 ( .A(p_input[730]), .B(p_input[714]), .Z(n2675) );
  XOR U2536 ( .A(n2676), .B(n2677), .Z(n2667) );
  AND U2537 ( .A(n2678), .B(n2679), .Z(n2677) );
  XOR U2538 ( .A(n2676), .B(n2521), .Z(n2679) );
  XNOR U2539 ( .A(p_input[745]), .B(n2680), .Z(n2521) );
  AND U2540 ( .A(n126), .B(n2681), .Z(n2680) );
  XOR U2541 ( .A(p_input[761]), .B(p_input[745]), .Z(n2681) );
  XNOR U2542 ( .A(n2518), .B(n2676), .Z(n2678) );
  XOR U2543 ( .A(n2682), .B(n2683), .Z(n2518) );
  AND U2544 ( .A(n124), .B(n2684), .Z(n2683) );
  XOR U2545 ( .A(p_input[729]), .B(p_input[713]), .Z(n2684) );
  XOR U2546 ( .A(n2685), .B(n2686), .Z(n2676) );
  AND U2547 ( .A(n2687), .B(n2688), .Z(n2686) );
  XOR U2548 ( .A(n2685), .B(n2533), .Z(n2688) );
  XNOR U2549 ( .A(p_input[744]), .B(n2689), .Z(n2533) );
  AND U2550 ( .A(n126), .B(n2690), .Z(n2689) );
  XOR U2551 ( .A(p_input[760]), .B(p_input[744]), .Z(n2690) );
  XNOR U2552 ( .A(n2530), .B(n2685), .Z(n2687) );
  XOR U2553 ( .A(n2691), .B(n2692), .Z(n2530) );
  AND U2554 ( .A(n124), .B(n2693), .Z(n2692) );
  XOR U2555 ( .A(p_input[728]), .B(p_input[712]), .Z(n2693) );
  XOR U2556 ( .A(n2694), .B(n2695), .Z(n2685) );
  AND U2557 ( .A(n2696), .B(n2697), .Z(n2695) );
  XOR U2558 ( .A(n2694), .B(n2545), .Z(n2697) );
  XNOR U2559 ( .A(p_input[743]), .B(n2698), .Z(n2545) );
  AND U2560 ( .A(n126), .B(n2699), .Z(n2698) );
  XOR U2561 ( .A(p_input[759]), .B(p_input[743]), .Z(n2699) );
  XNOR U2562 ( .A(n2542), .B(n2694), .Z(n2696) );
  XOR U2563 ( .A(n2700), .B(n2701), .Z(n2542) );
  AND U2564 ( .A(n124), .B(n2702), .Z(n2701) );
  XOR U2565 ( .A(p_input[727]), .B(p_input[711]), .Z(n2702) );
  XOR U2566 ( .A(n2703), .B(n2704), .Z(n2694) );
  AND U2567 ( .A(n2705), .B(n2706), .Z(n2704) );
  XOR U2568 ( .A(n2703), .B(n2557), .Z(n2706) );
  XNOR U2569 ( .A(p_input[742]), .B(n2707), .Z(n2557) );
  AND U2570 ( .A(n126), .B(n2708), .Z(n2707) );
  XOR U2571 ( .A(p_input[758]), .B(p_input[742]), .Z(n2708) );
  XNOR U2572 ( .A(n2554), .B(n2703), .Z(n2705) );
  XOR U2573 ( .A(n2709), .B(n2710), .Z(n2554) );
  AND U2574 ( .A(n124), .B(n2711), .Z(n2710) );
  XOR U2575 ( .A(p_input[726]), .B(p_input[710]), .Z(n2711) );
  XOR U2576 ( .A(n2712), .B(n2713), .Z(n2703) );
  AND U2577 ( .A(n2714), .B(n2715), .Z(n2713) );
  XOR U2578 ( .A(n2712), .B(n2569), .Z(n2715) );
  XNOR U2579 ( .A(p_input[741]), .B(n2716), .Z(n2569) );
  AND U2580 ( .A(n126), .B(n2717), .Z(n2716) );
  XOR U2581 ( .A(p_input[757]), .B(p_input[741]), .Z(n2717) );
  XNOR U2582 ( .A(n2566), .B(n2712), .Z(n2714) );
  XOR U2583 ( .A(n2718), .B(n2719), .Z(n2566) );
  AND U2584 ( .A(n124), .B(n2720), .Z(n2719) );
  XOR U2585 ( .A(p_input[725]), .B(p_input[709]), .Z(n2720) );
  XOR U2586 ( .A(n2721), .B(n2722), .Z(n2712) );
  AND U2587 ( .A(n2723), .B(n2724), .Z(n2722) );
  XOR U2588 ( .A(n2721), .B(n2581), .Z(n2724) );
  XNOR U2589 ( .A(p_input[740]), .B(n2725), .Z(n2581) );
  AND U2590 ( .A(n126), .B(n2726), .Z(n2725) );
  XOR U2591 ( .A(p_input[756]), .B(p_input[740]), .Z(n2726) );
  XNOR U2592 ( .A(n2578), .B(n2721), .Z(n2723) );
  XOR U2593 ( .A(n2727), .B(n2728), .Z(n2578) );
  AND U2594 ( .A(n124), .B(n2729), .Z(n2728) );
  XOR U2595 ( .A(p_input[724]), .B(p_input[708]), .Z(n2729) );
  XOR U2596 ( .A(n2730), .B(n2731), .Z(n2721) );
  AND U2597 ( .A(n2732), .B(n2733), .Z(n2731) );
  XOR U2598 ( .A(n2593), .B(n2730), .Z(n2733) );
  XNOR U2599 ( .A(p_input[739]), .B(n2734), .Z(n2593) );
  AND U2600 ( .A(n126), .B(n2735), .Z(n2734) );
  XOR U2601 ( .A(p_input[755]), .B(p_input[739]), .Z(n2735) );
  XNOR U2602 ( .A(n2730), .B(n2590), .Z(n2732) );
  XOR U2603 ( .A(n2736), .B(n2737), .Z(n2590) );
  AND U2604 ( .A(n124), .B(n2738), .Z(n2737) );
  XOR U2605 ( .A(p_input[723]), .B(p_input[707]), .Z(n2738) );
  XOR U2606 ( .A(n2739), .B(n2740), .Z(n2730) );
  AND U2607 ( .A(n2741), .B(n2742), .Z(n2740) );
  XOR U2608 ( .A(n2739), .B(n2605), .Z(n2742) );
  XNOR U2609 ( .A(p_input[738]), .B(n2743), .Z(n2605) );
  AND U2610 ( .A(n126), .B(n2744), .Z(n2743) );
  XOR U2611 ( .A(p_input[754]), .B(p_input[738]), .Z(n2744) );
  XNOR U2612 ( .A(n2602), .B(n2739), .Z(n2741) );
  XOR U2613 ( .A(n2745), .B(n2746), .Z(n2602) );
  AND U2614 ( .A(n124), .B(n2747), .Z(n2746) );
  XOR U2615 ( .A(p_input[722]), .B(p_input[706]), .Z(n2747) );
  XOR U2616 ( .A(n2748), .B(n2749), .Z(n2739) );
  AND U2617 ( .A(n2750), .B(n2751), .Z(n2749) );
  XNOR U2618 ( .A(n2752), .B(n2618), .Z(n2751) );
  XNOR U2619 ( .A(p_input[737]), .B(n2753), .Z(n2618) );
  AND U2620 ( .A(n126), .B(n2754), .Z(n2753) );
  XNOR U2621 ( .A(p_input[753]), .B(n2755), .Z(n2754) );
  IV U2622 ( .A(p_input[737]), .Z(n2755) );
  XNOR U2623 ( .A(n2615), .B(n2748), .Z(n2750) );
  XNOR U2624 ( .A(p_input[705]), .B(n2756), .Z(n2615) );
  AND U2625 ( .A(n124), .B(n2757), .Z(n2756) );
  XOR U2626 ( .A(p_input[721]), .B(p_input[705]), .Z(n2757) );
  IV U2627 ( .A(n2752), .Z(n2748) );
  AND U2628 ( .A(n2623), .B(n2626), .Z(n2752) );
  XOR U2629 ( .A(p_input[736]), .B(n2758), .Z(n2626) );
  AND U2630 ( .A(n126), .B(n2759), .Z(n2758) );
  XOR U2631 ( .A(p_input[752]), .B(p_input[736]), .Z(n2759) );
  XOR U2632 ( .A(n2760), .B(n2761), .Z(n126) );
  AND U2633 ( .A(n2762), .B(n2763), .Z(n2761) );
  XNOR U2634 ( .A(p_input[767]), .B(n2760), .Z(n2763) );
  XOR U2635 ( .A(n2760), .B(p_input[751]), .Z(n2762) );
  XOR U2636 ( .A(n2764), .B(n2765), .Z(n2760) );
  AND U2637 ( .A(n2766), .B(n2767), .Z(n2765) );
  XNOR U2638 ( .A(p_input[766]), .B(n2764), .Z(n2767) );
  XOR U2639 ( .A(n2764), .B(p_input[750]), .Z(n2766) );
  XOR U2640 ( .A(n2768), .B(n2769), .Z(n2764) );
  AND U2641 ( .A(n2770), .B(n2771), .Z(n2769) );
  XNOR U2642 ( .A(p_input[765]), .B(n2768), .Z(n2771) );
  XOR U2643 ( .A(n2768), .B(p_input[749]), .Z(n2770) );
  XOR U2644 ( .A(n2772), .B(n2773), .Z(n2768) );
  AND U2645 ( .A(n2774), .B(n2775), .Z(n2773) );
  XNOR U2646 ( .A(p_input[764]), .B(n2772), .Z(n2775) );
  XOR U2647 ( .A(n2772), .B(p_input[748]), .Z(n2774) );
  XOR U2648 ( .A(n2776), .B(n2777), .Z(n2772) );
  AND U2649 ( .A(n2778), .B(n2779), .Z(n2777) );
  XNOR U2650 ( .A(p_input[763]), .B(n2776), .Z(n2779) );
  XOR U2651 ( .A(n2776), .B(p_input[747]), .Z(n2778) );
  XOR U2652 ( .A(n2780), .B(n2781), .Z(n2776) );
  AND U2653 ( .A(n2782), .B(n2783), .Z(n2781) );
  XNOR U2654 ( .A(p_input[762]), .B(n2780), .Z(n2783) );
  XOR U2655 ( .A(n2780), .B(p_input[746]), .Z(n2782) );
  XOR U2656 ( .A(n2784), .B(n2785), .Z(n2780) );
  AND U2657 ( .A(n2786), .B(n2787), .Z(n2785) );
  XNOR U2658 ( .A(p_input[761]), .B(n2784), .Z(n2787) );
  XOR U2659 ( .A(n2784), .B(p_input[745]), .Z(n2786) );
  XOR U2660 ( .A(n2788), .B(n2789), .Z(n2784) );
  AND U2661 ( .A(n2790), .B(n2791), .Z(n2789) );
  XNOR U2662 ( .A(p_input[760]), .B(n2788), .Z(n2791) );
  XOR U2663 ( .A(n2788), .B(p_input[744]), .Z(n2790) );
  XOR U2664 ( .A(n2792), .B(n2793), .Z(n2788) );
  AND U2665 ( .A(n2794), .B(n2795), .Z(n2793) );
  XNOR U2666 ( .A(p_input[759]), .B(n2792), .Z(n2795) );
  XOR U2667 ( .A(n2792), .B(p_input[743]), .Z(n2794) );
  XOR U2668 ( .A(n2796), .B(n2797), .Z(n2792) );
  AND U2669 ( .A(n2798), .B(n2799), .Z(n2797) );
  XNOR U2670 ( .A(p_input[758]), .B(n2796), .Z(n2799) );
  XOR U2671 ( .A(n2796), .B(p_input[742]), .Z(n2798) );
  XOR U2672 ( .A(n2800), .B(n2801), .Z(n2796) );
  AND U2673 ( .A(n2802), .B(n2803), .Z(n2801) );
  XNOR U2674 ( .A(p_input[757]), .B(n2800), .Z(n2803) );
  XOR U2675 ( .A(n2800), .B(p_input[741]), .Z(n2802) );
  XOR U2676 ( .A(n2804), .B(n2805), .Z(n2800) );
  AND U2677 ( .A(n2806), .B(n2807), .Z(n2805) );
  XNOR U2678 ( .A(p_input[756]), .B(n2804), .Z(n2807) );
  XOR U2679 ( .A(n2804), .B(p_input[740]), .Z(n2806) );
  XOR U2680 ( .A(n2808), .B(n2809), .Z(n2804) );
  AND U2681 ( .A(n2810), .B(n2811), .Z(n2809) );
  XNOR U2682 ( .A(p_input[755]), .B(n2808), .Z(n2811) );
  XOR U2683 ( .A(n2808), .B(p_input[739]), .Z(n2810) );
  XOR U2684 ( .A(n2812), .B(n2813), .Z(n2808) );
  AND U2685 ( .A(n2814), .B(n2815), .Z(n2813) );
  XNOR U2686 ( .A(p_input[754]), .B(n2812), .Z(n2815) );
  XOR U2687 ( .A(n2812), .B(p_input[738]), .Z(n2814) );
  XNOR U2688 ( .A(n2816), .B(n2817), .Z(n2812) );
  AND U2689 ( .A(n2818), .B(n2819), .Z(n2817) );
  XOR U2690 ( .A(p_input[753]), .B(n2816), .Z(n2819) );
  XNOR U2691 ( .A(p_input[737]), .B(n2816), .Z(n2818) );
  AND U2692 ( .A(p_input[752]), .B(n2820), .Z(n2816) );
  IV U2693 ( .A(p_input[736]), .Z(n2820) );
  XNOR U2694 ( .A(p_input[704]), .B(n2821), .Z(n2623) );
  AND U2695 ( .A(n124), .B(n2822), .Z(n2821) );
  XOR U2696 ( .A(p_input[720]), .B(p_input[704]), .Z(n2822) );
  XOR U2697 ( .A(n2823), .B(n2824), .Z(n124) );
  AND U2698 ( .A(n2825), .B(n2826), .Z(n2824) );
  XNOR U2699 ( .A(p_input[735]), .B(n2823), .Z(n2826) );
  XOR U2700 ( .A(n2823), .B(p_input[719]), .Z(n2825) );
  XOR U2701 ( .A(n2827), .B(n2828), .Z(n2823) );
  AND U2702 ( .A(n2829), .B(n2830), .Z(n2828) );
  XNOR U2703 ( .A(p_input[734]), .B(n2827), .Z(n2830) );
  XNOR U2704 ( .A(n2827), .B(n2637), .Z(n2829) );
  IV U2705 ( .A(p_input[718]), .Z(n2637) );
  XOR U2706 ( .A(n2831), .B(n2832), .Z(n2827) );
  AND U2707 ( .A(n2833), .B(n2834), .Z(n2832) );
  XNOR U2708 ( .A(p_input[733]), .B(n2831), .Z(n2834) );
  XNOR U2709 ( .A(n2831), .B(n2646), .Z(n2833) );
  IV U2710 ( .A(p_input[717]), .Z(n2646) );
  XOR U2711 ( .A(n2835), .B(n2836), .Z(n2831) );
  AND U2712 ( .A(n2837), .B(n2838), .Z(n2836) );
  XNOR U2713 ( .A(p_input[732]), .B(n2835), .Z(n2838) );
  XNOR U2714 ( .A(n2835), .B(n2655), .Z(n2837) );
  IV U2715 ( .A(p_input[716]), .Z(n2655) );
  XOR U2716 ( .A(n2839), .B(n2840), .Z(n2835) );
  AND U2717 ( .A(n2841), .B(n2842), .Z(n2840) );
  XNOR U2718 ( .A(p_input[731]), .B(n2839), .Z(n2842) );
  XNOR U2719 ( .A(n2839), .B(n2664), .Z(n2841) );
  IV U2720 ( .A(p_input[715]), .Z(n2664) );
  XOR U2721 ( .A(n2843), .B(n2844), .Z(n2839) );
  AND U2722 ( .A(n2845), .B(n2846), .Z(n2844) );
  XNOR U2723 ( .A(p_input[730]), .B(n2843), .Z(n2846) );
  XNOR U2724 ( .A(n2843), .B(n2673), .Z(n2845) );
  IV U2725 ( .A(p_input[714]), .Z(n2673) );
  XOR U2726 ( .A(n2847), .B(n2848), .Z(n2843) );
  AND U2727 ( .A(n2849), .B(n2850), .Z(n2848) );
  XNOR U2728 ( .A(p_input[729]), .B(n2847), .Z(n2850) );
  XNOR U2729 ( .A(n2847), .B(n2682), .Z(n2849) );
  IV U2730 ( .A(p_input[713]), .Z(n2682) );
  XOR U2731 ( .A(n2851), .B(n2852), .Z(n2847) );
  AND U2732 ( .A(n2853), .B(n2854), .Z(n2852) );
  XNOR U2733 ( .A(p_input[728]), .B(n2851), .Z(n2854) );
  XNOR U2734 ( .A(n2851), .B(n2691), .Z(n2853) );
  IV U2735 ( .A(p_input[712]), .Z(n2691) );
  XOR U2736 ( .A(n2855), .B(n2856), .Z(n2851) );
  AND U2737 ( .A(n2857), .B(n2858), .Z(n2856) );
  XNOR U2738 ( .A(p_input[727]), .B(n2855), .Z(n2858) );
  XNOR U2739 ( .A(n2855), .B(n2700), .Z(n2857) );
  IV U2740 ( .A(p_input[711]), .Z(n2700) );
  XOR U2741 ( .A(n2859), .B(n2860), .Z(n2855) );
  AND U2742 ( .A(n2861), .B(n2862), .Z(n2860) );
  XNOR U2743 ( .A(p_input[726]), .B(n2859), .Z(n2862) );
  XNOR U2744 ( .A(n2859), .B(n2709), .Z(n2861) );
  IV U2745 ( .A(p_input[710]), .Z(n2709) );
  XOR U2746 ( .A(n2863), .B(n2864), .Z(n2859) );
  AND U2747 ( .A(n2865), .B(n2866), .Z(n2864) );
  XNOR U2748 ( .A(p_input[725]), .B(n2863), .Z(n2866) );
  XNOR U2749 ( .A(n2863), .B(n2718), .Z(n2865) );
  IV U2750 ( .A(p_input[709]), .Z(n2718) );
  XOR U2751 ( .A(n2867), .B(n2868), .Z(n2863) );
  AND U2752 ( .A(n2869), .B(n2870), .Z(n2868) );
  XNOR U2753 ( .A(p_input[724]), .B(n2867), .Z(n2870) );
  XNOR U2754 ( .A(n2867), .B(n2727), .Z(n2869) );
  IV U2755 ( .A(p_input[708]), .Z(n2727) );
  XOR U2756 ( .A(n2871), .B(n2872), .Z(n2867) );
  AND U2757 ( .A(n2873), .B(n2874), .Z(n2872) );
  XNOR U2758 ( .A(p_input[723]), .B(n2871), .Z(n2874) );
  XNOR U2759 ( .A(n2871), .B(n2736), .Z(n2873) );
  IV U2760 ( .A(p_input[707]), .Z(n2736) );
  XOR U2761 ( .A(n2875), .B(n2876), .Z(n2871) );
  AND U2762 ( .A(n2877), .B(n2878), .Z(n2876) );
  XNOR U2763 ( .A(p_input[722]), .B(n2875), .Z(n2878) );
  XNOR U2764 ( .A(n2875), .B(n2745), .Z(n2877) );
  IV U2765 ( .A(p_input[706]), .Z(n2745) );
  XNOR U2766 ( .A(n2879), .B(n2880), .Z(n2875) );
  AND U2767 ( .A(n2881), .B(n2882), .Z(n2880) );
  XOR U2768 ( .A(p_input[721]), .B(n2879), .Z(n2882) );
  XNOR U2769 ( .A(p_input[705]), .B(n2879), .Z(n2881) );
  AND U2770 ( .A(p_input[720]), .B(n2883), .Z(n2879) );
  IV U2771 ( .A(p_input[704]), .Z(n2883) );
  XOR U2772 ( .A(n2884), .B(n2885), .Z(n2442) );
  AND U2773 ( .A(n168), .B(n2886), .Z(n2885) );
  XNOR U2774 ( .A(n2887), .B(n2884), .Z(n2886) );
  XOR U2775 ( .A(n2888), .B(n2889), .Z(n168) );
  AND U2776 ( .A(n2890), .B(n2891), .Z(n2889) );
  XNOR U2777 ( .A(n2452), .B(n2888), .Z(n2891) );
  AND U2778 ( .A(p_input[703]), .B(p_input[687]), .Z(n2452) );
  XOR U2779 ( .A(n2888), .B(n2453), .Z(n2890) );
  AND U2780 ( .A(p_input[671]), .B(p_input[655]), .Z(n2453) );
  XOR U2781 ( .A(n2892), .B(n2893), .Z(n2888) );
  AND U2782 ( .A(n2894), .B(n2895), .Z(n2893) );
  XOR U2783 ( .A(n2892), .B(n2465), .Z(n2895) );
  XNOR U2784 ( .A(p_input[686]), .B(n2896), .Z(n2465) );
  AND U2785 ( .A(n130), .B(n2897), .Z(n2896) );
  XOR U2786 ( .A(p_input[702]), .B(p_input[686]), .Z(n2897) );
  XNOR U2787 ( .A(n2462), .B(n2892), .Z(n2894) );
  XOR U2788 ( .A(n2898), .B(n2899), .Z(n2462) );
  AND U2789 ( .A(n127), .B(n2900), .Z(n2899) );
  XOR U2790 ( .A(p_input[670]), .B(p_input[654]), .Z(n2900) );
  XOR U2791 ( .A(n2901), .B(n2902), .Z(n2892) );
  AND U2792 ( .A(n2903), .B(n2904), .Z(n2902) );
  XOR U2793 ( .A(n2901), .B(n2477), .Z(n2904) );
  XNOR U2794 ( .A(p_input[685]), .B(n2905), .Z(n2477) );
  AND U2795 ( .A(n130), .B(n2906), .Z(n2905) );
  XOR U2796 ( .A(p_input[701]), .B(p_input[685]), .Z(n2906) );
  XNOR U2797 ( .A(n2474), .B(n2901), .Z(n2903) );
  XOR U2798 ( .A(n2907), .B(n2908), .Z(n2474) );
  AND U2799 ( .A(n127), .B(n2909), .Z(n2908) );
  XOR U2800 ( .A(p_input[669]), .B(p_input[653]), .Z(n2909) );
  XOR U2801 ( .A(n2910), .B(n2911), .Z(n2901) );
  AND U2802 ( .A(n2912), .B(n2913), .Z(n2911) );
  XOR U2803 ( .A(n2910), .B(n2489), .Z(n2913) );
  XNOR U2804 ( .A(p_input[684]), .B(n2914), .Z(n2489) );
  AND U2805 ( .A(n130), .B(n2915), .Z(n2914) );
  XOR U2806 ( .A(p_input[700]), .B(p_input[684]), .Z(n2915) );
  XNOR U2807 ( .A(n2486), .B(n2910), .Z(n2912) );
  XOR U2808 ( .A(n2916), .B(n2917), .Z(n2486) );
  AND U2809 ( .A(n127), .B(n2918), .Z(n2917) );
  XOR U2810 ( .A(p_input[668]), .B(p_input[652]), .Z(n2918) );
  XOR U2811 ( .A(n2919), .B(n2920), .Z(n2910) );
  AND U2812 ( .A(n2921), .B(n2922), .Z(n2920) );
  XOR U2813 ( .A(n2919), .B(n2501), .Z(n2922) );
  XNOR U2814 ( .A(p_input[683]), .B(n2923), .Z(n2501) );
  AND U2815 ( .A(n130), .B(n2924), .Z(n2923) );
  XOR U2816 ( .A(p_input[699]), .B(p_input[683]), .Z(n2924) );
  XNOR U2817 ( .A(n2498), .B(n2919), .Z(n2921) );
  XOR U2818 ( .A(n2925), .B(n2926), .Z(n2498) );
  AND U2819 ( .A(n127), .B(n2927), .Z(n2926) );
  XOR U2820 ( .A(p_input[667]), .B(p_input[651]), .Z(n2927) );
  XOR U2821 ( .A(n2928), .B(n2929), .Z(n2919) );
  AND U2822 ( .A(n2930), .B(n2931), .Z(n2929) );
  XOR U2823 ( .A(n2928), .B(n2513), .Z(n2931) );
  XNOR U2824 ( .A(p_input[682]), .B(n2932), .Z(n2513) );
  AND U2825 ( .A(n130), .B(n2933), .Z(n2932) );
  XOR U2826 ( .A(p_input[698]), .B(p_input[682]), .Z(n2933) );
  XNOR U2827 ( .A(n2510), .B(n2928), .Z(n2930) );
  XOR U2828 ( .A(n2934), .B(n2935), .Z(n2510) );
  AND U2829 ( .A(n127), .B(n2936), .Z(n2935) );
  XOR U2830 ( .A(p_input[666]), .B(p_input[650]), .Z(n2936) );
  XOR U2831 ( .A(n2937), .B(n2938), .Z(n2928) );
  AND U2832 ( .A(n2939), .B(n2940), .Z(n2938) );
  XOR U2833 ( .A(n2937), .B(n2525), .Z(n2940) );
  XNOR U2834 ( .A(p_input[681]), .B(n2941), .Z(n2525) );
  AND U2835 ( .A(n130), .B(n2942), .Z(n2941) );
  XOR U2836 ( .A(p_input[697]), .B(p_input[681]), .Z(n2942) );
  XNOR U2837 ( .A(n2522), .B(n2937), .Z(n2939) );
  XOR U2838 ( .A(n2943), .B(n2944), .Z(n2522) );
  AND U2839 ( .A(n127), .B(n2945), .Z(n2944) );
  XOR U2840 ( .A(p_input[665]), .B(p_input[649]), .Z(n2945) );
  XOR U2841 ( .A(n2946), .B(n2947), .Z(n2937) );
  AND U2842 ( .A(n2948), .B(n2949), .Z(n2947) );
  XOR U2843 ( .A(n2946), .B(n2537), .Z(n2949) );
  XNOR U2844 ( .A(p_input[680]), .B(n2950), .Z(n2537) );
  AND U2845 ( .A(n130), .B(n2951), .Z(n2950) );
  XOR U2846 ( .A(p_input[696]), .B(p_input[680]), .Z(n2951) );
  XNOR U2847 ( .A(n2534), .B(n2946), .Z(n2948) );
  XOR U2848 ( .A(n2952), .B(n2953), .Z(n2534) );
  AND U2849 ( .A(n127), .B(n2954), .Z(n2953) );
  XOR U2850 ( .A(p_input[664]), .B(p_input[648]), .Z(n2954) );
  XOR U2851 ( .A(n2955), .B(n2956), .Z(n2946) );
  AND U2852 ( .A(n2957), .B(n2958), .Z(n2956) );
  XOR U2853 ( .A(n2955), .B(n2549), .Z(n2958) );
  XNOR U2854 ( .A(p_input[679]), .B(n2959), .Z(n2549) );
  AND U2855 ( .A(n130), .B(n2960), .Z(n2959) );
  XOR U2856 ( .A(p_input[695]), .B(p_input[679]), .Z(n2960) );
  XNOR U2857 ( .A(n2546), .B(n2955), .Z(n2957) );
  XOR U2858 ( .A(n2961), .B(n2962), .Z(n2546) );
  AND U2859 ( .A(n127), .B(n2963), .Z(n2962) );
  XOR U2860 ( .A(p_input[663]), .B(p_input[647]), .Z(n2963) );
  XOR U2861 ( .A(n2964), .B(n2965), .Z(n2955) );
  AND U2862 ( .A(n2966), .B(n2967), .Z(n2965) );
  XOR U2863 ( .A(n2964), .B(n2561), .Z(n2967) );
  XNOR U2864 ( .A(p_input[678]), .B(n2968), .Z(n2561) );
  AND U2865 ( .A(n130), .B(n2969), .Z(n2968) );
  XOR U2866 ( .A(p_input[694]), .B(p_input[678]), .Z(n2969) );
  XNOR U2867 ( .A(n2558), .B(n2964), .Z(n2966) );
  XOR U2868 ( .A(n2970), .B(n2971), .Z(n2558) );
  AND U2869 ( .A(n127), .B(n2972), .Z(n2971) );
  XOR U2870 ( .A(p_input[662]), .B(p_input[646]), .Z(n2972) );
  XOR U2871 ( .A(n2973), .B(n2974), .Z(n2964) );
  AND U2872 ( .A(n2975), .B(n2976), .Z(n2974) );
  XOR U2873 ( .A(n2973), .B(n2573), .Z(n2976) );
  XNOR U2874 ( .A(p_input[677]), .B(n2977), .Z(n2573) );
  AND U2875 ( .A(n130), .B(n2978), .Z(n2977) );
  XOR U2876 ( .A(p_input[693]), .B(p_input[677]), .Z(n2978) );
  XNOR U2877 ( .A(n2570), .B(n2973), .Z(n2975) );
  XOR U2878 ( .A(n2979), .B(n2980), .Z(n2570) );
  AND U2879 ( .A(n127), .B(n2981), .Z(n2980) );
  XOR U2880 ( .A(p_input[661]), .B(p_input[645]), .Z(n2981) );
  XOR U2881 ( .A(n2982), .B(n2983), .Z(n2973) );
  AND U2882 ( .A(n2984), .B(n2985), .Z(n2983) );
  XOR U2883 ( .A(n2982), .B(n2585), .Z(n2985) );
  XNOR U2884 ( .A(p_input[676]), .B(n2986), .Z(n2585) );
  AND U2885 ( .A(n130), .B(n2987), .Z(n2986) );
  XOR U2886 ( .A(p_input[692]), .B(p_input[676]), .Z(n2987) );
  XNOR U2887 ( .A(n2582), .B(n2982), .Z(n2984) );
  XOR U2888 ( .A(n2988), .B(n2989), .Z(n2582) );
  AND U2889 ( .A(n127), .B(n2990), .Z(n2989) );
  XOR U2890 ( .A(p_input[660]), .B(p_input[644]), .Z(n2990) );
  XOR U2891 ( .A(n2991), .B(n2992), .Z(n2982) );
  AND U2892 ( .A(n2993), .B(n2994), .Z(n2992) );
  XOR U2893 ( .A(n2597), .B(n2991), .Z(n2994) );
  XNOR U2894 ( .A(p_input[675]), .B(n2995), .Z(n2597) );
  AND U2895 ( .A(n130), .B(n2996), .Z(n2995) );
  XOR U2896 ( .A(p_input[691]), .B(p_input[675]), .Z(n2996) );
  XNOR U2897 ( .A(n2991), .B(n2594), .Z(n2993) );
  XOR U2898 ( .A(n2997), .B(n2998), .Z(n2594) );
  AND U2899 ( .A(n127), .B(n2999), .Z(n2998) );
  XOR U2900 ( .A(p_input[659]), .B(p_input[643]), .Z(n2999) );
  XOR U2901 ( .A(n3000), .B(n3001), .Z(n2991) );
  AND U2902 ( .A(n3002), .B(n3003), .Z(n3001) );
  XOR U2903 ( .A(n3000), .B(n2609), .Z(n3003) );
  XNOR U2904 ( .A(p_input[674]), .B(n3004), .Z(n2609) );
  AND U2905 ( .A(n130), .B(n3005), .Z(n3004) );
  XOR U2906 ( .A(p_input[690]), .B(p_input[674]), .Z(n3005) );
  XNOR U2907 ( .A(n2606), .B(n3000), .Z(n3002) );
  XOR U2908 ( .A(n3006), .B(n3007), .Z(n2606) );
  AND U2909 ( .A(n127), .B(n3008), .Z(n3007) );
  XOR U2910 ( .A(p_input[658]), .B(p_input[642]), .Z(n3008) );
  XOR U2911 ( .A(n3009), .B(n3010), .Z(n3000) );
  AND U2912 ( .A(n3011), .B(n3012), .Z(n3010) );
  XNOR U2913 ( .A(n3013), .B(n2622), .Z(n3012) );
  XNOR U2914 ( .A(p_input[673]), .B(n3014), .Z(n2622) );
  AND U2915 ( .A(n130), .B(n3015), .Z(n3014) );
  XNOR U2916 ( .A(p_input[689]), .B(n3016), .Z(n3015) );
  IV U2917 ( .A(p_input[673]), .Z(n3016) );
  XNOR U2918 ( .A(n2619), .B(n3009), .Z(n3011) );
  XNOR U2919 ( .A(p_input[641]), .B(n3017), .Z(n2619) );
  AND U2920 ( .A(n127), .B(n3018), .Z(n3017) );
  XOR U2921 ( .A(p_input[657]), .B(p_input[641]), .Z(n3018) );
  IV U2922 ( .A(n3013), .Z(n3009) );
  AND U2923 ( .A(n2884), .B(n2887), .Z(n3013) );
  XOR U2924 ( .A(p_input[672]), .B(n3019), .Z(n2887) );
  AND U2925 ( .A(n130), .B(n3020), .Z(n3019) );
  XOR U2926 ( .A(p_input[688]), .B(p_input[672]), .Z(n3020) );
  XOR U2927 ( .A(n3021), .B(n3022), .Z(n130) );
  AND U2928 ( .A(n3023), .B(n3024), .Z(n3022) );
  XNOR U2929 ( .A(p_input[703]), .B(n3021), .Z(n3024) );
  XOR U2930 ( .A(n3021), .B(p_input[687]), .Z(n3023) );
  XOR U2931 ( .A(n3025), .B(n3026), .Z(n3021) );
  AND U2932 ( .A(n3027), .B(n3028), .Z(n3026) );
  XNOR U2933 ( .A(p_input[702]), .B(n3025), .Z(n3028) );
  XOR U2934 ( .A(n3025), .B(p_input[686]), .Z(n3027) );
  XOR U2935 ( .A(n3029), .B(n3030), .Z(n3025) );
  AND U2936 ( .A(n3031), .B(n3032), .Z(n3030) );
  XNOR U2937 ( .A(p_input[701]), .B(n3029), .Z(n3032) );
  XOR U2938 ( .A(n3029), .B(p_input[685]), .Z(n3031) );
  XOR U2939 ( .A(n3033), .B(n3034), .Z(n3029) );
  AND U2940 ( .A(n3035), .B(n3036), .Z(n3034) );
  XNOR U2941 ( .A(p_input[700]), .B(n3033), .Z(n3036) );
  XOR U2942 ( .A(n3033), .B(p_input[684]), .Z(n3035) );
  XOR U2943 ( .A(n3037), .B(n3038), .Z(n3033) );
  AND U2944 ( .A(n3039), .B(n3040), .Z(n3038) );
  XNOR U2945 ( .A(p_input[699]), .B(n3037), .Z(n3040) );
  XOR U2946 ( .A(n3037), .B(p_input[683]), .Z(n3039) );
  XOR U2947 ( .A(n3041), .B(n3042), .Z(n3037) );
  AND U2948 ( .A(n3043), .B(n3044), .Z(n3042) );
  XNOR U2949 ( .A(p_input[698]), .B(n3041), .Z(n3044) );
  XOR U2950 ( .A(n3041), .B(p_input[682]), .Z(n3043) );
  XOR U2951 ( .A(n3045), .B(n3046), .Z(n3041) );
  AND U2952 ( .A(n3047), .B(n3048), .Z(n3046) );
  XNOR U2953 ( .A(p_input[697]), .B(n3045), .Z(n3048) );
  XOR U2954 ( .A(n3045), .B(p_input[681]), .Z(n3047) );
  XOR U2955 ( .A(n3049), .B(n3050), .Z(n3045) );
  AND U2956 ( .A(n3051), .B(n3052), .Z(n3050) );
  XNOR U2957 ( .A(p_input[696]), .B(n3049), .Z(n3052) );
  XOR U2958 ( .A(n3049), .B(p_input[680]), .Z(n3051) );
  XOR U2959 ( .A(n3053), .B(n3054), .Z(n3049) );
  AND U2960 ( .A(n3055), .B(n3056), .Z(n3054) );
  XNOR U2961 ( .A(p_input[695]), .B(n3053), .Z(n3056) );
  XOR U2962 ( .A(n3053), .B(p_input[679]), .Z(n3055) );
  XOR U2963 ( .A(n3057), .B(n3058), .Z(n3053) );
  AND U2964 ( .A(n3059), .B(n3060), .Z(n3058) );
  XNOR U2965 ( .A(p_input[694]), .B(n3057), .Z(n3060) );
  XOR U2966 ( .A(n3057), .B(p_input[678]), .Z(n3059) );
  XOR U2967 ( .A(n3061), .B(n3062), .Z(n3057) );
  AND U2968 ( .A(n3063), .B(n3064), .Z(n3062) );
  XNOR U2969 ( .A(p_input[693]), .B(n3061), .Z(n3064) );
  XOR U2970 ( .A(n3061), .B(p_input[677]), .Z(n3063) );
  XOR U2971 ( .A(n3065), .B(n3066), .Z(n3061) );
  AND U2972 ( .A(n3067), .B(n3068), .Z(n3066) );
  XNOR U2973 ( .A(p_input[692]), .B(n3065), .Z(n3068) );
  XOR U2974 ( .A(n3065), .B(p_input[676]), .Z(n3067) );
  XOR U2975 ( .A(n3069), .B(n3070), .Z(n3065) );
  AND U2976 ( .A(n3071), .B(n3072), .Z(n3070) );
  XNOR U2977 ( .A(p_input[691]), .B(n3069), .Z(n3072) );
  XOR U2978 ( .A(n3069), .B(p_input[675]), .Z(n3071) );
  XOR U2979 ( .A(n3073), .B(n3074), .Z(n3069) );
  AND U2980 ( .A(n3075), .B(n3076), .Z(n3074) );
  XNOR U2981 ( .A(p_input[690]), .B(n3073), .Z(n3076) );
  XOR U2982 ( .A(n3073), .B(p_input[674]), .Z(n3075) );
  XNOR U2983 ( .A(n3077), .B(n3078), .Z(n3073) );
  AND U2984 ( .A(n3079), .B(n3080), .Z(n3078) );
  XOR U2985 ( .A(p_input[689]), .B(n3077), .Z(n3080) );
  XNOR U2986 ( .A(p_input[673]), .B(n3077), .Z(n3079) );
  AND U2987 ( .A(p_input[688]), .B(n3081), .Z(n3077) );
  IV U2988 ( .A(p_input[672]), .Z(n3081) );
  XNOR U2989 ( .A(p_input[640]), .B(n3082), .Z(n2884) );
  AND U2990 ( .A(n127), .B(n3083), .Z(n3082) );
  XOR U2991 ( .A(p_input[656]), .B(p_input[640]), .Z(n3083) );
  XOR U2992 ( .A(n3084), .B(n3085), .Z(n127) );
  AND U2993 ( .A(n3086), .B(n3087), .Z(n3085) );
  XNOR U2994 ( .A(p_input[671]), .B(n3084), .Z(n3087) );
  XOR U2995 ( .A(n3084), .B(p_input[655]), .Z(n3086) );
  XOR U2996 ( .A(n3088), .B(n3089), .Z(n3084) );
  AND U2997 ( .A(n3090), .B(n3091), .Z(n3089) );
  XNOR U2998 ( .A(p_input[670]), .B(n3088), .Z(n3091) );
  XNOR U2999 ( .A(n3088), .B(n2898), .Z(n3090) );
  IV U3000 ( .A(p_input[654]), .Z(n2898) );
  XOR U3001 ( .A(n3092), .B(n3093), .Z(n3088) );
  AND U3002 ( .A(n3094), .B(n3095), .Z(n3093) );
  XNOR U3003 ( .A(p_input[669]), .B(n3092), .Z(n3095) );
  XNOR U3004 ( .A(n3092), .B(n2907), .Z(n3094) );
  IV U3005 ( .A(p_input[653]), .Z(n2907) );
  XOR U3006 ( .A(n3096), .B(n3097), .Z(n3092) );
  AND U3007 ( .A(n3098), .B(n3099), .Z(n3097) );
  XNOR U3008 ( .A(p_input[668]), .B(n3096), .Z(n3099) );
  XNOR U3009 ( .A(n3096), .B(n2916), .Z(n3098) );
  IV U3010 ( .A(p_input[652]), .Z(n2916) );
  XOR U3011 ( .A(n3100), .B(n3101), .Z(n3096) );
  AND U3012 ( .A(n3102), .B(n3103), .Z(n3101) );
  XNOR U3013 ( .A(p_input[667]), .B(n3100), .Z(n3103) );
  XNOR U3014 ( .A(n3100), .B(n2925), .Z(n3102) );
  IV U3015 ( .A(p_input[651]), .Z(n2925) );
  XOR U3016 ( .A(n3104), .B(n3105), .Z(n3100) );
  AND U3017 ( .A(n3106), .B(n3107), .Z(n3105) );
  XNOR U3018 ( .A(p_input[666]), .B(n3104), .Z(n3107) );
  XNOR U3019 ( .A(n3104), .B(n2934), .Z(n3106) );
  IV U3020 ( .A(p_input[650]), .Z(n2934) );
  XOR U3021 ( .A(n3108), .B(n3109), .Z(n3104) );
  AND U3022 ( .A(n3110), .B(n3111), .Z(n3109) );
  XNOR U3023 ( .A(p_input[665]), .B(n3108), .Z(n3111) );
  XNOR U3024 ( .A(n3108), .B(n2943), .Z(n3110) );
  IV U3025 ( .A(p_input[649]), .Z(n2943) );
  XOR U3026 ( .A(n3112), .B(n3113), .Z(n3108) );
  AND U3027 ( .A(n3114), .B(n3115), .Z(n3113) );
  XNOR U3028 ( .A(p_input[664]), .B(n3112), .Z(n3115) );
  XNOR U3029 ( .A(n3112), .B(n2952), .Z(n3114) );
  IV U3030 ( .A(p_input[648]), .Z(n2952) );
  XOR U3031 ( .A(n3116), .B(n3117), .Z(n3112) );
  AND U3032 ( .A(n3118), .B(n3119), .Z(n3117) );
  XNOR U3033 ( .A(p_input[663]), .B(n3116), .Z(n3119) );
  XNOR U3034 ( .A(n3116), .B(n2961), .Z(n3118) );
  IV U3035 ( .A(p_input[647]), .Z(n2961) );
  XOR U3036 ( .A(n3120), .B(n3121), .Z(n3116) );
  AND U3037 ( .A(n3122), .B(n3123), .Z(n3121) );
  XNOR U3038 ( .A(p_input[662]), .B(n3120), .Z(n3123) );
  XNOR U3039 ( .A(n3120), .B(n2970), .Z(n3122) );
  IV U3040 ( .A(p_input[646]), .Z(n2970) );
  XOR U3041 ( .A(n3124), .B(n3125), .Z(n3120) );
  AND U3042 ( .A(n3126), .B(n3127), .Z(n3125) );
  XNOR U3043 ( .A(p_input[661]), .B(n3124), .Z(n3127) );
  XNOR U3044 ( .A(n3124), .B(n2979), .Z(n3126) );
  IV U3045 ( .A(p_input[645]), .Z(n2979) );
  XOR U3046 ( .A(n3128), .B(n3129), .Z(n3124) );
  AND U3047 ( .A(n3130), .B(n3131), .Z(n3129) );
  XNOR U3048 ( .A(p_input[660]), .B(n3128), .Z(n3131) );
  XNOR U3049 ( .A(n3128), .B(n2988), .Z(n3130) );
  IV U3050 ( .A(p_input[644]), .Z(n2988) );
  XOR U3051 ( .A(n3132), .B(n3133), .Z(n3128) );
  AND U3052 ( .A(n3134), .B(n3135), .Z(n3133) );
  XNOR U3053 ( .A(p_input[659]), .B(n3132), .Z(n3135) );
  XNOR U3054 ( .A(n3132), .B(n2997), .Z(n3134) );
  IV U3055 ( .A(p_input[643]), .Z(n2997) );
  XOR U3056 ( .A(n3136), .B(n3137), .Z(n3132) );
  AND U3057 ( .A(n3138), .B(n3139), .Z(n3137) );
  XNOR U3058 ( .A(p_input[658]), .B(n3136), .Z(n3139) );
  XNOR U3059 ( .A(n3136), .B(n3006), .Z(n3138) );
  IV U3060 ( .A(p_input[642]), .Z(n3006) );
  XNOR U3061 ( .A(n3140), .B(n3141), .Z(n3136) );
  AND U3062 ( .A(n3142), .B(n3143), .Z(n3141) );
  XOR U3063 ( .A(p_input[657]), .B(n3140), .Z(n3143) );
  XNOR U3064 ( .A(p_input[641]), .B(n3140), .Z(n3142) );
  AND U3065 ( .A(p_input[656]), .B(n3144), .Z(n3140) );
  IV U3066 ( .A(p_input[640]), .Z(n3144) );
  XOR U3067 ( .A(n3145), .B(n3146), .Z(n2260) );
  AND U3068 ( .A(n247), .B(n3147), .Z(n3146) );
  XNOR U3069 ( .A(n3148), .B(n3145), .Z(n3147) );
  XOR U3070 ( .A(n3149), .B(n3150), .Z(n247) );
  AND U3071 ( .A(n3151), .B(n3152), .Z(n3150) );
  XNOR U3072 ( .A(n2272), .B(n3149), .Z(n3152) );
  AND U3073 ( .A(n3153), .B(n3154), .Z(n2272) );
  XOR U3074 ( .A(n3149), .B(n2271), .Z(n3151) );
  AND U3075 ( .A(n3155), .B(n3156), .Z(n2271) );
  XOR U3076 ( .A(n3157), .B(n3158), .Z(n3149) );
  AND U3077 ( .A(n3159), .B(n3160), .Z(n3158) );
  XOR U3078 ( .A(n3157), .B(n2284), .Z(n3160) );
  XOR U3079 ( .A(n3161), .B(n3162), .Z(n2284) );
  AND U3080 ( .A(n174), .B(n3163), .Z(n3162) );
  XOR U3081 ( .A(n3164), .B(n3161), .Z(n3163) );
  XNOR U3082 ( .A(n2281), .B(n3157), .Z(n3159) );
  XOR U3083 ( .A(n3165), .B(n3166), .Z(n2281) );
  AND U3084 ( .A(n171), .B(n3167), .Z(n3166) );
  XOR U3085 ( .A(n3168), .B(n3165), .Z(n3167) );
  XOR U3086 ( .A(n3169), .B(n3170), .Z(n3157) );
  AND U3087 ( .A(n3171), .B(n3172), .Z(n3170) );
  XOR U3088 ( .A(n3169), .B(n2296), .Z(n3172) );
  XOR U3089 ( .A(n3173), .B(n3174), .Z(n2296) );
  AND U3090 ( .A(n174), .B(n3175), .Z(n3174) );
  XOR U3091 ( .A(n3176), .B(n3173), .Z(n3175) );
  XNOR U3092 ( .A(n2293), .B(n3169), .Z(n3171) );
  XOR U3093 ( .A(n3177), .B(n3178), .Z(n2293) );
  AND U3094 ( .A(n171), .B(n3179), .Z(n3178) );
  XOR U3095 ( .A(n3180), .B(n3177), .Z(n3179) );
  XOR U3096 ( .A(n3181), .B(n3182), .Z(n3169) );
  AND U3097 ( .A(n3183), .B(n3184), .Z(n3182) );
  XOR U3098 ( .A(n3181), .B(n2308), .Z(n3184) );
  XOR U3099 ( .A(n3185), .B(n3186), .Z(n2308) );
  AND U3100 ( .A(n174), .B(n3187), .Z(n3186) );
  XOR U3101 ( .A(n3188), .B(n3185), .Z(n3187) );
  XNOR U3102 ( .A(n2305), .B(n3181), .Z(n3183) );
  XOR U3103 ( .A(n3189), .B(n3190), .Z(n2305) );
  AND U3104 ( .A(n171), .B(n3191), .Z(n3190) );
  XOR U3105 ( .A(n3192), .B(n3189), .Z(n3191) );
  XOR U3106 ( .A(n3193), .B(n3194), .Z(n3181) );
  AND U3107 ( .A(n3195), .B(n3196), .Z(n3194) );
  XOR U3108 ( .A(n3193), .B(n2320), .Z(n3196) );
  XOR U3109 ( .A(n3197), .B(n3198), .Z(n2320) );
  AND U3110 ( .A(n174), .B(n3199), .Z(n3198) );
  XOR U3111 ( .A(n3200), .B(n3197), .Z(n3199) );
  XNOR U3112 ( .A(n2317), .B(n3193), .Z(n3195) );
  XOR U3113 ( .A(n3201), .B(n3202), .Z(n2317) );
  AND U3114 ( .A(n171), .B(n3203), .Z(n3202) );
  XOR U3115 ( .A(n3204), .B(n3201), .Z(n3203) );
  XOR U3116 ( .A(n3205), .B(n3206), .Z(n3193) );
  AND U3117 ( .A(n3207), .B(n3208), .Z(n3206) );
  XOR U3118 ( .A(n3205), .B(n2332), .Z(n3208) );
  XOR U3119 ( .A(n3209), .B(n3210), .Z(n2332) );
  AND U3120 ( .A(n174), .B(n3211), .Z(n3210) );
  XOR U3121 ( .A(n3212), .B(n3209), .Z(n3211) );
  XNOR U3122 ( .A(n2329), .B(n3205), .Z(n3207) );
  XOR U3123 ( .A(n3213), .B(n3214), .Z(n2329) );
  AND U3124 ( .A(n171), .B(n3215), .Z(n3214) );
  XOR U3125 ( .A(n3216), .B(n3213), .Z(n3215) );
  XOR U3126 ( .A(n3217), .B(n3218), .Z(n3205) );
  AND U3127 ( .A(n3219), .B(n3220), .Z(n3218) );
  XOR U3128 ( .A(n3217), .B(n2344), .Z(n3220) );
  XOR U3129 ( .A(n3221), .B(n3222), .Z(n2344) );
  AND U3130 ( .A(n174), .B(n3223), .Z(n3222) );
  XOR U3131 ( .A(n3224), .B(n3221), .Z(n3223) );
  XNOR U3132 ( .A(n2341), .B(n3217), .Z(n3219) );
  XOR U3133 ( .A(n3225), .B(n3226), .Z(n2341) );
  AND U3134 ( .A(n171), .B(n3227), .Z(n3226) );
  XOR U3135 ( .A(n3228), .B(n3225), .Z(n3227) );
  XOR U3136 ( .A(n3229), .B(n3230), .Z(n3217) );
  AND U3137 ( .A(n3231), .B(n3232), .Z(n3230) );
  XOR U3138 ( .A(n3229), .B(n2356), .Z(n3232) );
  XOR U3139 ( .A(n3233), .B(n3234), .Z(n2356) );
  AND U3140 ( .A(n174), .B(n3235), .Z(n3234) );
  XOR U3141 ( .A(n3236), .B(n3233), .Z(n3235) );
  XNOR U3142 ( .A(n2353), .B(n3229), .Z(n3231) );
  XOR U3143 ( .A(n3237), .B(n3238), .Z(n2353) );
  AND U3144 ( .A(n171), .B(n3239), .Z(n3238) );
  XOR U3145 ( .A(n3240), .B(n3237), .Z(n3239) );
  XOR U3146 ( .A(n3241), .B(n3242), .Z(n3229) );
  AND U3147 ( .A(n3243), .B(n3244), .Z(n3242) );
  XOR U3148 ( .A(n3241), .B(n2368), .Z(n3244) );
  XOR U3149 ( .A(n3245), .B(n3246), .Z(n2368) );
  AND U3150 ( .A(n174), .B(n3247), .Z(n3246) );
  XOR U3151 ( .A(n3248), .B(n3245), .Z(n3247) );
  XNOR U3152 ( .A(n2365), .B(n3241), .Z(n3243) );
  XOR U3153 ( .A(n3249), .B(n3250), .Z(n2365) );
  AND U3154 ( .A(n171), .B(n3251), .Z(n3250) );
  XOR U3155 ( .A(n3252), .B(n3249), .Z(n3251) );
  XOR U3156 ( .A(n3253), .B(n3254), .Z(n3241) );
  AND U3157 ( .A(n3255), .B(n3256), .Z(n3254) );
  XOR U3158 ( .A(n3253), .B(n2380), .Z(n3256) );
  XOR U3159 ( .A(n3257), .B(n3258), .Z(n2380) );
  AND U3160 ( .A(n174), .B(n3259), .Z(n3258) );
  XOR U3161 ( .A(n3260), .B(n3257), .Z(n3259) );
  XNOR U3162 ( .A(n2377), .B(n3253), .Z(n3255) );
  XOR U3163 ( .A(n3261), .B(n3262), .Z(n2377) );
  AND U3164 ( .A(n171), .B(n3263), .Z(n3262) );
  XOR U3165 ( .A(n3264), .B(n3261), .Z(n3263) );
  XOR U3166 ( .A(n3265), .B(n3266), .Z(n3253) );
  AND U3167 ( .A(n3267), .B(n3268), .Z(n3266) );
  XOR U3168 ( .A(n3265), .B(n2392), .Z(n3268) );
  XOR U3169 ( .A(n3269), .B(n3270), .Z(n2392) );
  AND U3170 ( .A(n174), .B(n3271), .Z(n3270) );
  XOR U3171 ( .A(n3272), .B(n3269), .Z(n3271) );
  XNOR U3172 ( .A(n2389), .B(n3265), .Z(n3267) );
  XOR U3173 ( .A(n3273), .B(n3274), .Z(n2389) );
  AND U3174 ( .A(n171), .B(n3275), .Z(n3274) );
  XOR U3175 ( .A(n3276), .B(n3273), .Z(n3275) );
  XOR U3176 ( .A(n3277), .B(n3278), .Z(n3265) );
  AND U3177 ( .A(n3279), .B(n3280), .Z(n3278) );
  XOR U3178 ( .A(n3277), .B(n2404), .Z(n3280) );
  XOR U3179 ( .A(n3281), .B(n3282), .Z(n2404) );
  AND U3180 ( .A(n174), .B(n3283), .Z(n3282) );
  XOR U3181 ( .A(n3284), .B(n3281), .Z(n3283) );
  XNOR U3182 ( .A(n2401), .B(n3277), .Z(n3279) );
  XOR U3183 ( .A(n3285), .B(n3286), .Z(n2401) );
  AND U3184 ( .A(n171), .B(n3287), .Z(n3286) );
  XOR U3185 ( .A(n3288), .B(n3285), .Z(n3287) );
  XOR U3186 ( .A(n3289), .B(n3290), .Z(n3277) );
  AND U3187 ( .A(n3291), .B(n3292), .Z(n3290) );
  XOR U3188 ( .A(n2416), .B(n3289), .Z(n3292) );
  XOR U3189 ( .A(n3293), .B(n3294), .Z(n2416) );
  AND U3190 ( .A(n174), .B(n3295), .Z(n3294) );
  XOR U3191 ( .A(n3293), .B(n3296), .Z(n3295) );
  XNOR U3192 ( .A(n3289), .B(n2413), .Z(n3291) );
  XOR U3193 ( .A(n3297), .B(n3298), .Z(n2413) );
  AND U3194 ( .A(n171), .B(n3299), .Z(n3298) );
  XOR U3195 ( .A(n3297), .B(n3300), .Z(n3299) );
  XOR U3196 ( .A(n3301), .B(n3302), .Z(n3289) );
  AND U3197 ( .A(n3303), .B(n3304), .Z(n3302) );
  XOR U3198 ( .A(n3301), .B(n2428), .Z(n3304) );
  XOR U3199 ( .A(n3305), .B(n3306), .Z(n2428) );
  AND U3200 ( .A(n174), .B(n3307), .Z(n3306) );
  XOR U3201 ( .A(n3308), .B(n3305), .Z(n3307) );
  XNOR U3202 ( .A(n2425), .B(n3301), .Z(n3303) );
  XOR U3203 ( .A(n3309), .B(n3310), .Z(n2425) );
  AND U3204 ( .A(n171), .B(n3311), .Z(n3310) );
  XOR U3205 ( .A(n3312), .B(n3309), .Z(n3311) );
  XOR U3206 ( .A(n3313), .B(n3314), .Z(n3301) );
  AND U3207 ( .A(n3315), .B(n3316), .Z(n3314) );
  XNOR U3208 ( .A(n3317), .B(n2441), .Z(n3316) );
  XOR U3209 ( .A(n3318), .B(n3319), .Z(n2441) );
  AND U3210 ( .A(n174), .B(n3320), .Z(n3319) );
  XOR U3211 ( .A(n3321), .B(n3318), .Z(n3320) );
  XNOR U3212 ( .A(n2438), .B(n3313), .Z(n3315) );
  XOR U3213 ( .A(n3322), .B(n3323), .Z(n2438) );
  AND U3214 ( .A(n171), .B(n3324), .Z(n3323) );
  XOR U3215 ( .A(n3325), .B(n3322), .Z(n3324) );
  IV U3216 ( .A(n3317), .Z(n3313) );
  AND U3217 ( .A(n3145), .B(n3148), .Z(n3317) );
  XNOR U3218 ( .A(n3326), .B(n3327), .Z(n3148) );
  AND U3219 ( .A(n174), .B(n3328), .Z(n3327) );
  XNOR U3220 ( .A(n3329), .B(n3326), .Z(n3328) );
  XOR U3221 ( .A(n3330), .B(n3331), .Z(n174) );
  AND U3222 ( .A(n3332), .B(n3333), .Z(n3331) );
  XNOR U3223 ( .A(n3153), .B(n3330), .Z(n3333) );
  AND U3224 ( .A(p_input[639]), .B(p_input[623]), .Z(n3153) );
  XOR U3225 ( .A(n3330), .B(n3154), .Z(n3332) );
  AND U3226 ( .A(p_input[607]), .B(p_input[591]), .Z(n3154) );
  XOR U3227 ( .A(n3334), .B(n3335), .Z(n3330) );
  AND U3228 ( .A(n3336), .B(n3337), .Z(n3335) );
  XOR U3229 ( .A(n3334), .B(n3164), .Z(n3337) );
  XNOR U3230 ( .A(p_input[622]), .B(n3338), .Z(n3164) );
  AND U3231 ( .A(n138), .B(n3339), .Z(n3338) );
  XOR U3232 ( .A(p_input[638]), .B(p_input[622]), .Z(n3339) );
  XNOR U3233 ( .A(n3161), .B(n3334), .Z(n3336) );
  XOR U3234 ( .A(n3340), .B(n3341), .Z(n3161) );
  AND U3235 ( .A(n136), .B(n3342), .Z(n3341) );
  XOR U3236 ( .A(p_input[606]), .B(p_input[590]), .Z(n3342) );
  XOR U3237 ( .A(n3343), .B(n3344), .Z(n3334) );
  AND U3238 ( .A(n3345), .B(n3346), .Z(n3344) );
  XOR U3239 ( .A(n3343), .B(n3176), .Z(n3346) );
  XNOR U3240 ( .A(p_input[621]), .B(n3347), .Z(n3176) );
  AND U3241 ( .A(n138), .B(n3348), .Z(n3347) );
  XOR U3242 ( .A(p_input[637]), .B(p_input[621]), .Z(n3348) );
  XNOR U3243 ( .A(n3173), .B(n3343), .Z(n3345) );
  XOR U3244 ( .A(n3349), .B(n3350), .Z(n3173) );
  AND U3245 ( .A(n136), .B(n3351), .Z(n3350) );
  XOR U3246 ( .A(p_input[605]), .B(p_input[589]), .Z(n3351) );
  XOR U3247 ( .A(n3352), .B(n3353), .Z(n3343) );
  AND U3248 ( .A(n3354), .B(n3355), .Z(n3353) );
  XOR U3249 ( .A(n3352), .B(n3188), .Z(n3355) );
  XNOR U3250 ( .A(p_input[620]), .B(n3356), .Z(n3188) );
  AND U3251 ( .A(n138), .B(n3357), .Z(n3356) );
  XOR U3252 ( .A(p_input[636]), .B(p_input[620]), .Z(n3357) );
  XNOR U3253 ( .A(n3185), .B(n3352), .Z(n3354) );
  XOR U3254 ( .A(n3358), .B(n3359), .Z(n3185) );
  AND U3255 ( .A(n136), .B(n3360), .Z(n3359) );
  XOR U3256 ( .A(p_input[604]), .B(p_input[588]), .Z(n3360) );
  XOR U3257 ( .A(n3361), .B(n3362), .Z(n3352) );
  AND U3258 ( .A(n3363), .B(n3364), .Z(n3362) );
  XOR U3259 ( .A(n3361), .B(n3200), .Z(n3364) );
  XNOR U3260 ( .A(p_input[619]), .B(n3365), .Z(n3200) );
  AND U3261 ( .A(n138), .B(n3366), .Z(n3365) );
  XOR U3262 ( .A(p_input[635]), .B(p_input[619]), .Z(n3366) );
  XNOR U3263 ( .A(n3197), .B(n3361), .Z(n3363) );
  XOR U3264 ( .A(n3367), .B(n3368), .Z(n3197) );
  AND U3265 ( .A(n136), .B(n3369), .Z(n3368) );
  XOR U3266 ( .A(p_input[603]), .B(p_input[587]), .Z(n3369) );
  XOR U3267 ( .A(n3370), .B(n3371), .Z(n3361) );
  AND U3268 ( .A(n3372), .B(n3373), .Z(n3371) );
  XOR U3269 ( .A(n3370), .B(n3212), .Z(n3373) );
  XNOR U3270 ( .A(p_input[618]), .B(n3374), .Z(n3212) );
  AND U3271 ( .A(n138), .B(n3375), .Z(n3374) );
  XOR U3272 ( .A(p_input[634]), .B(p_input[618]), .Z(n3375) );
  XNOR U3273 ( .A(n3209), .B(n3370), .Z(n3372) );
  XOR U3274 ( .A(n3376), .B(n3377), .Z(n3209) );
  AND U3275 ( .A(n136), .B(n3378), .Z(n3377) );
  XOR U3276 ( .A(p_input[602]), .B(p_input[586]), .Z(n3378) );
  XOR U3277 ( .A(n3379), .B(n3380), .Z(n3370) );
  AND U3278 ( .A(n3381), .B(n3382), .Z(n3380) );
  XOR U3279 ( .A(n3379), .B(n3224), .Z(n3382) );
  XNOR U3280 ( .A(p_input[617]), .B(n3383), .Z(n3224) );
  AND U3281 ( .A(n138), .B(n3384), .Z(n3383) );
  XOR U3282 ( .A(p_input[633]), .B(p_input[617]), .Z(n3384) );
  XNOR U3283 ( .A(n3221), .B(n3379), .Z(n3381) );
  XOR U3284 ( .A(n3385), .B(n3386), .Z(n3221) );
  AND U3285 ( .A(n136), .B(n3387), .Z(n3386) );
  XOR U3286 ( .A(p_input[601]), .B(p_input[585]), .Z(n3387) );
  XOR U3287 ( .A(n3388), .B(n3389), .Z(n3379) );
  AND U3288 ( .A(n3390), .B(n3391), .Z(n3389) );
  XOR U3289 ( .A(n3388), .B(n3236), .Z(n3391) );
  XNOR U3290 ( .A(p_input[616]), .B(n3392), .Z(n3236) );
  AND U3291 ( .A(n138), .B(n3393), .Z(n3392) );
  XOR U3292 ( .A(p_input[632]), .B(p_input[616]), .Z(n3393) );
  XNOR U3293 ( .A(n3233), .B(n3388), .Z(n3390) );
  XOR U3294 ( .A(n3394), .B(n3395), .Z(n3233) );
  AND U3295 ( .A(n136), .B(n3396), .Z(n3395) );
  XOR U3296 ( .A(p_input[600]), .B(p_input[584]), .Z(n3396) );
  XOR U3297 ( .A(n3397), .B(n3398), .Z(n3388) );
  AND U3298 ( .A(n3399), .B(n3400), .Z(n3398) );
  XOR U3299 ( .A(n3397), .B(n3248), .Z(n3400) );
  XNOR U3300 ( .A(p_input[615]), .B(n3401), .Z(n3248) );
  AND U3301 ( .A(n138), .B(n3402), .Z(n3401) );
  XOR U3302 ( .A(p_input[631]), .B(p_input[615]), .Z(n3402) );
  XNOR U3303 ( .A(n3245), .B(n3397), .Z(n3399) );
  XOR U3304 ( .A(n3403), .B(n3404), .Z(n3245) );
  AND U3305 ( .A(n136), .B(n3405), .Z(n3404) );
  XOR U3306 ( .A(p_input[599]), .B(p_input[583]), .Z(n3405) );
  XOR U3307 ( .A(n3406), .B(n3407), .Z(n3397) );
  AND U3308 ( .A(n3408), .B(n3409), .Z(n3407) );
  XOR U3309 ( .A(n3406), .B(n3260), .Z(n3409) );
  XNOR U3310 ( .A(p_input[614]), .B(n3410), .Z(n3260) );
  AND U3311 ( .A(n138), .B(n3411), .Z(n3410) );
  XOR U3312 ( .A(p_input[630]), .B(p_input[614]), .Z(n3411) );
  XNOR U3313 ( .A(n3257), .B(n3406), .Z(n3408) );
  XOR U3314 ( .A(n3412), .B(n3413), .Z(n3257) );
  AND U3315 ( .A(n136), .B(n3414), .Z(n3413) );
  XOR U3316 ( .A(p_input[598]), .B(p_input[582]), .Z(n3414) );
  XOR U3317 ( .A(n3415), .B(n3416), .Z(n3406) );
  AND U3318 ( .A(n3417), .B(n3418), .Z(n3416) );
  XOR U3319 ( .A(n3415), .B(n3272), .Z(n3418) );
  XNOR U3320 ( .A(p_input[613]), .B(n3419), .Z(n3272) );
  AND U3321 ( .A(n138), .B(n3420), .Z(n3419) );
  XOR U3322 ( .A(p_input[629]), .B(p_input[613]), .Z(n3420) );
  XNOR U3323 ( .A(n3269), .B(n3415), .Z(n3417) );
  XOR U3324 ( .A(n3421), .B(n3422), .Z(n3269) );
  AND U3325 ( .A(n136), .B(n3423), .Z(n3422) );
  XOR U3326 ( .A(p_input[597]), .B(p_input[581]), .Z(n3423) );
  XOR U3327 ( .A(n3424), .B(n3425), .Z(n3415) );
  AND U3328 ( .A(n3426), .B(n3427), .Z(n3425) );
  XOR U3329 ( .A(n3424), .B(n3284), .Z(n3427) );
  XNOR U3330 ( .A(p_input[612]), .B(n3428), .Z(n3284) );
  AND U3331 ( .A(n138), .B(n3429), .Z(n3428) );
  XOR U3332 ( .A(p_input[628]), .B(p_input[612]), .Z(n3429) );
  XNOR U3333 ( .A(n3281), .B(n3424), .Z(n3426) );
  XOR U3334 ( .A(n3430), .B(n3431), .Z(n3281) );
  AND U3335 ( .A(n136), .B(n3432), .Z(n3431) );
  XOR U3336 ( .A(p_input[596]), .B(p_input[580]), .Z(n3432) );
  XOR U3337 ( .A(n3433), .B(n3434), .Z(n3424) );
  AND U3338 ( .A(n3435), .B(n3436), .Z(n3434) );
  XOR U3339 ( .A(n3296), .B(n3433), .Z(n3436) );
  XNOR U3340 ( .A(p_input[611]), .B(n3437), .Z(n3296) );
  AND U3341 ( .A(n138), .B(n3438), .Z(n3437) );
  XOR U3342 ( .A(p_input[627]), .B(p_input[611]), .Z(n3438) );
  XNOR U3343 ( .A(n3433), .B(n3293), .Z(n3435) );
  XOR U3344 ( .A(n3439), .B(n3440), .Z(n3293) );
  AND U3345 ( .A(n136), .B(n3441), .Z(n3440) );
  XOR U3346 ( .A(p_input[595]), .B(p_input[579]), .Z(n3441) );
  XOR U3347 ( .A(n3442), .B(n3443), .Z(n3433) );
  AND U3348 ( .A(n3444), .B(n3445), .Z(n3443) );
  XOR U3349 ( .A(n3442), .B(n3308), .Z(n3445) );
  XNOR U3350 ( .A(p_input[610]), .B(n3446), .Z(n3308) );
  AND U3351 ( .A(n138), .B(n3447), .Z(n3446) );
  XOR U3352 ( .A(p_input[626]), .B(p_input[610]), .Z(n3447) );
  XNOR U3353 ( .A(n3305), .B(n3442), .Z(n3444) );
  XOR U3354 ( .A(n3448), .B(n3449), .Z(n3305) );
  AND U3355 ( .A(n136), .B(n3450), .Z(n3449) );
  XOR U3356 ( .A(p_input[594]), .B(p_input[578]), .Z(n3450) );
  XOR U3357 ( .A(n3451), .B(n3452), .Z(n3442) );
  AND U3358 ( .A(n3453), .B(n3454), .Z(n3452) );
  XNOR U3359 ( .A(n3455), .B(n3321), .Z(n3454) );
  XNOR U3360 ( .A(p_input[609]), .B(n3456), .Z(n3321) );
  AND U3361 ( .A(n138), .B(n3457), .Z(n3456) );
  XNOR U3362 ( .A(p_input[625]), .B(n3458), .Z(n3457) );
  IV U3363 ( .A(p_input[609]), .Z(n3458) );
  XNOR U3364 ( .A(n3318), .B(n3451), .Z(n3453) );
  XNOR U3365 ( .A(p_input[577]), .B(n3459), .Z(n3318) );
  AND U3366 ( .A(n136), .B(n3460), .Z(n3459) );
  XOR U3367 ( .A(p_input[593]), .B(p_input[577]), .Z(n3460) );
  IV U3368 ( .A(n3455), .Z(n3451) );
  AND U3369 ( .A(n3326), .B(n3329), .Z(n3455) );
  XOR U3370 ( .A(p_input[608]), .B(n3461), .Z(n3329) );
  AND U3371 ( .A(n138), .B(n3462), .Z(n3461) );
  XOR U3372 ( .A(p_input[624]), .B(p_input[608]), .Z(n3462) );
  XOR U3373 ( .A(n3463), .B(n3464), .Z(n138) );
  AND U3374 ( .A(n3465), .B(n3466), .Z(n3464) );
  XNOR U3375 ( .A(p_input[639]), .B(n3463), .Z(n3466) );
  XOR U3376 ( .A(n3463), .B(p_input[623]), .Z(n3465) );
  XOR U3377 ( .A(n3467), .B(n3468), .Z(n3463) );
  AND U3378 ( .A(n3469), .B(n3470), .Z(n3468) );
  XNOR U3379 ( .A(p_input[638]), .B(n3467), .Z(n3470) );
  XOR U3380 ( .A(n3467), .B(p_input[622]), .Z(n3469) );
  XOR U3381 ( .A(n3471), .B(n3472), .Z(n3467) );
  AND U3382 ( .A(n3473), .B(n3474), .Z(n3472) );
  XNOR U3383 ( .A(p_input[637]), .B(n3471), .Z(n3474) );
  XOR U3384 ( .A(n3471), .B(p_input[621]), .Z(n3473) );
  XOR U3385 ( .A(n3475), .B(n3476), .Z(n3471) );
  AND U3386 ( .A(n3477), .B(n3478), .Z(n3476) );
  XNOR U3387 ( .A(p_input[636]), .B(n3475), .Z(n3478) );
  XOR U3388 ( .A(n3475), .B(p_input[620]), .Z(n3477) );
  XOR U3389 ( .A(n3479), .B(n3480), .Z(n3475) );
  AND U3390 ( .A(n3481), .B(n3482), .Z(n3480) );
  XNOR U3391 ( .A(p_input[635]), .B(n3479), .Z(n3482) );
  XOR U3392 ( .A(n3479), .B(p_input[619]), .Z(n3481) );
  XOR U3393 ( .A(n3483), .B(n3484), .Z(n3479) );
  AND U3394 ( .A(n3485), .B(n3486), .Z(n3484) );
  XNOR U3395 ( .A(p_input[634]), .B(n3483), .Z(n3486) );
  XOR U3396 ( .A(n3483), .B(p_input[618]), .Z(n3485) );
  XOR U3397 ( .A(n3487), .B(n3488), .Z(n3483) );
  AND U3398 ( .A(n3489), .B(n3490), .Z(n3488) );
  XNOR U3399 ( .A(p_input[633]), .B(n3487), .Z(n3490) );
  XOR U3400 ( .A(n3487), .B(p_input[617]), .Z(n3489) );
  XOR U3401 ( .A(n3491), .B(n3492), .Z(n3487) );
  AND U3402 ( .A(n3493), .B(n3494), .Z(n3492) );
  XNOR U3403 ( .A(p_input[632]), .B(n3491), .Z(n3494) );
  XOR U3404 ( .A(n3491), .B(p_input[616]), .Z(n3493) );
  XOR U3405 ( .A(n3495), .B(n3496), .Z(n3491) );
  AND U3406 ( .A(n3497), .B(n3498), .Z(n3496) );
  XNOR U3407 ( .A(p_input[631]), .B(n3495), .Z(n3498) );
  XOR U3408 ( .A(n3495), .B(p_input[615]), .Z(n3497) );
  XOR U3409 ( .A(n3499), .B(n3500), .Z(n3495) );
  AND U3410 ( .A(n3501), .B(n3502), .Z(n3500) );
  XNOR U3411 ( .A(p_input[630]), .B(n3499), .Z(n3502) );
  XOR U3412 ( .A(n3499), .B(p_input[614]), .Z(n3501) );
  XOR U3413 ( .A(n3503), .B(n3504), .Z(n3499) );
  AND U3414 ( .A(n3505), .B(n3506), .Z(n3504) );
  XNOR U3415 ( .A(p_input[629]), .B(n3503), .Z(n3506) );
  XOR U3416 ( .A(n3503), .B(p_input[613]), .Z(n3505) );
  XOR U3417 ( .A(n3507), .B(n3508), .Z(n3503) );
  AND U3418 ( .A(n3509), .B(n3510), .Z(n3508) );
  XNOR U3419 ( .A(p_input[628]), .B(n3507), .Z(n3510) );
  XOR U3420 ( .A(n3507), .B(p_input[612]), .Z(n3509) );
  XOR U3421 ( .A(n3511), .B(n3512), .Z(n3507) );
  AND U3422 ( .A(n3513), .B(n3514), .Z(n3512) );
  XNOR U3423 ( .A(p_input[627]), .B(n3511), .Z(n3514) );
  XOR U3424 ( .A(n3511), .B(p_input[611]), .Z(n3513) );
  XOR U3425 ( .A(n3515), .B(n3516), .Z(n3511) );
  AND U3426 ( .A(n3517), .B(n3518), .Z(n3516) );
  XNOR U3427 ( .A(p_input[626]), .B(n3515), .Z(n3518) );
  XOR U3428 ( .A(n3515), .B(p_input[610]), .Z(n3517) );
  XNOR U3429 ( .A(n3519), .B(n3520), .Z(n3515) );
  AND U3430 ( .A(n3521), .B(n3522), .Z(n3520) );
  XOR U3431 ( .A(p_input[625]), .B(n3519), .Z(n3522) );
  XNOR U3432 ( .A(p_input[609]), .B(n3519), .Z(n3521) );
  AND U3433 ( .A(p_input[624]), .B(n3523), .Z(n3519) );
  IV U3434 ( .A(p_input[608]), .Z(n3523) );
  XNOR U3435 ( .A(p_input[576]), .B(n3524), .Z(n3326) );
  AND U3436 ( .A(n136), .B(n3525), .Z(n3524) );
  XOR U3437 ( .A(p_input[592]), .B(p_input[576]), .Z(n3525) );
  XOR U3438 ( .A(n3526), .B(n3527), .Z(n136) );
  AND U3439 ( .A(n3528), .B(n3529), .Z(n3527) );
  XNOR U3440 ( .A(p_input[607]), .B(n3526), .Z(n3529) );
  XOR U3441 ( .A(n3526), .B(p_input[591]), .Z(n3528) );
  XOR U3442 ( .A(n3530), .B(n3531), .Z(n3526) );
  AND U3443 ( .A(n3532), .B(n3533), .Z(n3531) );
  XNOR U3444 ( .A(p_input[606]), .B(n3530), .Z(n3533) );
  XNOR U3445 ( .A(n3530), .B(n3340), .Z(n3532) );
  IV U3446 ( .A(p_input[590]), .Z(n3340) );
  XOR U3447 ( .A(n3534), .B(n3535), .Z(n3530) );
  AND U3448 ( .A(n3536), .B(n3537), .Z(n3535) );
  XNOR U3449 ( .A(p_input[605]), .B(n3534), .Z(n3537) );
  XNOR U3450 ( .A(n3534), .B(n3349), .Z(n3536) );
  IV U3451 ( .A(p_input[589]), .Z(n3349) );
  XOR U3452 ( .A(n3538), .B(n3539), .Z(n3534) );
  AND U3453 ( .A(n3540), .B(n3541), .Z(n3539) );
  XNOR U3454 ( .A(p_input[604]), .B(n3538), .Z(n3541) );
  XNOR U3455 ( .A(n3538), .B(n3358), .Z(n3540) );
  IV U3456 ( .A(p_input[588]), .Z(n3358) );
  XOR U3457 ( .A(n3542), .B(n3543), .Z(n3538) );
  AND U3458 ( .A(n3544), .B(n3545), .Z(n3543) );
  XNOR U3459 ( .A(p_input[603]), .B(n3542), .Z(n3545) );
  XNOR U3460 ( .A(n3542), .B(n3367), .Z(n3544) );
  IV U3461 ( .A(p_input[587]), .Z(n3367) );
  XOR U3462 ( .A(n3546), .B(n3547), .Z(n3542) );
  AND U3463 ( .A(n3548), .B(n3549), .Z(n3547) );
  XNOR U3464 ( .A(p_input[602]), .B(n3546), .Z(n3549) );
  XNOR U3465 ( .A(n3546), .B(n3376), .Z(n3548) );
  IV U3466 ( .A(p_input[586]), .Z(n3376) );
  XOR U3467 ( .A(n3550), .B(n3551), .Z(n3546) );
  AND U3468 ( .A(n3552), .B(n3553), .Z(n3551) );
  XNOR U3469 ( .A(p_input[601]), .B(n3550), .Z(n3553) );
  XNOR U3470 ( .A(n3550), .B(n3385), .Z(n3552) );
  IV U3471 ( .A(p_input[585]), .Z(n3385) );
  XOR U3472 ( .A(n3554), .B(n3555), .Z(n3550) );
  AND U3473 ( .A(n3556), .B(n3557), .Z(n3555) );
  XNOR U3474 ( .A(p_input[600]), .B(n3554), .Z(n3557) );
  XNOR U3475 ( .A(n3554), .B(n3394), .Z(n3556) );
  IV U3476 ( .A(p_input[584]), .Z(n3394) );
  XOR U3477 ( .A(n3558), .B(n3559), .Z(n3554) );
  AND U3478 ( .A(n3560), .B(n3561), .Z(n3559) );
  XNOR U3479 ( .A(p_input[599]), .B(n3558), .Z(n3561) );
  XNOR U3480 ( .A(n3558), .B(n3403), .Z(n3560) );
  IV U3481 ( .A(p_input[583]), .Z(n3403) );
  XOR U3482 ( .A(n3562), .B(n3563), .Z(n3558) );
  AND U3483 ( .A(n3564), .B(n3565), .Z(n3563) );
  XNOR U3484 ( .A(p_input[598]), .B(n3562), .Z(n3565) );
  XNOR U3485 ( .A(n3562), .B(n3412), .Z(n3564) );
  IV U3486 ( .A(p_input[582]), .Z(n3412) );
  XOR U3487 ( .A(n3566), .B(n3567), .Z(n3562) );
  AND U3488 ( .A(n3568), .B(n3569), .Z(n3567) );
  XNOR U3489 ( .A(p_input[597]), .B(n3566), .Z(n3569) );
  XNOR U3490 ( .A(n3566), .B(n3421), .Z(n3568) );
  IV U3491 ( .A(p_input[581]), .Z(n3421) );
  XOR U3492 ( .A(n3570), .B(n3571), .Z(n3566) );
  AND U3493 ( .A(n3572), .B(n3573), .Z(n3571) );
  XNOR U3494 ( .A(p_input[596]), .B(n3570), .Z(n3573) );
  XNOR U3495 ( .A(n3570), .B(n3430), .Z(n3572) );
  IV U3496 ( .A(p_input[580]), .Z(n3430) );
  XOR U3497 ( .A(n3574), .B(n3575), .Z(n3570) );
  AND U3498 ( .A(n3576), .B(n3577), .Z(n3575) );
  XNOR U3499 ( .A(p_input[595]), .B(n3574), .Z(n3577) );
  XNOR U3500 ( .A(n3574), .B(n3439), .Z(n3576) );
  IV U3501 ( .A(p_input[579]), .Z(n3439) );
  XOR U3502 ( .A(n3578), .B(n3579), .Z(n3574) );
  AND U3503 ( .A(n3580), .B(n3581), .Z(n3579) );
  XNOR U3504 ( .A(p_input[594]), .B(n3578), .Z(n3581) );
  XNOR U3505 ( .A(n3578), .B(n3448), .Z(n3580) );
  IV U3506 ( .A(p_input[578]), .Z(n3448) );
  XNOR U3507 ( .A(n3582), .B(n3583), .Z(n3578) );
  AND U3508 ( .A(n3584), .B(n3585), .Z(n3583) );
  XOR U3509 ( .A(p_input[593]), .B(n3582), .Z(n3585) );
  XNOR U3510 ( .A(p_input[577]), .B(n3582), .Z(n3584) );
  AND U3511 ( .A(p_input[592]), .B(n3586), .Z(n3582) );
  IV U3512 ( .A(p_input[576]), .Z(n3586) );
  XOR U3513 ( .A(n3587), .B(n3588), .Z(n3145) );
  AND U3514 ( .A(n171), .B(n3589), .Z(n3588) );
  XNOR U3515 ( .A(n3590), .B(n3587), .Z(n3589) );
  XOR U3516 ( .A(n3591), .B(n3592), .Z(n171) );
  AND U3517 ( .A(n3593), .B(n3594), .Z(n3592) );
  XNOR U3518 ( .A(n3156), .B(n3591), .Z(n3594) );
  AND U3519 ( .A(p_input[575]), .B(p_input[559]), .Z(n3156) );
  XOR U3520 ( .A(n3591), .B(n3155), .Z(n3593) );
  AND U3521 ( .A(p_input[527]), .B(p_input[543]), .Z(n3155) );
  XOR U3522 ( .A(n3595), .B(n3596), .Z(n3591) );
  AND U3523 ( .A(n3597), .B(n3598), .Z(n3596) );
  XOR U3524 ( .A(n3595), .B(n3168), .Z(n3598) );
  XNOR U3525 ( .A(p_input[558]), .B(n3599), .Z(n3168) );
  AND U3526 ( .A(n142), .B(n3600), .Z(n3599) );
  XOR U3527 ( .A(p_input[574]), .B(p_input[558]), .Z(n3600) );
  XNOR U3528 ( .A(n3165), .B(n3595), .Z(n3597) );
  XOR U3529 ( .A(n3601), .B(n3602), .Z(n3165) );
  AND U3530 ( .A(n139), .B(n3603), .Z(n3602) );
  XOR U3531 ( .A(p_input[542]), .B(p_input[526]), .Z(n3603) );
  XOR U3532 ( .A(n3604), .B(n3605), .Z(n3595) );
  AND U3533 ( .A(n3606), .B(n3607), .Z(n3605) );
  XOR U3534 ( .A(n3604), .B(n3180), .Z(n3607) );
  XNOR U3535 ( .A(p_input[557]), .B(n3608), .Z(n3180) );
  AND U3536 ( .A(n142), .B(n3609), .Z(n3608) );
  XOR U3537 ( .A(p_input[573]), .B(p_input[557]), .Z(n3609) );
  XNOR U3538 ( .A(n3177), .B(n3604), .Z(n3606) );
  XOR U3539 ( .A(n3610), .B(n3611), .Z(n3177) );
  AND U3540 ( .A(n139), .B(n3612), .Z(n3611) );
  XOR U3541 ( .A(p_input[541]), .B(p_input[525]), .Z(n3612) );
  XOR U3542 ( .A(n3613), .B(n3614), .Z(n3604) );
  AND U3543 ( .A(n3615), .B(n3616), .Z(n3614) );
  XOR U3544 ( .A(n3613), .B(n3192), .Z(n3616) );
  XNOR U3545 ( .A(p_input[556]), .B(n3617), .Z(n3192) );
  AND U3546 ( .A(n142), .B(n3618), .Z(n3617) );
  XOR U3547 ( .A(p_input[572]), .B(p_input[556]), .Z(n3618) );
  XNOR U3548 ( .A(n3189), .B(n3613), .Z(n3615) );
  XOR U3549 ( .A(n3619), .B(n3620), .Z(n3189) );
  AND U3550 ( .A(n139), .B(n3621), .Z(n3620) );
  XOR U3551 ( .A(p_input[540]), .B(p_input[524]), .Z(n3621) );
  XOR U3552 ( .A(n3622), .B(n3623), .Z(n3613) );
  AND U3553 ( .A(n3624), .B(n3625), .Z(n3623) );
  XOR U3554 ( .A(n3622), .B(n3204), .Z(n3625) );
  XNOR U3555 ( .A(p_input[555]), .B(n3626), .Z(n3204) );
  AND U3556 ( .A(n142), .B(n3627), .Z(n3626) );
  XOR U3557 ( .A(p_input[571]), .B(p_input[555]), .Z(n3627) );
  XNOR U3558 ( .A(n3201), .B(n3622), .Z(n3624) );
  XOR U3559 ( .A(n3628), .B(n3629), .Z(n3201) );
  AND U3560 ( .A(n139), .B(n3630), .Z(n3629) );
  XOR U3561 ( .A(p_input[539]), .B(p_input[523]), .Z(n3630) );
  XOR U3562 ( .A(n3631), .B(n3632), .Z(n3622) );
  AND U3563 ( .A(n3633), .B(n3634), .Z(n3632) );
  XOR U3564 ( .A(n3631), .B(n3216), .Z(n3634) );
  XNOR U3565 ( .A(p_input[554]), .B(n3635), .Z(n3216) );
  AND U3566 ( .A(n142), .B(n3636), .Z(n3635) );
  XOR U3567 ( .A(p_input[570]), .B(p_input[554]), .Z(n3636) );
  XNOR U3568 ( .A(n3213), .B(n3631), .Z(n3633) );
  XOR U3569 ( .A(n3637), .B(n3638), .Z(n3213) );
  AND U3570 ( .A(n139), .B(n3639), .Z(n3638) );
  XOR U3571 ( .A(p_input[538]), .B(p_input[522]), .Z(n3639) );
  XOR U3572 ( .A(n3640), .B(n3641), .Z(n3631) );
  AND U3573 ( .A(n3642), .B(n3643), .Z(n3641) );
  XOR U3574 ( .A(n3640), .B(n3228), .Z(n3643) );
  XNOR U3575 ( .A(p_input[553]), .B(n3644), .Z(n3228) );
  AND U3576 ( .A(n142), .B(n3645), .Z(n3644) );
  XOR U3577 ( .A(p_input[569]), .B(p_input[553]), .Z(n3645) );
  XNOR U3578 ( .A(n3225), .B(n3640), .Z(n3642) );
  XOR U3579 ( .A(n3646), .B(n3647), .Z(n3225) );
  AND U3580 ( .A(n139), .B(n3648), .Z(n3647) );
  XOR U3581 ( .A(p_input[537]), .B(p_input[521]), .Z(n3648) );
  XOR U3582 ( .A(n3649), .B(n3650), .Z(n3640) );
  AND U3583 ( .A(n3651), .B(n3652), .Z(n3650) );
  XOR U3584 ( .A(n3649), .B(n3240), .Z(n3652) );
  XNOR U3585 ( .A(p_input[552]), .B(n3653), .Z(n3240) );
  AND U3586 ( .A(n142), .B(n3654), .Z(n3653) );
  XOR U3587 ( .A(p_input[568]), .B(p_input[552]), .Z(n3654) );
  XNOR U3588 ( .A(n3237), .B(n3649), .Z(n3651) );
  XOR U3589 ( .A(n3655), .B(n3656), .Z(n3237) );
  AND U3590 ( .A(n139), .B(n3657), .Z(n3656) );
  XOR U3591 ( .A(p_input[536]), .B(p_input[520]), .Z(n3657) );
  XOR U3592 ( .A(n3658), .B(n3659), .Z(n3649) );
  AND U3593 ( .A(n3660), .B(n3661), .Z(n3659) );
  XOR U3594 ( .A(n3658), .B(n3252), .Z(n3661) );
  XNOR U3595 ( .A(p_input[551]), .B(n3662), .Z(n3252) );
  AND U3596 ( .A(n142), .B(n3663), .Z(n3662) );
  XOR U3597 ( .A(p_input[567]), .B(p_input[551]), .Z(n3663) );
  XNOR U3598 ( .A(n3249), .B(n3658), .Z(n3660) );
  XOR U3599 ( .A(n3664), .B(n3665), .Z(n3249) );
  AND U3600 ( .A(n139), .B(n3666), .Z(n3665) );
  XOR U3601 ( .A(p_input[535]), .B(p_input[519]), .Z(n3666) );
  XOR U3602 ( .A(n3667), .B(n3668), .Z(n3658) );
  AND U3603 ( .A(n3669), .B(n3670), .Z(n3668) );
  XOR U3604 ( .A(n3667), .B(n3264), .Z(n3670) );
  XNOR U3605 ( .A(p_input[550]), .B(n3671), .Z(n3264) );
  AND U3606 ( .A(n142), .B(n3672), .Z(n3671) );
  XOR U3607 ( .A(p_input[566]), .B(p_input[550]), .Z(n3672) );
  XNOR U3608 ( .A(n3261), .B(n3667), .Z(n3669) );
  XOR U3609 ( .A(n3673), .B(n3674), .Z(n3261) );
  AND U3610 ( .A(n139), .B(n3675), .Z(n3674) );
  XOR U3611 ( .A(p_input[534]), .B(p_input[518]), .Z(n3675) );
  XOR U3612 ( .A(n3676), .B(n3677), .Z(n3667) );
  AND U3613 ( .A(n3678), .B(n3679), .Z(n3677) );
  XOR U3614 ( .A(n3676), .B(n3276), .Z(n3679) );
  XNOR U3615 ( .A(p_input[549]), .B(n3680), .Z(n3276) );
  AND U3616 ( .A(n142), .B(n3681), .Z(n3680) );
  XOR U3617 ( .A(p_input[565]), .B(p_input[549]), .Z(n3681) );
  XNOR U3618 ( .A(n3273), .B(n3676), .Z(n3678) );
  XOR U3619 ( .A(n3682), .B(n3683), .Z(n3273) );
  AND U3620 ( .A(n139), .B(n3684), .Z(n3683) );
  XOR U3621 ( .A(p_input[533]), .B(p_input[517]), .Z(n3684) );
  XOR U3622 ( .A(n3685), .B(n3686), .Z(n3676) );
  AND U3623 ( .A(n3687), .B(n3688), .Z(n3686) );
  XOR U3624 ( .A(n3685), .B(n3288), .Z(n3688) );
  XNOR U3625 ( .A(p_input[548]), .B(n3689), .Z(n3288) );
  AND U3626 ( .A(n142), .B(n3690), .Z(n3689) );
  XOR U3627 ( .A(p_input[564]), .B(p_input[548]), .Z(n3690) );
  XNOR U3628 ( .A(n3285), .B(n3685), .Z(n3687) );
  XOR U3629 ( .A(n3691), .B(n3692), .Z(n3285) );
  AND U3630 ( .A(n139), .B(n3693), .Z(n3692) );
  XOR U3631 ( .A(p_input[532]), .B(p_input[516]), .Z(n3693) );
  XOR U3632 ( .A(n3694), .B(n3695), .Z(n3685) );
  AND U3633 ( .A(n3696), .B(n3697), .Z(n3695) );
  XOR U3634 ( .A(n3300), .B(n3694), .Z(n3697) );
  XNOR U3635 ( .A(p_input[547]), .B(n3698), .Z(n3300) );
  AND U3636 ( .A(n142), .B(n3699), .Z(n3698) );
  XOR U3637 ( .A(p_input[563]), .B(p_input[547]), .Z(n3699) );
  XNOR U3638 ( .A(n3694), .B(n3297), .Z(n3696) );
  XOR U3639 ( .A(n3700), .B(n3701), .Z(n3297) );
  AND U3640 ( .A(n139), .B(n3702), .Z(n3701) );
  XOR U3641 ( .A(p_input[531]), .B(p_input[515]), .Z(n3702) );
  XOR U3642 ( .A(n3703), .B(n3704), .Z(n3694) );
  AND U3643 ( .A(n3705), .B(n3706), .Z(n3704) );
  XOR U3644 ( .A(n3703), .B(n3312), .Z(n3706) );
  XNOR U3645 ( .A(p_input[546]), .B(n3707), .Z(n3312) );
  AND U3646 ( .A(n142), .B(n3708), .Z(n3707) );
  XOR U3647 ( .A(p_input[562]), .B(p_input[546]), .Z(n3708) );
  XNOR U3648 ( .A(n3309), .B(n3703), .Z(n3705) );
  XOR U3649 ( .A(n3709), .B(n3710), .Z(n3309) );
  AND U3650 ( .A(n139), .B(n3711), .Z(n3710) );
  XOR U3651 ( .A(p_input[530]), .B(p_input[514]), .Z(n3711) );
  XOR U3652 ( .A(n3712), .B(n3713), .Z(n3703) );
  AND U3653 ( .A(n3714), .B(n3715), .Z(n3713) );
  XNOR U3654 ( .A(n3716), .B(n3325), .Z(n3715) );
  XNOR U3655 ( .A(p_input[545]), .B(n3717), .Z(n3325) );
  AND U3656 ( .A(n142), .B(n3718), .Z(n3717) );
  XNOR U3657 ( .A(p_input[561]), .B(n3719), .Z(n3718) );
  IV U3658 ( .A(p_input[545]), .Z(n3719) );
  XNOR U3659 ( .A(n3322), .B(n3712), .Z(n3714) );
  XNOR U3660 ( .A(p_input[513]), .B(n3720), .Z(n3322) );
  AND U3661 ( .A(n139), .B(n3721), .Z(n3720) );
  XOR U3662 ( .A(p_input[529]), .B(p_input[513]), .Z(n3721) );
  IV U3663 ( .A(n3716), .Z(n3712) );
  AND U3664 ( .A(n3587), .B(n3590), .Z(n3716) );
  XOR U3665 ( .A(p_input[544]), .B(n3722), .Z(n3590) );
  AND U3666 ( .A(n142), .B(n3723), .Z(n3722) );
  XOR U3667 ( .A(p_input[560]), .B(p_input[544]), .Z(n3723) );
  XOR U3668 ( .A(n3724), .B(n3725), .Z(n142) );
  AND U3669 ( .A(n3726), .B(n3727), .Z(n3725) );
  XNOR U3670 ( .A(p_input[575]), .B(n3724), .Z(n3727) );
  XOR U3671 ( .A(n3724), .B(p_input[559]), .Z(n3726) );
  XOR U3672 ( .A(n3728), .B(n3729), .Z(n3724) );
  AND U3673 ( .A(n3730), .B(n3731), .Z(n3729) );
  XNOR U3674 ( .A(p_input[574]), .B(n3728), .Z(n3731) );
  XOR U3675 ( .A(n3728), .B(p_input[558]), .Z(n3730) );
  XOR U3676 ( .A(n3732), .B(n3733), .Z(n3728) );
  AND U3677 ( .A(n3734), .B(n3735), .Z(n3733) );
  XNOR U3678 ( .A(p_input[573]), .B(n3732), .Z(n3735) );
  XOR U3679 ( .A(n3732), .B(p_input[557]), .Z(n3734) );
  XOR U3680 ( .A(n3736), .B(n3737), .Z(n3732) );
  AND U3681 ( .A(n3738), .B(n3739), .Z(n3737) );
  XNOR U3682 ( .A(p_input[572]), .B(n3736), .Z(n3739) );
  XOR U3683 ( .A(n3736), .B(p_input[556]), .Z(n3738) );
  XOR U3684 ( .A(n3740), .B(n3741), .Z(n3736) );
  AND U3685 ( .A(n3742), .B(n3743), .Z(n3741) );
  XNOR U3686 ( .A(p_input[571]), .B(n3740), .Z(n3743) );
  XOR U3687 ( .A(n3740), .B(p_input[555]), .Z(n3742) );
  XOR U3688 ( .A(n3744), .B(n3745), .Z(n3740) );
  AND U3689 ( .A(n3746), .B(n3747), .Z(n3745) );
  XNOR U3690 ( .A(p_input[570]), .B(n3744), .Z(n3747) );
  XOR U3691 ( .A(n3744), .B(p_input[554]), .Z(n3746) );
  XOR U3692 ( .A(n3748), .B(n3749), .Z(n3744) );
  AND U3693 ( .A(n3750), .B(n3751), .Z(n3749) );
  XNOR U3694 ( .A(p_input[569]), .B(n3748), .Z(n3751) );
  XOR U3695 ( .A(n3748), .B(p_input[553]), .Z(n3750) );
  XOR U3696 ( .A(n3752), .B(n3753), .Z(n3748) );
  AND U3697 ( .A(n3754), .B(n3755), .Z(n3753) );
  XNOR U3698 ( .A(p_input[568]), .B(n3752), .Z(n3755) );
  XOR U3699 ( .A(n3752), .B(p_input[552]), .Z(n3754) );
  XOR U3700 ( .A(n3756), .B(n3757), .Z(n3752) );
  AND U3701 ( .A(n3758), .B(n3759), .Z(n3757) );
  XNOR U3702 ( .A(p_input[567]), .B(n3756), .Z(n3759) );
  XOR U3703 ( .A(n3756), .B(p_input[551]), .Z(n3758) );
  XOR U3704 ( .A(n3760), .B(n3761), .Z(n3756) );
  AND U3705 ( .A(n3762), .B(n3763), .Z(n3761) );
  XNOR U3706 ( .A(p_input[566]), .B(n3760), .Z(n3763) );
  XOR U3707 ( .A(n3760), .B(p_input[550]), .Z(n3762) );
  XOR U3708 ( .A(n3764), .B(n3765), .Z(n3760) );
  AND U3709 ( .A(n3766), .B(n3767), .Z(n3765) );
  XNOR U3710 ( .A(p_input[565]), .B(n3764), .Z(n3767) );
  XOR U3711 ( .A(n3764), .B(p_input[549]), .Z(n3766) );
  XOR U3712 ( .A(n3768), .B(n3769), .Z(n3764) );
  AND U3713 ( .A(n3770), .B(n3771), .Z(n3769) );
  XNOR U3714 ( .A(p_input[564]), .B(n3768), .Z(n3771) );
  XOR U3715 ( .A(n3768), .B(p_input[548]), .Z(n3770) );
  XOR U3716 ( .A(n3772), .B(n3773), .Z(n3768) );
  AND U3717 ( .A(n3774), .B(n3775), .Z(n3773) );
  XNOR U3718 ( .A(p_input[563]), .B(n3772), .Z(n3775) );
  XOR U3719 ( .A(n3772), .B(p_input[547]), .Z(n3774) );
  XOR U3720 ( .A(n3776), .B(n3777), .Z(n3772) );
  AND U3721 ( .A(n3778), .B(n3779), .Z(n3777) );
  XNOR U3722 ( .A(p_input[562]), .B(n3776), .Z(n3779) );
  XOR U3723 ( .A(n3776), .B(p_input[546]), .Z(n3778) );
  XNOR U3724 ( .A(n3780), .B(n3781), .Z(n3776) );
  AND U3725 ( .A(n3782), .B(n3783), .Z(n3781) );
  XOR U3726 ( .A(p_input[561]), .B(n3780), .Z(n3783) );
  XNOR U3727 ( .A(p_input[545]), .B(n3780), .Z(n3782) );
  AND U3728 ( .A(p_input[560]), .B(n3784), .Z(n3780) );
  IV U3729 ( .A(p_input[544]), .Z(n3784) );
  XNOR U3730 ( .A(p_input[512]), .B(n3785), .Z(n3587) );
  AND U3731 ( .A(n139), .B(n3786), .Z(n3785) );
  XOR U3732 ( .A(p_input[528]), .B(p_input[512]), .Z(n3786) );
  XOR U3733 ( .A(n3787), .B(n3788), .Z(n139) );
  AND U3734 ( .A(n3789), .B(n3790), .Z(n3788) );
  XNOR U3735 ( .A(p_input[543]), .B(n3787), .Z(n3790) );
  XOR U3736 ( .A(n3787), .B(p_input[527]), .Z(n3789) );
  XOR U3737 ( .A(n3791), .B(n3792), .Z(n3787) );
  AND U3738 ( .A(n3793), .B(n3794), .Z(n3792) );
  XNOR U3739 ( .A(p_input[542]), .B(n3791), .Z(n3794) );
  XNOR U3740 ( .A(n3791), .B(n3601), .Z(n3793) );
  IV U3741 ( .A(p_input[526]), .Z(n3601) );
  XOR U3742 ( .A(n3795), .B(n3796), .Z(n3791) );
  AND U3743 ( .A(n3797), .B(n3798), .Z(n3796) );
  XNOR U3744 ( .A(p_input[541]), .B(n3795), .Z(n3798) );
  XNOR U3745 ( .A(n3795), .B(n3610), .Z(n3797) );
  IV U3746 ( .A(p_input[525]), .Z(n3610) );
  XOR U3747 ( .A(n3799), .B(n3800), .Z(n3795) );
  AND U3748 ( .A(n3801), .B(n3802), .Z(n3800) );
  XNOR U3749 ( .A(p_input[540]), .B(n3799), .Z(n3802) );
  XNOR U3750 ( .A(n3799), .B(n3619), .Z(n3801) );
  IV U3751 ( .A(p_input[524]), .Z(n3619) );
  XOR U3752 ( .A(n3803), .B(n3804), .Z(n3799) );
  AND U3753 ( .A(n3805), .B(n3806), .Z(n3804) );
  XNOR U3754 ( .A(p_input[539]), .B(n3803), .Z(n3806) );
  XNOR U3755 ( .A(n3803), .B(n3628), .Z(n3805) );
  IV U3756 ( .A(p_input[523]), .Z(n3628) );
  XOR U3757 ( .A(n3807), .B(n3808), .Z(n3803) );
  AND U3758 ( .A(n3809), .B(n3810), .Z(n3808) );
  XNOR U3759 ( .A(p_input[538]), .B(n3807), .Z(n3810) );
  XNOR U3760 ( .A(n3807), .B(n3637), .Z(n3809) );
  IV U3761 ( .A(p_input[522]), .Z(n3637) );
  XOR U3762 ( .A(n3811), .B(n3812), .Z(n3807) );
  AND U3763 ( .A(n3813), .B(n3814), .Z(n3812) );
  XNOR U3764 ( .A(p_input[537]), .B(n3811), .Z(n3814) );
  XNOR U3765 ( .A(n3811), .B(n3646), .Z(n3813) );
  IV U3766 ( .A(p_input[521]), .Z(n3646) );
  XOR U3767 ( .A(n3815), .B(n3816), .Z(n3811) );
  AND U3768 ( .A(n3817), .B(n3818), .Z(n3816) );
  XNOR U3769 ( .A(p_input[536]), .B(n3815), .Z(n3818) );
  XNOR U3770 ( .A(n3815), .B(n3655), .Z(n3817) );
  IV U3771 ( .A(p_input[520]), .Z(n3655) );
  XOR U3772 ( .A(n3819), .B(n3820), .Z(n3815) );
  AND U3773 ( .A(n3821), .B(n3822), .Z(n3820) );
  XNOR U3774 ( .A(p_input[535]), .B(n3819), .Z(n3822) );
  XNOR U3775 ( .A(n3819), .B(n3664), .Z(n3821) );
  IV U3776 ( .A(p_input[519]), .Z(n3664) );
  XOR U3777 ( .A(n3823), .B(n3824), .Z(n3819) );
  AND U3778 ( .A(n3825), .B(n3826), .Z(n3824) );
  XNOR U3779 ( .A(p_input[534]), .B(n3823), .Z(n3826) );
  XNOR U3780 ( .A(n3823), .B(n3673), .Z(n3825) );
  IV U3781 ( .A(p_input[518]), .Z(n3673) );
  XOR U3782 ( .A(n3827), .B(n3828), .Z(n3823) );
  AND U3783 ( .A(n3829), .B(n3830), .Z(n3828) );
  XNOR U3784 ( .A(p_input[533]), .B(n3827), .Z(n3830) );
  XNOR U3785 ( .A(n3827), .B(n3682), .Z(n3829) );
  IV U3786 ( .A(p_input[517]), .Z(n3682) );
  XOR U3787 ( .A(n3831), .B(n3832), .Z(n3827) );
  AND U3788 ( .A(n3833), .B(n3834), .Z(n3832) );
  XNOR U3789 ( .A(p_input[532]), .B(n3831), .Z(n3834) );
  XNOR U3790 ( .A(n3831), .B(n3691), .Z(n3833) );
  IV U3791 ( .A(p_input[516]), .Z(n3691) );
  XOR U3792 ( .A(n3835), .B(n3836), .Z(n3831) );
  AND U3793 ( .A(n3837), .B(n3838), .Z(n3836) );
  XNOR U3794 ( .A(p_input[531]), .B(n3835), .Z(n3838) );
  XNOR U3795 ( .A(n3835), .B(n3700), .Z(n3837) );
  IV U3796 ( .A(p_input[515]), .Z(n3700) );
  XOR U3797 ( .A(n3839), .B(n3840), .Z(n3835) );
  AND U3798 ( .A(n3841), .B(n3842), .Z(n3840) );
  XNOR U3799 ( .A(p_input[530]), .B(n3839), .Z(n3842) );
  XNOR U3800 ( .A(n3839), .B(n3709), .Z(n3841) );
  IV U3801 ( .A(p_input[514]), .Z(n3709) );
  XNOR U3802 ( .A(n3843), .B(n3844), .Z(n3839) );
  AND U3803 ( .A(n3845), .B(n3846), .Z(n3844) );
  XOR U3804 ( .A(p_input[529]), .B(n3843), .Z(n3846) );
  XNOR U3805 ( .A(p_input[513]), .B(n3843), .Z(n3845) );
  AND U3806 ( .A(p_input[528]), .B(n3847), .Z(n3843) );
  IV U3807 ( .A(p_input[512]), .Z(n3847) );
  XOR U3808 ( .A(n3848), .B(n3849), .Z(n16) );
  AND U3809 ( .A(n299), .B(n3850), .Z(n3849) );
  XNOR U3810 ( .A(n3851), .B(n3848), .Z(n3850) );
  XOR U3811 ( .A(n3852), .B(n3853), .Z(n299) );
  AND U3812 ( .A(n3854), .B(n3855), .Z(n3853) );
  XOR U3813 ( .A(n3852), .B(n318), .Z(n3855) );
  XNOR U3814 ( .A(n3856), .B(n3857), .Z(n318) );
  AND U3815 ( .A(n3858), .B(n290), .Z(n3857) );
  AND U3816 ( .A(n3856), .B(n3859), .Z(n3858) );
  XNOR U3817 ( .A(n315), .B(n3852), .Z(n3854) );
  XOR U3818 ( .A(n3860), .B(n3861), .Z(n315) );
  AND U3819 ( .A(n3862), .B(n287), .Z(n3861) );
  NOR U3820 ( .A(n3860), .B(n3863), .Z(n3862) );
  XOR U3821 ( .A(n3864), .B(n3865), .Z(n3852) );
  AND U3822 ( .A(n3866), .B(n3867), .Z(n3865) );
  XOR U3823 ( .A(n3864), .B(n330), .Z(n3867) );
  XOR U3824 ( .A(n3868), .B(n3869), .Z(n330) );
  AND U3825 ( .A(n290), .B(n3870), .Z(n3869) );
  XOR U3826 ( .A(n3871), .B(n3868), .Z(n3870) );
  XNOR U3827 ( .A(n327), .B(n3864), .Z(n3866) );
  XOR U3828 ( .A(n3872), .B(n3873), .Z(n327) );
  AND U3829 ( .A(n287), .B(n3874), .Z(n3873) );
  XOR U3830 ( .A(n3875), .B(n3872), .Z(n3874) );
  XOR U3831 ( .A(n3876), .B(n3877), .Z(n3864) );
  AND U3832 ( .A(n3878), .B(n3879), .Z(n3877) );
  XOR U3833 ( .A(n3876), .B(n342), .Z(n3879) );
  XOR U3834 ( .A(n3880), .B(n3881), .Z(n342) );
  AND U3835 ( .A(n290), .B(n3882), .Z(n3881) );
  XOR U3836 ( .A(n3883), .B(n3880), .Z(n3882) );
  XNOR U3837 ( .A(n339), .B(n3876), .Z(n3878) );
  XOR U3838 ( .A(n3884), .B(n3885), .Z(n339) );
  AND U3839 ( .A(n287), .B(n3886), .Z(n3885) );
  XOR U3840 ( .A(n3887), .B(n3884), .Z(n3886) );
  XOR U3841 ( .A(n3888), .B(n3889), .Z(n3876) );
  AND U3842 ( .A(n3890), .B(n3891), .Z(n3889) );
  XOR U3843 ( .A(n3888), .B(n354), .Z(n3891) );
  XOR U3844 ( .A(n3892), .B(n3893), .Z(n354) );
  AND U3845 ( .A(n290), .B(n3894), .Z(n3893) );
  XOR U3846 ( .A(n3895), .B(n3892), .Z(n3894) );
  XNOR U3847 ( .A(n351), .B(n3888), .Z(n3890) );
  XOR U3848 ( .A(n3896), .B(n3897), .Z(n351) );
  AND U3849 ( .A(n287), .B(n3898), .Z(n3897) );
  XOR U3850 ( .A(n3899), .B(n3896), .Z(n3898) );
  XOR U3851 ( .A(n3900), .B(n3901), .Z(n3888) );
  AND U3852 ( .A(n3902), .B(n3903), .Z(n3901) );
  XOR U3853 ( .A(n3900), .B(n366), .Z(n3903) );
  XOR U3854 ( .A(n3904), .B(n3905), .Z(n366) );
  AND U3855 ( .A(n290), .B(n3906), .Z(n3905) );
  XOR U3856 ( .A(n3907), .B(n3904), .Z(n3906) );
  XNOR U3857 ( .A(n363), .B(n3900), .Z(n3902) );
  XOR U3858 ( .A(n3908), .B(n3909), .Z(n363) );
  AND U3859 ( .A(n287), .B(n3910), .Z(n3909) );
  XOR U3860 ( .A(n3911), .B(n3908), .Z(n3910) );
  XOR U3861 ( .A(n3912), .B(n3913), .Z(n3900) );
  AND U3862 ( .A(n3914), .B(n3915), .Z(n3913) );
  XOR U3863 ( .A(n3912), .B(n378), .Z(n3915) );
  XOR U3864 ( .A(n3916), .B(n3917), .Z(n378) );
  AND U3865 ( .A(n290), .B(n3918), .Z(n3917) );
  XOR U3866 ( .A(n3919), .B(n3916), .Z(n3918) );
  XNOR U3867 ( .A(n375), .B(n3912), .Z(n3914) );
  XOR U3868 ( .A(n3920), .B(n3921), .Z(n375) );
  AND U3869 ( .A(n287), .B(n3922), .Z(n3921) );
  XOR U3870 ( .A(n3923), .B(n3920), .Z(n3922) );
  XOR U3871 ( .A(n3924), .B(n3925), .Z(n3912) );
  AND U3872 ( .A(n3926), .B(n3927), .Z(n3925) );
  XOR U3873 ( .A(n3924), .B(n390), .Z(n3927) );
  XOR U3874 ( .A(n3928), .B(n3929), .Z(n390) );
  AND U3875 ( .A(n290), .B(n3930), .Z(n3929) );
  XOR U3876 ( .A(n3931), .B(n3928), .Z(n3930) );
  XNOR U3877 ( .A(n387), .B(n3924), .Z(n3926) );
  XOR U3878 ( .A(n3932), .B(n3933), .Z(n387) );
  AND U3879 ( .A(n287), .B(n3934), .Z(n3933) );
  XOR U3880 ( .A(n3935), .B(n3932), .Z(n3934) );
  XOR U3881 ( .A(n3936), .B(n3937), .Z(n3924) );
  AND U3882 ( .A(n3938), .B(n3939), .Z(n3937) );
  XOR U3883 ( .A(n3936), .B(n402), .Z(n3939) );
  XOR U3884 ( .A(n3940), .B(n3941), .Z(n402) );
  AND U3885 ( .A(n290), .B(n3942), .Z(n3941) );
  XOR U3886 ( .A(n3943), .B(n3940), .Z(n3942) );
  XNOR U3887 ( .A(n399), .B(n3936), .Z(n3938) );
  XOR U3888 ( .A(n3944), .B(n3945), .Z(n399) );
  AND U3889 ( .A(n287), .B(n3946), .Z(n3945) );
  XOR U3890 ( .A(n3947), .B(n3944), .Z(n3946) );
  XOR U3891 ( .A(n3948), .B(n3949), .Z(n3936) );
  AND U3892 ( .A(n3950), .B(n3951), .Z(n3949) );
  XOR U3893 ( .A(n3948), .B(n414), .Z(n3951) );
  XOR U3894 ( .A(n3952), .B(n3953), .Z(n414) );
  AND U3895 ( .A(n290), .B(n3954), .Z(n3953) );
  XOR U3896 ( .A(n3955), .B(n3952), .Z(n3954) );
  XNOR U3897 ( .A(n411), .B(n3948), .Z(n3950) );
  XOR U3898 ( .A(n3956), .B(n3957), .Z(n411) );
  AND U3899 ( .A(n287), .B(n3958), .Z(n3957) );
  XOR U3900 ( .A(n3959), .B(n3956), .Z(n3958) );
  XOR U3901 ( .A(n3960), .B(n3961), .Z(n3948) );
  AND U3902 ( .A(n3962), .B(n3963), .Z(n3961) );
  XOR U3903 ( .A(n3960), .B(n426), .Z(n3963) );
  XOR U3904 ( .A(n3964), .B(n3965), .Z(n426) );
  AND U3905 ( .A(n290), .B(n3966), .Z(n3965) );
  XOR U3906 ( .A(n3967), .B(n3964), .Z(n3966) );
  XNOR U3907 ( .A(n423), .B(n3960), .Z(n3962) );
  XOR U3908 ( .A(n3968), .B(n3969), .Z(n423) );
  AND U3909 ( .A(n287), .B(n3970), .Z(n3969) );
  XOR U3910 ( .A(n3971), .B(n3968), .Z(n3970) );
  XOR U3911 ( .A(n3972), .B(n3973), .Z(n3960) );
  AND U3912 ( .A(n3974), .B(n3975), .Z(n3973) );
  XOR U3913 ( .A(n3972), .B(n438), .Z(n3975) );
  XOR U3914 ( .A(n3976), .B(n3977), .Z(n438) );
  AND U3915 ( .A(n290), .B(n3978), .Z(n3977) );
  XOR U3916 ( .A(n3979), .B(n3976), .Z(n3978) );
  XNOR U3917 ( .A(n435), .B(n3972), .Z(n3974) );
  XOR U3918 ( .A(n3980), .B(n3981), .Z(n435) );
  AND U3919 ( .A(n287), .B(n3982), .Z(n3981) );
  XOR U3920 ( .A(n3983), .B(n3980), .Z(n3982) );
  XOR U3921 ( .A(n3984), .B(n3985), .Z(n3972) );
  AND U3922 ( .A(n3986), .B(n3987), .Z(n3985) );
  XOR U3923 ( .A(n3984), .B(n450), .Z(n3987) );
  XOR U3924 ( .A(n3988), .B(n3989), .Z(n450) );
  AND U3925 ( .A(n290), .B(n3990), .Z(n3989) );
  XOR U3926 ( .A(n3991), .B(n3988), .Z(n3990) );
  XNOR U3927 ( .A(n447), .B(n3984), .Z(n3986) );
  XOR U3928 ( .A(n3992), .B(n3993), .Z(n447) );
  AND U3929 ( .A(n287), .B(n3994), .Z(n3993) );
  XOR U3930 ( .A(n3995), .B(n3992), .Z(n3994) );
  XOR U3931 ( .A(n3996), .B(n3997), .Z(n3984) );
  AND U3932 ( .A(n3998), .B(n3999), .Z(n3997) );
  XOR U3933 ( .A(n462), .B(n3996), .Z(n3999) );
  XOR U3934 ( .A(n4000), .B(n4001), .Z(n462) );
  AND U3935 ( .A(n290), .B(n4002), .Z(n4001) );
  XOR U3936 ( .A(n4000), .B(n4003), .Z(n4002) );
  XNOR U3937 ( .A(n3996), .B(n459), .Z(n3998) );
  XOR U3938 ( .A(n4004), .B(n4005), .Z(n459) );
  AND U3939 ( .A(n287), .B(n4006), .Z(n4005) );
  XOR U3940 ( .A(n4004), .B(n4007), .Z(n4006) );
  XOR U3941 ( .A(n4008), .B(n4009), .Z(n3996) );
  AND U3942 ( .A(n4010), .B(n4011), .Z(n4009) );
  XOR U3943 ( .A(n4008), .B(n474), .Z(n4011) );
  XOR U3944 ( .A(n4012), .B(n4013), .Z(n474) );
  AND U3945 ( .A(n290), .B(n4014), .Z(n4013) );
  XOR U3946 ( .A(n4015), .B(n4012), .Z(n4014) );
  XNOR U3947 ( .A(n471), .B(n4008), .Z(n4010) );
  XOR U3948 ( .A(n4016), .B(n4017), .Z(n471) );
  AND U3949 ( .A(n287), .B(n4018), .Z(n4017) );
  XOR U3950 ( .A(n4019), .B(n4016), .Z(n4018) );
  XOR U3951 ( .A(n4020), .B(n4021), .Z(n4008) );
  AND U3952 ( .A(n4022), .B(n4023), .Z(n4021) );
  XNOR U3953 ( .A(n4024), .B(n486), .Z(n4023) );
  XOR U3954 ( .A(n4025), .B(n4026), .Z(n486) );
  AND U3955 ( .A(n290), .B(n4027), .Z(n4026) );
  XOR U3956 ( .A(n4028), .B(n4025), .Z(n4027) );
  XNOR U3957 ( .A(n483), .B(n4020), .Z(n4022) );
  XOR U3958 ( .A(n4029), .B(n4030), .Z(n483) );
  AND U3959 ( .A(n287), .B(n4031), .Z(n4030) );
  XOR U3960 ( .A(n4032), .B(n4029), .Z(n4031) );
  IV U3961 ( .A(n4024), .Z(n4020) );
  AND U3962 ( .A(n3848), .B(n3851), .Z(n4024) );
  XNOR U3963 ( .A(n4033), .B(n4034), .Z(n3851) );
  AND U3964 ( .A(n290), .B(n4035), .Z(n4034) );
  XNOR U3965 ( .A(n4036), .B(n4033), .Z(n4035) );
  XOR U3966 ( .A(n4037), .B(n4038), .Z(n290) );
  AND U3967 ( .A(n4039), .B(n4040), .Z(n4038) );
  XOR U3968 ( .A(n3859), .B(n4037), .Z(n4040) );
  IV U3969 ( .A(n4041), .Z(n3859) );
  AND U3970 ( .A(n4042), .B(n4043), .Z(n4041) );
  XOR U3971 ( .A(n4037), .B(n3856), .Z(n4039) );
  AND U3972 ( .A(n4044), .B(n4045), .Z(n3856) );
  XOR U3973 ( .A(n4046), .B(n4047), .Z(n4037) );
  AND U3974 ( .A(n4048), .B(n4049), .Z(n4047) );
  XOR U3975 ( .A(n4046), .B(n3871), .Z(n4049) );
  XOR U3976 ( .A(n4050), .B(n4051), .Z(n3871) );
  AND U3977 ( .A(n258), .B(n4052), .Z(n4051) );
  XOR U3978 ( .A(n4053), .B(n4050), .Z(n4052) );
  XNOR U3979 ( .A(n3868), .B(n4046), .Z(n4048) );
  XOR U3980 ( .A(n4054), .B(n4055), .Z(n3868) );
  AND U3981 ( .A(n256), .B(n4056), .Z(n4055) );
  XOR U3982 ( .A(n4057), .B(n4054), .Z(n4056) );
  XOR U3983 ( .A(n4058), .B(n4059), .Z(n4046) );
  AND U3984 ( .A(n4060), .B(n4061), .Z(n4059) );
  XOR U3985 ( .A(n4058), .B(n3883), .Z(n4061) );
  XOR U3986 ( .A(n4062), .B(n4063), .Z(n3883) );
  AND U3987 ( .A(n258), .B(n4064), .Z(n4063) );
  XOR U3988 ( .A(n4065), .B(n4062), .Z(n4064) );
  XNOR U3989 ( .A(n3880), .B(n4058), .Z(n4060) );
  XOR U3990 ( .A(n4066), .B(n4067), .Z(n3880) );
  AND U3991 ( .A(n256), .B(n4068), .Z(n4067) );
  XOR U3992 ( .A(n4069), .B(n4066), .Z(n4068) );
  XOR U3993 ( .A(n4070), .B(n4071), .Z(n4058) );
  AND U3994 ( .A(n4072), .B(n4073), .Z(n4071) );
  XOR U3995 ( .A(n4070), .B(n3895), .Z(n4073) );
  XOR U3996 ( .A(n4074), .B(n4075), .Z(n3895) );
  AND U3997 ( .A(n258), .B(n4076), .Z(n4075) );
  XOR U3998 ( .A(n4077), .B(n4074), .Z(n4076) );
  XNOR U3999 ( .A(n3892), .B(n4070), .Z(n4072) );
  XOR U4000 ( .A(n4078), .B(n4079), .Z(n3892) );
  AND U4001 ( .A(n256), .B(n4080), .Z(n4079) );
  XOR U4002 ( .A(n4081), .B(n4078), .Z(n4080) );
  XOR U4003 ( .A(n4082), .B(n4083), .Z(n4070) );
  AND U4004 ( .A(n4084), .B(n4085), .Z(n4083) );
  XOR U4005 ( .A(n4082), .B(n3907), .Z(n4085) );
  XOR U4006 ( .A(n4086), .B(n4087), .Z(n3907) );
  AND U4007 ( .A(n258), .B(n4088), .Z(n4087) );
  XOR U4008 ( .A(n4089), .B(n4086), .Z(n4088) );
  XNOR U4009 ( .A(n3904), .B(n4082), .Z(n4084) );
  XOR U4010 ( .A(n4090), .B(n4091), .Z(n3904) );
  AND U4011 ( .A(n256), .B(n4092), .Z(n4091) );
  XOR U4012 ( .A(n4093), .B(n4090), .Z(n4092) );
  XOR U4013 ( .A(n4094), .B(n4095), .Z(n4082) );
  AND U4014 ( .A(n4096), .B(n4097), .Z(n4095) );
  XOR U4015 ( .A(n4094), .B(n3919), .Z(n4097) );
  XOR U4016 ( .A(n4098), .B(n4099), .Z(n3919) );
  AND U4017 ( .A(n258), .B(n4100), .Z(n4099) );
  XOR U4018 ( .A(n4101), .B(n4098), .Z(n4100) );
  XNOR U4019 ( .A(n3916), .B(n4094), .Z(n4096) );
  XOR U4020 ( .A(n4102), .B(n4103), .Z(n3916) );
  AND U4021 ( .A(n256), .B(n4104), .Z(n4103) );
  XOR U4022 ( .A(n4105), .B(n4102), .Z(n4104) );
  XOR U4023 ( .A(n4106), .B(n4107), .Z(n4094) );
  AND U4024 ( .A(n4108), .B(n4109), .Z(n4107) );
  XOR U4025 ( .A(n4106), .B(n3931), .Z(n4109) );
  XOR U4026 ( .A(n4110), .B(n4111), .Z(n3931) );
  AND U4027 ( .A(n258), .B(n4112), .Z(n4111) );
  XOR U4028 ( .A(n4113), .B(n4110), .Z(n4112) );
  XNOR U4029 ( .A(n3928), .B(n4106), .Z(n4108) );
  XOR U4030 ( .A(n4114), .B(n4115), .Z(n3928) );
  AND U4031 ( .A(n256), .B(n4116), .Z(n4115) );
  XOR U4032 ( .A(n4117), .B(n4114), .Z(n4116) );
  XOR U4033 ( .A(n4118), .B(n4119), .Z(n4106) );
  AND U4034 ( .A(n4120), .B(n4121), .Z(n4119) );
  XOR U4035 ( .A(n4118), .B(n3943), .Z(n4121) );
  XOR U4036 ( .A(n4122), .B(n4123), .Z(n3943) );
  AND U4037 ( .A(n258), .B(n4124), .Z(n4123) );
  XOR U4038 ( .A(n4125), .B(n4122), .Z(n4124) );
  XNOR U4039 ( .A(n3940), .B(n4118), .Z(n4120) );
  XOR U4040 ( .A(n4126), .B(n4127), .Z(n3940) );
  AND U4041 ( .A(n256), .B(n4128), .Z(n4127) );
  XOR U4042 ( .A(n4129), .B(n4126), .Z(n4128) );
  XOR U4043 ( .A(n4130), .B(n4131), .Z(n4118) );
  AND U4044 ( .A(n4132), .B(n4133), .Z(n4131) );
  XOR U4045 ( .A(n4130), .B(n3955), .Z(n4133) );
  XOR U4046 ( .A(n4134), .B(n4135), .Z(n3955) );
  AND U4047 ( .A(n258), .B(n4136), .Z(n4135) );
  XOR U4048 ( .A(n4137), .B(n4134), .Z(n4136) );
  XNOR U4049 ( .A(n3952), .B(n4130), .Z(n4132) );
  XOR U4050 ( .A(n4138), .B(n4139), .Z(n3952) );
  AND U4051 ( .A(n256), .B(n4140), .Z(n4139) );
  XOR U4052 ( .A(n4141), .B(n4138), .Z(n4140) );
  XOR U4053 ( .A(n4142), .B(n4143), .Z(n4130) );
  AND U4054 ( .A(n4144), .B(n4145), .Z(n4143) );
  XOR U4055 ( .A(n4142), .B(n3967), .Z(n4145) );
  XOR U4056 ( .A(n4146), .B(n4147), .Z(n3967) );
  AND U4057 ( .A(n258), .B(n4148), .Z(n4147) );
  XOR U4058 ( .A(n4149), .B(n4146), .Z(n4148) );
  XNOR U4059 ( .A(n3964), .B(n4142), .Z(n4144) );
  XOR U4060 ( .A(n4150), .B(n4151), .Z(n3964) );
  AND U4061 ( .A(n256), .B(n4152), .Z(n4151) );
  XOR U4062 ( .A(n4153), .B(n4150), .Z(n4152) );
  XOR U4063 ( .A(n4154), .B(n4155), .Z(n4142) );
  AND U4064 ( .A(n4156), .B(n4157), .Z(n4155) );
  XOR U4065 ( .A(n4154), .B(n3979), .Z(n4157) );
  XOR U4066 ( .A(n4158), .B(n4159), .Z(n3979) );
  AND U4067 ( .A(n258), .B(n4160), .Z(n4159) );
  XOR U4068 ( .A(n4161), .B(n4158), .Z(n4160) );
  XNOR U4069 ( .A(n3976), .B(n4154), .Z(n4156) );
  XOR U4070 ( .A(n4162), .B(n4163), .Z(n3976) );
  AND U4071 ( .A(n256), .B(n4164), .Z(n4163) );
  XOR U4072 ( .A(n4165), .B(n4162), .Z(n4164) );
  XOR U4073 ( .A(n4166), .B(n4167), .Z(n4154) );
  AND U4074 ( .A(n4168), .B(n4169), .Z(n4167) );
  XOR U4075 ( .A(n4166), .B(n3991), .Z(n4169) );
  XOR U4076 ( .A(n4170), .B(n4171), .Z(n3991) );
  AND U4077 ( .A(n258), .B(n4172), .Z(n4171) );
  XOR U4078 ( .A(n4173), .B(n4170), .Z(n4172) );
  XNOR U4079 ( .A(n3988), .B(n4166), .Z(n4168) );
  XOR U4080 ( .A(n4174), .B(n4175), .Z(n3988) );
  AND U4081 ( .A(n256), .B(n4176), .Z(n4175) );
  XOR U4082 ( .A(n4177), .B(n4174), .Z(n4176) );
  XOR U4083 ( .A(n4178), .B(n4179), .Z(n4166) );
  AND U4084 ( .A(n4180), .B(n4181), .Z(n4179) );
  XOR U4085 ( .A(n4003), .B(n4178), .Z(n4181) );
  XOR U4086 ( .A(n4182), .B(n4183), .Z(n4003) );
  AND U4087 ( .A(n258), .B(n4184), .Z(n4183) );
  XOR U4088 ( .A(n4182), .B(n4185), .Z(n4184) );
  XNOR U4089 ( .A(n4178), .B(n4000), .Z(n4180) );
  XOR U4090 ( .A(n4186), .B(n4187), .Z(n4000) );
  AND U4091 ( .A(n256), .B(n4188), .Z(n4187) );
  XOR U4092 ( .A(n4186), .B(n4189), .Z(n4188) );
  XOR U4093 ( .A(n4190), .B(n4191), .Z(n4178) );
  AND U4094 ( .A(n4192), .B(n4193), .Z(n4191) );
  XOR U4095 ( .A(n4190), .B(n4015), .Z(n4193) );
  XOR U4096 ( .A(n4194), .B(n4195), .Z(n4015) );
  AND U4097 ( .A(n258), .B(n4196), .Z(n4195) );
  XOR U4098 ( .A(n4197), .B(n4194), .Z(n4196) );
  XNOR U4099 ( .A(n4012), .B(n4190), .Z(n4192) );
  XOR U4100 ( .A(n4198), .B(n4199), .Z(n4012) );
  AND U4101 ( .A(n256), .B(n4200), .Z(n4199) );
  XOR U4102 ( .A(n4201), .B(n4198), .Z(n4200) );
  XOR U4103 ( .A(n4202), .B(n4203), .Z(n4190) );
  AND U4104 ( .A(n4204), .B(n4205), .Z(n4203) );
  XNOR U4105 ( .A(n4206), .B(n4028), .Z(n4205) );
  XOR U4106 ( .A(n4207), .B(n4208), .Z(n4028) );
  AND U4107 ( .A(n258), .B(n4209), .Z(n4208) );
  XOR U4108 ( .A(n4210), .B(n4207), .Z(n4209) );
  XNOR U4109 ( .A(n4025), .B(n4202), .Z(n4204) );
  XOR U4110 ( .A(n4211), .B(n4212), .Z(n4025) );
  AND U4111 ( .A(n256), .B(n4213), .Z(n4212) );
  XOR U4112 ( .A(n4214), .B(n4211), .Z(n4213) );
  IV U4113 ( .A(n4206), .Z(n4202) );
  AND U4114 ( .A(n4033), .B(n4036), .Z(n4206) );
  XNOR U4115 ( .A(n4215), .B(n4216), .Z(n4036) );
  AND U4116 ( .A(n258), .B(n4217), .Z(n4216) );
  XNOR U4117 ( .A(n4218), .B(n4215), .Z(n4217) );
  XOR U4118 ( .A(n4219), .B(n4220), .Z(n258) );
  AND U4119 ( .A(n4221), .B(n4222), .Z(n4220) );
  XNOR U4120 ( .A(n4042), .B(n4219), .Z(n4222) );
  AND U4121 ( .A(n4223), .B(n4224), .Z(n4042) );
  XOR U4122 ( .A(n4219), .B(n4043), .Z(n4221) );
  AND U4123 ( .A(n4225), .B(n4226), .Z(n4043) );
  XOR U4124 ( .A(n4227), .B(n4228), .Z(n4219) );
  AND U4125 ( .A(n4229), .B(n4230), .Z(n4228) );
  XOR U4126 ( .A(n4227), .B(n4053), .Z(n4230) );
  XOR U4127 ( .A(n4231), .B(n4232), .Z(n4053) );
  AND U4128 ( .A(n186), .B(n4233), .Z(n4232) );
  XOR U4129 ( .A(n4234), .B(n4231), .Z(n4233) );
  XNOR U4130 ( .A(n4050), .B(n4227), .Z(n4229) );
  XOR U4131 ( .A(n4235), .B(n4236), .Z(n4050) );
  AND U4132 ( .A(n184), .B(n4237), .Z(n4236) );
  XOR U4133 ( .A(n4238), .B(n4235), .Z(n4237) );
  XOR U4134 ( .A(n4239), .B(n4240), .Z(n4227) );
  AND U4135 ( .A(n4241), .B(n4242), .Z(n4240) );
  XOR U4136 ( .A(n4239), .B(n4065), .Z(n4242) );
  XOR U4137 ( .A(n4243), .B(n4244), .Z(n4065) );
  AND U4138 ( .A(n186), .B(n4245), .Z(n4244) );
  XOR U4139 ( .A(n4246), .B(n4243), .Z(n4245) );
  XNOR U4140 ( .A(n4062), .B(n4239), .Z(n4241) );
  XOR U4141 ( .A(n4247), .B(n4248), .Z(n4062) );
  AND U4142 ( .A(n184), .B(n4249), .Z(n4248) );
  XOR U4143 ( .A(n4250), .B(n4247), .Z(n4249) );
  XOR U4144 ( .A(n4251), .B(n4252), .Z(n4239) );
  AND U4145 ( .A(n4253), .B(n4254), .Z(n4252) );
  XOR U4146 ( .A(n4251), .B(n4077), .Z(n4254) );
  XOR U4147 ( .A(n4255), .B(n4256), .Z(n4077) );
  AND U4148 ( .A(n186), .B(n4257), .Z(n4256) );
  XOR U4149 ( .A(n4258), .B(n4255), .Z(n4257) );
  XNOR U4150 ( .A(n4074), .B(n4251), .Z(n4253) );
  XOR U4151 ( .A(n4259), .B(n4260), .Z(n4074) );
  AND U4152 ( .A(n184), .B(n4261), .Z(n4260) );
  XOR U4153 ( .A(n4262), .B(n4259), .Z(n4261) );
  XOR U4154 ( .A(n4263), .B(n4264), .Z(n4251) );
  AND U4155 ( .A(n4265), .B(n4266), .Z(n4264) );
  XOR U4156 ( .A(n4263), .B(n4089), .Z(n4266) );
  XOR U4157 ( .A(n4267), .B(n4268), .Z(n4089) );
  AND U4158 ( .A(n186), .B(n4269), .Z(n4268) );
  XOR U4159 ( .A(n4270), .B(n4267), .Z(n4269) );
  XNOR U4160 ( .A(n4086), .B(n4263), .Z(n4265) );
  XOR U4161 ( .A(n4271), .B(n4272), .Z(n4086) );
  AND U4162 ( .A(n184), .B(n4273), .Z(n4272) );
  XOR U4163 ( .A(n4274), .B(n4271), .Z(n4273) );
  XOR U4164 ( .A(n4275), .B(n4276), .Z(n4263) );
  AND U4165 ( .A(n4277), .B(n4278), .Z(n4276) );
  XOR U4166 ( .A(n4275), .B(n4101), .Z(n4278) );
  XOR U4167 ( .A(n4279), .B(n4280), .Z(n4101) );
  AND U4168 ( .A(n186), .B(n4281), .Z(n4280) );
  XOR U4169 ( .A(n4282), .B(n4279), .Z(n4281) );
  XNOR U4170 ( .A(n4098), .B(n4275), .Z(n4277) );
  XOR U4171 ( .A(n4283), .B(n4284), .Z(n4098) );
  AND U4172 ( .A(n184), .B(n4285), .Z(n4284) );
  XOR U4173 ( .A(n4286), .B(n4283), .Z(n4285) );
  XOR U4174 ( .A(n4287), .B(n4288), .Z(n4275) );
  AND U4175 ( .A(n4289), .B(n4290), .Z(n4288) );
  XOR U4176 ( .A(n4287), .B(n4113), .Z(n4290) );
  XOR U4177 ( .A(n4291), .B(n4292), .Z(n4113) );
  AND U4178 ( .A(n186), .B(n4293), .Z(n4292) );
  XOR U4179 ( .A(n4294), .B(n4291), .Z(n4293) );
  XNOR U4180 ( .A(n4110), .B(n4287), .Z(n4289) );
  XOR U4181 ( .A(n4295), .B(n4296), .Z(n4110) );
  AND U4182 ( .A(n184), .B(n4297), .Z(n4296) );
  XOR U4183 ( .A(n4298), .B(n4295), .Z(n4297) );
  XOR U4184 ( .A(n4299), .B(n4300), .Z(n4287) );
  AND U4185 ( .A(n4301), .B(n4302), .Z(n4300) );
  XOR U4186 ( .A(n4299), .B(n4125), .Z(n4302) );
  XOR U4187 ( .A(n4303), .B(n4304), .Z(n4125) );
  AND U4188 ( .A(n186), .B(n4305), .Z(n4304) );
  XOR U4189 ( .A(n4306), .B(n4303), .Z(n4305) );
  XNOR U4190 ( .A(n4122), .B(n4299), .Z(n4301) );
  XOR U4191 ( .A(n4307), .B(n4308), .Z(n4122) );
  AND U4192 ( .A(n184), .B(n4309), .Z(n4308) );
  XOR U4193 ( .A(n4310), .B(n4307), .Z(n4309) );
  XOR U4194 ( .A(n4311), .B(n4312), .Z(n4299) );
  AND U4195 ( .A(n4313), .B(n4314), .Z(n4312) );
  XOR U4196 ( .A(n4311), .B(n4137), .Z(n4314) );
  XOR U4197 ( .A(n4315), .B(n4316), .Z(n4137) );
  AND U4198 ( .A(n186), .B(n4317), .Z(n4316) );
  XOR U4199 ( .A(n4318), .B(n4315), .Z(n4317) );
  XNOR U4200 ( .A(n4134), .B(n4311), .Z(n4313) );
  XOR U4201 ( .A(n4319), .B(n4320), .Z(n4134) );
  AND U4202 ( .A(n184), .B(n4321), .Z(n4320) );
  XOR U4203 ( .A(n4322), .B(n4319), .Z(n4321) );
  XOR U4204 ( .A(n4323), .B(n4324), .Z(n4311) );
  AND U4205 ( .A(n4325), .B(n4326), .Z(n4324) );
  XOR U4206 ( .A(n4323), .B(n4149), .Z(n4326) );
  XOR U4207 ( .A(n4327), .B(n4328), .Z(n4149) );
  AND U4208 ( .A(n186), .B(n4329), .Z(n4328) );
  XOR U4209 ( .A(n4330), .B(n4327), .Z(n4329) );
  XNOR U4210 ( .A(n4146), .B(n4323), .Z(n4325) );
  XOR U4211 ( .A(n4331), .B(n4332), .Z(n4146) );
  AND U4212 ( .A(n184), .B(n4333), .Z(n4332) );
  XOR U4213 ( .A(n4334), .B(n4331), .Z(n4333) );
  XOR U4214 ( .A(n4335), .B(n4336), .Z(n4323) );
  AND U4215 ( .A(n4337), .B(n4338), .Z(n4336) );
  XOR U4216 ( .A(n4335), .B(n4161), .Z(n4338) );
  XOR U4217 ( .A(n4339), .B(n4340), .Z(n4161) );
  AND U4218 ( .A(n186), .B(n4341), .Z(n4340) );
  XOR U4219 ( .A(n4342), .B(n4339), .Z(n4341) );
  XNOR U4220 ( .A(n4158), .B(n4335), .Z(n4337) );
  XOR U4221 ( .A(n4343), .B(n4344), .Z(n4158) );
  AND U4222 ( .A(n184), .B(n4345), .Z(n4344) );
  XOR U4223 ( .A(n4346), .B(n4343), .Z(n4345) );
  XOR U4224 ( .A(n4347), .B(n4348), .Z(n4335) );
  AND U4225 ( .A(n4349), .B(n4350), .Z(n4348) );
  XOR U4226 ( .A(n4347), .B(n4173), .Z(n4350) );
  XOR U4227 ( .A(n4351), .B(n4352), .Z(n4173) );
  AND U4228 ( .A(n186), .B(n4353), .Z(n4352) );
  XOR U4229 ( .A(n4354), .B(n4351), .Z(n4353) );
  XNOR U4230 ( .A(n4170), .B(n4347), .Z(n4349) );
  XOR U4231 ( .A(n4355), .B(n4356), .Z(n4170) );
  AND U4232 ( .A(n184), .B(n4357), .Z(n4356) );
  XOR U4233 ( .A(n4358), .B(n4355), .Z(n4357) );
  XOR U4234 ( .A(n4359), .B(n4360), .Z(n4347) );
  AND U4235 ( .A(n4361), .B(n4362), .Z(n4360) );
  XOR U4236 ( .A(n4185), .B(n4359), .Z(n4362) );
  XOR U4237 ( .A(n4363), .B(n4364), .Z(n4185) );
  AND U4238 ( .A(n186), .B(n4365), .Z(n4364) );
  XOR U4239 ( .A(n4363), .B(n4366), .Z(n4365) );
  XNOR U4240 ( .A(n4359), .B(n4182), .Z(n4361) );
  XOR U4241 ( .A(n4367), .B(n4368), .Z(n4182) );
  AND U4242 ( .A(n184), .B(n4369), .Z(n4368) );
  XOR U4243 ( .A(n4367), .B(n4370), .Z(n4369) );
  XOR U4244 ( .A(n4371), .B(n4372), .Z(n4359) );
  AND U4245 ( .A(n4373), .B(n4374), .Z(n4372) );
  XOR U4246 ( .A(n4371), .B(n4197), .Z(n4374) );
  XOR U4247 ( .A(n4375), .B(n4376), .Z(n4197) );
  AND U4248 ( .A(n186), .B(n4377), .Z(n4376) );
  XOR U4249 ( .A(n4378), .B(n4375), .Z(n4377) );
  XNOR U4250 ( .A(n4194), .B(n4371), .Z(n4373) );
  XOR U4251 ( .A(n4379), .B(n4380), .Z(n4194) );
  AND U4252 ( .A(n184), .B(n4381), .Z(n4380) );
  XOR U4253 ( .A(n4382), .B(n4379), .Z(n4381) );
  XOR U4254 ( .A(n4383), .B(n4384), .Z(n4371) );
  AND U4255 ( .A(n4385), .B(n4386), .Z(n4384) );
  XNOR U4256 ( .A(n4387), .B(n4210), .Z(n4386) );
  XOR U4257 ( .A(n4388), .B(n4389), .Z(n4210) );
  AND U4258 ( .A(n186), .B(n4390), .Z(n4389) );
  XOR U4259 ( .A(n4391), .B(n4388), .Z(n4390) );
  XNOR U4260 ( .A(n4207), .B(n4383), .Z(n4385) );
  XOR U4261 ( .A(n4392), .B(n4393), .Z(n4207) );
  AND U4262 ( .A(n184), .B(n4394), .Z(n4393) );
  XOR U4263 ( .A(n4395), .B(n4392), .Z(n4394) );
  IV U4264 ( .A(n4387), .Z(n4383) );
  AND U4265 ( .A(n4215), .B(n4218), .Z(n4387) );
  XNOR U4266 ( .A(n4396), .B(n4397), .Z(n4218) );
  AND U4267 ( .A(n186), .B(n4398), .Z(n4397) );
  XNOR U4268 ( .A(n4399), .B(n4396), .Z(n4398) );
  XOR U4269 ( .A(n4400), .B(n4401), .Z(n186) );
  AND U4270 ( .A(n4402), .B(n4403), .Z(n4401) );
  XNOR U4271 ( .A(n4223), .B(n4400), .Z(n4403) );
  AND U4272 ( .A(p_input[511]), .B(p_input[495]), .Z(n4223) );
  XOR U4273 ( .A(n4400), .B(n4224), .Z(n4402) );
  AND U4274 ( .A(p_input[479]), .B(p_input[463]), .Z(n4224) );
  XOR U4275 ( .A(n4404), .B(n4405), .Z(n4400) );
  AND U4276 ( .A(n4406), .B(n4407), .Z(n4405) );
  XOR U4277 ( .A(n4404), .B(n4234), .Z(n4407) );
  XNOR U4278 ( .A(p_input[494]), .B(n4408), .Z(n4234) );
  AND U4279 ( .A(n218), .B(n4409), .Z(n4408) );
  XOR U4280 ( .A(p_input[510]), .B(p_input[494]), .Z(n4409) );
  XNOR U4281 ( .A(n4231), .B(n4404), .Z(n4406) );
  XOR U4282 ( .A(n4410), .B(n4411), .Z(n4231) );
  AND U4283 ( .A(n216), .B(n4412), .Z(n4411) );
  XOR U4284 ( .A(p_input[478]), .B(p_input[462]), .Z(n4412) );
  XOR U4285 ( .A(n4413), .B(n4414), .Z(n4404) );
  AND U4286 ( .A(n4415), .B(n4416), .Z(n4414) );
  XOR U4287 ( .A(n4413), .B(n4246), .Z(n4416) );
  XNOR U4288 ( .A(p_input[493]), .B(n4417), .Z(n4246) );
  AND U4289 ( .A(n218), .B(n4418), .Z(n4417) );
  XOR U4290 ( .A(p_input[509]), .B(p_input[493]), .Z(n4418) );
  XNOR U4291 ( .A(n4243), .B(n4413), .Z(n4415) );
  XOR U4292 ( .A(n4419), .B(n4420), .Z(n4243) );
  AND U4293 ( .A(n216), .B(n4421), .Z(n4420) );
  XOR U4294 ( .A(p_input[477]), .B(p_input[461]), .Z(n4421) );
  XOR U4295 ( .A(n4422), .B(n4423), .Z(n4413) );
  AND U4296 ( .A(n4424), .B(n4425), .Z(n4423) );
  XOR U4297 ( .A(n4422), .B(n4258), .Z(n4425) );
  XNOR U4298 ( .A(p_input[492]), .B(n4426), .Z(n4258) );
  AND U4299 ( .A(n218), .B(n4427), .Z(n4426) );
  XOR U4300 ( .A(p_input[508]), .B(p_input[492]), .Z(n4427) );
  XNOR U4301 ( .A(n4255), .B(n4422), .Z(n4424) );
  XOR U4302 ( .A(n4428), .B(n4429), .Z(n4255) );
  AND U4303 ( .A(n216), .B(n4430), .Z(n4429) );
  XOR U4304 ( .A(p_input[476]), .B(p_input[460]), .Z(n4430) );
  XOR U4305 ( .A(n4431), .B(n4432), .Z(n4422) );
  AND U4306 ( .A(n4433), .B(n4434), .Z(n4432) );
  XOR U4307 ( .A(n4431), .B(n4270), .Z(n4434) );
  XNOR U4308 ( .A(p_input[491]), .B(n4435), .Z(n4270) );
  AND U4309 ( .A(n218), .B(n4436), .Z(n4435) );
  XOR U4310 ( .A(p_input[507]), .B(p_input[491]), .Z(n4436) );
  XNOR U4311 ( .A(n4267), .B(n4431), .Z(n4433) );
  XOR U4312 ( .A(n4437), .B(n4438), .Z(n4267) );
  AND U4313 ( .A(n216), .B(n4439), .Z(n4438) );
  XOR U4314 ( .A(p_input[475]), .B(p_input[459]), .Z(n4439) );
  XOR U4315 ( .A(n4440), .B(n4441), .Z(n4431) );
  AND U4316 ( .A(n4442), .B(n4443), .Z(n4441) );
  XOR U4317 ( .A(n4440), .B(n4282), .Z(n4443) );
  XNOR U4318 ( .A(p_input[490]), .B(n4444), .Z(n4282) );
  AND U4319 ( .A(n218), .B(n4445), .Z(n4444) );
  XOR U4320 ( .A(p_input[506]), .B(p_input[490]), .Z(n4445) );
  XNOR U4321 ( .A(n4279), .B(n4440), .Z(n4442) );
  XOR U4322 ( .A(n4446), .B(n4447), .Z(n4279) );
  AND U4323 ( .A(n216), .B(n4448), .Z(n4447) );
  XOR U4324 ( .A(p_input[474]), .B(p_input[458]), .Z(n4448) );
  XOR U4325 ( .A(n4449), .B(n4450), .Z(n4440) );
  AND U4326 ( .A(n4451), .B(n4452), .Z(n4450) );
  XOR U4327 ( .A(n4449), .B(n4294), .Z(n4452) );
  XNOR U4328 ( .A(p_input[489]), .B(n4453), .Z(n4294) );
  AND U4329 ( .A(n218), .B(n4454), .Z(n4453) );
  XOR U4330 ( .A(p_input[505]), .B(p_input[489]), .Z(n4454) );
  XNOR U4331 ( .A(n4291), .B(n4449), .Z(n4451) );
  XOR U4332 ( .A(n4455), .B(n4456), .Z(n4291) );
  AND U4333 ( .A(n216), .B(n4457), .Z(n4456) );
  XOR U4334 ( .A(p_input[473]), .B(p_input[457]), .Z(n4457) );
  XOR U4335 ( .A(n4458), .B(n4459), .Z(n4449) );
  AND U4336 ( .A(n4460), .B(n4461), .Z(n4459) );
  XOR U4337 ( .A(n4458), .B(n4306), .Z(n4461) );
  XNOR U4338 ( .A(p_input[488]), .B(n4462), .Z(n4306) );
  AND U4339 ( .A(n218), .B(n4463), .Z(n4462) );
  XOR U4340 ( .A(p_input[504]), .B(p_input[488]), .Z(n4463) );
  XNOR U4341 ( .A(n4303), .B(n4458), .Z(n4460) );
  XOR U4342 ( .A(n4464), .B(n4465), .Z(n4303) );
  AND U4343 ( .A(n216), .B(n4466), .Z(n4465) );
  XOR U4344 ( .A(p_input[472]), .B(p_input[456]), .Z(n4466) );
  XOR U4345 ( .A(n4467), .B(n4468), .Z(n4458) );
  AND U4346 ( .A(n4469), .B(n4470), .Z(n4468) );
  XOR U4347 ( .A(n4467), .B(n4318), .Z(n4470) );
  XNOR U4348 ( .A(p_input[487]), .B(n4471), .Z(n4318) );
  AND U4349 ( .A(n218), .B(n4472), .Z(n4471) );
  XOR U4350 ( .A(p_input[503]), .B(p_input[487]), .Z(n4472) );
  XNOR U4351 ( .A(n4315), .B(n4467), .Z(n4469) );
  XOR U4352 ( .A(n4473), .B(n4474), .Z(n4315) );
  AND U4353 ( .A(n216), .B(n4475), .Z(n4474) );
  XOR U4354 ( .A(p_input[471]), .B(p_input[455]), .Z(n4475) );
  XOR U4355 ( .A(n4476), .B(n4477), .Z(n4467) );
  AND U4356 ( .A(n4478), .B(n4479), .Z(n4477) );
  XOR U4357 ( .A(n4476), .B(n4330), .Z(n4479) );
  XNOR U4358 ( .A(p_input[486]), .B(n4480), .Z(n4330) );
  AND U4359 ( .A(n218), .B(n4481), .Z(n4480) );
  XOR U4360 ( .A(p_input[502]), .B(p_input[486]), .Z(n4481) );
  XNOR U4361 ( .A(n4327), .B(n4476), .Z(n4478) );
  XOR U4362 ( .A(n4482), .B(n4483), .Z(n4327) );
  AND U4363 ( .A(n216), .B(n4484), .Z(n4483) );
  XOR U4364 ( .A(p_input[470]), .B(p_input[454]), .Z(n4484) );
  XOR U4365 ( .A(n4485), .B(n4486), .Z(n4476) );
  AND U4366 ( .A(n4487), .B(n4488), .Z(n4486) );
  XOR U4367 ( .A(n4485), .B(n4342), .Z(n4488) );
  XNOR U4368 ( .A(p_input[485]), .B(n4489), .Z(n4342) );
  AND U4369 ( .A(n218), .B(n4490), .Z(n4489) );
  XOR U4370 ( .A(p_input[501]), .B(p_input[485]), .Z(n4490) );
  XNOR U4371 ( .A(n4339), .B(n4485), .Z(n4487) );
  XOR U4372 ( .A(n4491), .B(n4492), .Z(n4339) );
  AND U4373 ( .A(n216), .B(n4493), .Z(n4492) );
  XOR U4374 ( .A(p_input[469]), .B(p_input[453]), .Z(n4493) );
  XOR U4375 ( .A(n4494), .B(n4495), .Z(n4485) );
  AND U4376 ( .A(n4496), .B(n4497), .Z(n4495) );
  XOR U4377 ( .A(n4494), .B(n4354), .Z(n4497) );
  XNOR U4378 ( .A(p_input[484]), .B(n4498), .Z(n4354) );
  AND U4379 ( .A(n218), .B(n4499), .Z(n4498) );
  XOR U4380 ( .A(p_input[500]), .B(p_input[484]), .Z(n4499) );
  XNOR U4381 ( .A(n4351), .B(n4494), .Z(n4496) );
  XOR U4382 ( .A(n4500), .B(n4501), .Z(n4351) );
  AND U4383 ( .A(n216), .B(n4502), .Z(n4501) );
  XOR U4384 ( .A(p_input[468]), .B(p_input[452]), .Z(n4502) );
  XOR U4385 ( .A(n4503), .B(n4504), .Z(n4494) );
  AND U4386 ( .A(n4505), .B(n4506), .Z(n4504) );
  XOR U4387 ( .A(n4366), .B(n4503), .Z(n4506) );
  XNOR U4388 ( .A(p_input[483]), .B(n4507), .Z(n4366) );
  AND U4389 ( .A(n218), .B(n4508), .Z(n4507) );
  XOR U4390 ( .A(p_input[499]), .B(p_input[483]), .Z(n4508) );
  XNOR U4391 ( .A(n4503), .B(n4363), .Z(n4505) );
  XOR U4392 ( .A(n4509), .B(n4510), .Z(n4363) );
  AND U4393 ( .A(n216), .B(n4511), .Z(n4510) );
  XOR U4394 ( .A(p_input[467]), .B(p_input[451]), .Z(n4511) );
  XOR U4395 ( .A(n4512), .B(n4513), .Z(n4503) );
  AND U4396 ( .A(n4514), .B(n4515), .Z(n4513) );
  XOR U4397 ( .A(n4512), .B(n4378), .Z(n4515) );
  XNOR U4398 ( .A(p_input[482]), .B(n4516), .Z(n4378) );
  AND U4399 ( .A(n218), .B(n4517), .Z(n4516) );
  XOR U4400 ( .A(p_input[498]), .B(p_input[482]), .Z(n4517) );
  XNOR U4401 ( .A(n4375), .B(n4512), .Z(n4514) );
  XOR U4402 ( .A(n4518), .B(n4519), .Z(n4375) );
  AND U4403 ( .A(n216), .B(n4520), .Z(n4519) );
  XOR U4404 ( .A(p_input[466]), .B(p_input[450]), .Z(n4520) );
  XOR U4405 ( .A(n4521), .B(n4522), .Z(n4512) );
  AND U4406 ( .A(n4523), .B(n4524), .Z(n4522) );
  XNOR U4407 ( .A(n4525), .B(n4391), .Z(n4524) );
  XNOR U4408 ( .A(p_input[481]), .B(n4526), .Z(n4391) );
  AND U4409 ( .A(n218), .B(n4527), .Z(n4526) );
  XNOR U4410 ( .A(p_input[497]), .B(n4528), .Z(n4527) );
  IV U4411 ( .A(p_input[481]), .Z(n4528) );
  XNOR U4412 ( .A(n4388), .B(n4521), .Z(n4523) );
  XNOR U4413 ( .A(p_input[449]), .B(n4529), .Z(n4388) );
  AND U4414 ( .A(n216), .B(n4530), .Z(n4529) );
  XOR U4415 ( .A(p_input[465]), .B(p_input[449]), .Z(n4530) );
  IV U4416 ( .A(n4525), .Z(n4521) );
  AND U4417 ( .A(n4396), .B(n4399), .Z(n4525) );
  XOR U4418 ( .A(p_input[480]), .B(n4531), .Z(n4399) );
  AND U4419 ( .A(n218), .B(n4532), .Z(n4531) );
  XOR U4420 ( .A(p_input[496]), .B(p_input[480]), .Z(n4532) );
  XOR U4421 ( .A(n4533), .B(n4534), .Z(n218) );
  AND U4422 ( .A(n4535), .B(n4536), .Z(n4534) );
  XNOR U4423 ( .A(p_input[511]), .B(n4533), .Z(n4536) );
  XOR U4424 ( .A(n4533), .B(p_input[495]), .Z(n4535) );
  XOR U4425 ( .A(n4537), .B(n4538), .Z(n4533) );
  AND U4426 ( .A(n4539), .B(n4540), .Z(n4538) );
  XNOR U4427 ( .A(p_input[510]), .B(n4537), .Z(n4540) );
  XOR U4428 ( .A(n4537), .B(p_input[494]), .Z(n4539) );
  XOR U4429 ( .A(n4541), .B(n4542), .Z(n4537) );
  AND U4430 ( .A(n4543), .B(n4544), .Z(n4542) );
  XNOR U4431 ( .A(p_input[509]), .B(n4541), .Z(n4544) );
  XOR U4432 ( .A(n4541), .B(p_input[493]), .Z(n4543) );
  XOR U4433 ( .A(n4545), .B(n4546), .Z(n4541) );
  AND U4434 ( .A(n4547), .B(n4548), .Z(n4546) );
  XNOR U4435 ( .A(p_input[508]), .B(n4545), .Z(n4548) );
  XOR U4436 ( .A(n4545), .B(p_input[492]), .Z(n4547) );
  XOR U4437 ( .A(n4549), .B(n4550), .Z(n4545) );
  AND U4438 ( .A(n4551), .B(n4552), .Z(n4550) );
  XNOR U4439 ( .A(p_input[507]), .B(n4549), .Z(n4552) );
  XOR U4440 ( .A(n4549), .B(p_input[491]), .Z(n4551) );
  XOR U4441 ( .A(n4553), .B(n4554), .Z(n4549) );
  AND U4442 ( .A(n4555), .B(n4556), .Z(n4554) );
  XNOR U4443 ( .A(p_input[506]), .B(n4553), .Z(n4556) );
  XOR U4444 ( .A(n4553), .B(p_input[490]), .Z(n4555) );
  XOR U4445 ( .A(n4557), .B(n4558), .Z(n4553) );
  AND U4446 ( .A(n4559), .B(n4560), .Z(n4558) );
  XNOR U4447 ( .A(p_input[505]), .B(n4557), .Z(n4560) );
  XOR U4448 ( .A(n4557), .B(p_input[489]), .Z(n4559) );
  XOR U4449 ( .A(n4561), .B(n4562), .Z(n4557) );
  AND U4450 ( .A(n4563), .B(n4564), .Z(n4562) );
  XNOR U4451 ( .A(p_input[504]), .B(n4561), .Z(n4564) );
  XOR U4452 ( .A(n4561), .B(p_input[488]), .Z(n4563) );
  XOR U4453 ( .A(n4565), .B(n4566), .Z(n4561) );
  AND U4454 ( .A(n4567), .B(n4568), .Z(n4566) );
  XNOR U4455 ( .A(p_input[503]), .B(n4565), .Z(n4568) );
  XOR U4456 ( .A(n4565), .B(p_input[487]), .Z(n4567) );
  XOR U4457 ( .A(n4569), .B(n4570), .Z(n4565) );
  AND U4458 ( .A(n4571), .B(n4572), .Z(n4570) );
  XNOR U4459 ( .A(p_input[502]), .B(n4569), .Z(n4572) );
  XOR U4460 ( .A(n4569), .B(p_input[486]), .Z(n4571) );
  XOR U4461 ( .A(n4573), .B(n4574), .Z(n4569) );
  AND U4462 ( .A(n4575), .B(n4576), .Z(n4574) );
  XNOR U4463 ( .A(p_input[501]), .B(n4573), .Z(n4576) );
  XOR U4464 ( .A(n4573), .B(p_input[485]), .Z(n4575) );
  XOR U4465 ( .A(n4577), .B(n4578), .Z(n4573) );
  AND U4466 ( .A(n4579), .B(n4580), .Z(n4578) );
  XNOR U4467 ( .A(p_input[500]), .B(n4577), .Z(n4580) );
  XOR U4468 ( .A(n4577), .B(p_input[484]), .Z(n4579) );
  XOR U4469 ( .A(n4581), .B(n4582), .Z(n4577) );
  AND U4470 ( .A(n4583), .B(n4584), .Z(n4582) );
  XNOR U4471 ( .A(p_input[499]), .B(n4581), .Z(n4584) );
  XOR U4472 ( .A(n4581), .B(p_input[483]), .Z(n4583) );
  XOR U4473 ( .A(n4585), .B(n4586), .Z(n4581) );
  AND U4474 ( .A(n4587), .B(n4588), .Z(n4586) );
  XNOR U4475 ( .A(p_input[498]), .B(n4585), .Z(n4588) );
  XOR U4476 ( .A(n4585), .B(p_input[482]), .Z(n4587) );
  XNOR U4477 ( .A(n4589), .B(n4590), .Z(n4585) );
  AND U4478 ( .A(n4591), .B(n4592), .Z(n4590) );
  XOR U4479 ( .A(p_input[497]), .B(n4589), .Z(n4592) );
  XNOR U4480 ( .A(p_input[481]), .B(n4589), .Z(n4591) );
  AND U4481 ( .A(p_input[496]), .B(n4593), .Z(n4589) );
  IV U4482 ( .A(p_input[480]), .Z(n4593) );
  XNOR U4483 ( .A(p_input[448]), .B(n4594), .Z(n4396) );
  AND U4484 ( .A(n216), .B(n4595), .Z(n4594) );
  XOR U4485 ( .A(p_input[464]), .B(p_input[448]), .Z(n4595) );
  XOR U4486 ( .A(n4596), .B(n4597), .Z(n216) );
  AND U4487 ( .A(n4598), .B(n4599), .Z(n4597) );
  XNOR U4488 ( .A(p_input[479]), .B(n4596), .Z(n4599) );
  XOR U4489 ( .A(n4596), .B(p_input[463]), .Z(n4598) );
  XOR U4490 ( .A(n4600), .B(n4601), .Z(n4596) );
  AND U4491 ( .A(n4602), .B(n4603), .Z(n4601) );
  XNOR U4492 ( .A(p_input[478]), .B(n4600), .Z(n4603) );
  XNOR U4493 ( .A(n4600), .B(n4410), .Z(n4602) );
  IV U4494 ( .A(p_input[462]), .Z(n4410) );
  XOR U4495 ( .A(n4604), .B(n4605), .Z(n4600) );
  AND U4496 ( .A(n4606), .B(n4607), .Z(n4605) );
  XNOR U4497 ( .A(p_input[477]), .B(n4604), .Z(n4607) );
  XNOR U4498 ( .A(n4604), .B(n4419), .Z(n4606) );
  IV U4499 ( .A(p_input[461]), .Z(n4419) );
  XOR U4500 ( .A(n4608), .B(n4609), .Z(n4604) );
  AND U4501 ( .A(n4610), .B(n4611), .Z(n4609) );
  XNOR U4502 ( .A(p_input[476]), .B(n4608), .Z(n4611) );
  XNOR U4503 ( .A(n4608), .B(n4428), .Z(n4610) );
  IV U4504 ( .A(p_input[460]), .Z(n4428) );
  XOR U4505 ( .A(n4612), .B(n4613), .Z(n4608) );
  AND U4506 ( .A(n4614), .B(n4615), .Z(n4613) );
  XNOR U4507 ( .A(p_input[475]), .B(n4612), .Z(n4615) );
  XNOR U4508 ( .A(n4612), .B(n4437), .Z(n4614) );
  IV U4509 ( .A(p_input[459]), .Z(n4437) );
  XOR U4510 ( .A(n4616), .B(n4617), .Z(n4612) );
  AND U4511 ( .A(n4618), .B(n4619), .Z(n4617) );
  XNOR U4512 ( .A(p_input[474]), .B(n4616), .Z(n4619) );
  XNOR U4513 ( .A(n4616), .B(n4446), .Z(n4618) );
  IV U4514 ( .A(p_input[458]), .Z(n4446) );
  XOR U4515 ( .A(n4620), .B(n4621), .Z(n4616) );
  AND U4516 ( .A(n4622), .B(n4623), .Z(n4621) );
  XNOR U4517 ( .A(p_input[473]), .B(n4620), .Z(n4623) );
  XNOR U4518 ( .A(n4620), .B(n4455), .Z(n4622) );
  IV U4519 ( .A(p_input[457]), .Z(n4455) );
  XOR U4520 ( .A(n4624), .B(n4625), .Z(n4620) );
  AND U4521 ( .A(n4626), .B(n4627), .Z(n4625) );
  XNOR U4522 ( .A(p_input[472]), .B(n4624), .Z(n4627) );
  XNOR U4523 ( .A(n4624), .B(n4464), .Z(n4626) );
  IV U4524 ( .A(p_input[456]), .Z(n4464) );
  XOR U4525 ( .A(n4628), .B(n4629), .Z(n4624) );
  AND U4526 ( .A(n4630), .B(n4631), .Z(n4629) );
  XNOR U4527 ( .A(p_input[471]), .B(n4628), .Z(n4631) );
  XNOR U4528 ( .A(n4628), .B(n4473), .Z(n4630) );
  IV U4529 ( .A(p_input[455]), .Z(n4473) );
  XOR U4530 ( .A(n4632), .B(n4633), .Z(n4628) );
  AND U4531 ( .A(n4634), .B(n4635), .Z(n4633) );
  XNOR U4532 ( .A(p_input[470]), .B(n4632), .Z(n4635) );
  XNOR U4533 ( .A(n4632), .B(n4482), .Z(n4634) );
  IV U4534 ( .A(p_input[454]), .Z(n4482) );
  XOR U4535 ( .A(n4636), .B(n4637), .Z(n4632) );
  AND U4536 ( .A(n4638), .B(n4639), .Z(n4637) );
  XNOR U4537 ( .A(p_input[469]), .B(n4636), .Z(n4639) );
  XNOR U4538 ( .A(n4636), .B(n4491), .Z(n4638) );
  IV U4539 ( .A(p_input[453]), .Z(n4491) );
  XOR U4540 ( .A(n4640), .B(n4641), .Z(n4636) );
  AND U4541 ( .A(n4642), .B(n4643), .Z(n4641) );
  XNOR U4542 ( .A(p_input[468]), .B(n4640), .Z(n4643) );
  XNOR U4543 ( .A(n4640), .B(n4500), .Z(n4642) );
  IV U4544 ( .A(p_input[452]), .Z(n4500) );
  XOR U4545 ( .A(n4644), .B(n4645), .Z(n4640) );
  AND U4546 ( .A(n4646), .B(n4647), .Z(n4645) );
  XNOR U4547 ( .A(p_input[467]), .B(n4644), .Z(n4647) );
  XNOR U4548 ( .A(n4644), .B(n4509), .Z(n4646) );
  IV U4549 ( .A(p_input[451]), .Z(n4509) );
  XOR U4550 ( .A(n4648), .B(n4649), .Z(n4644) );
  AND U4551 ( .A(n4650), .B(n4651), .Z(n4649) );
  XNOR U4552 ( .A(p_input[466]), .B(n4648), .Z(n4651) );
  XNOR U4553 ( .A(n4648), .B(n4518), .Z(n4650) );
  IV U4554 ( .A(p_input[450]), .Z(n4518) );
  XNOR U4555 ( .A(n4652), .B(n4653), .Z(n4648) );
  AND U4556 ( .A(n4654), .B(n4655), .Z(n4653) );
  XOR U4557 ( .A(p_input[465]), .B(n4652), .Z(n4655) );
  XNOR U4558 ( .A(p_input[449]), .B(n4652), .Z(n4654) );
  AND U4559 ( .A(p_input[464]), .B(n4656), .Z(n4652) );
  IV U4560 ( .A(p_input[448]), .Z(n4656) );
  XOR U4561 ( .A(n4657), .B(n4658), .Z(n4215) );
  AND U4562 ( .A(n184), .B(n4659), .Z(n4658) );
  XNOR U4563 ( .A(n4660), .B(n4657), .Z(n4659) );
  XOR U4564 ( .A(n4661), .B(n4662), .Z(n184) );
  AND U4565 ( .A(n4663), .B(n4664), .Z(n4662) );
  XNOR U4566 ( .A(n4225), .B(n4661), .Z(n4664) );
  AND U4567 ( .A(p_input[447]), .B(p_input[431]), .Z(n4225) );
  XOR U4568 ( .A(n4661), .B(n4226), .Z(n4663) );
  AND U4569 ( .A(p_input[415]), .B(p_input[399]), .Z(n4226) );
  XOR U4570 ( .A(n4665), .B(n4666), .Z(n4661) );
  AND U4571 ( .A(n4667), .B(n4668), .Z(n4666) );
  XOR U4572 ( .A(n4665), .B(n4238), .Z(n4668) );
  XNOR U4573 ( .A(p_input[430]), .B(n4669), .Z(n4238) );
  AND U4574 ( .A(n222), .B(n4670), .Z(n4669) );
  XOR U4575 ( .A(p_input[446]), .B(p_input[430]), .Z(n4670) );
  XNOR U4576 ( .A(n4235), .B(n4665), .Z(n4667) );
  XOR U4577 ( .A(n4671), .B(n4672), .Z(n4235) );
  AND U4578 ( .A(n219), .B(n4673), .Z(n4672) );
  XOR U4579 ( .A(p_input[414]), .B(p_input[398]), .Z(n4673) );
  XOR U4580 ( .A(n4674), .B(n4675), .Z(n4665) );
  AND U4581 ( .A(n4676), .B(n4677), .Z(n4675) );
  XOR U4582 ( .A(n4674), .B(n4250), .Z(n4677) );
  XNOR U4583 ( .A(p_input[429]), .B(n4678), .Z(n4250) );
  AND U4584 ( .A(n222), .B(n4679), .Z(n4678) );
  XOR U4585 ( .A(p_input[445]), .B(p_input[429]), .Z(n4679) );
  XNOR U4586 ( .A(n4247), .B(n4674), .Z(n4676) );
  XOR U4587 ( .A(n4680), .B(n4681), .Z(n4247) );
  AND U4588 ( .A(n219), .B(n4682), .Z(n4681) );
  XOR U4589 ( .A(p_input[413]), .B(p_input[397]), .Z(n4682) );
  XOR U4590 ( .A(n4683), .B(n4684), .Z(n4674) );
  AND U4591 ( .A(n4685), .B(n4686), .Z(n4684) );
  XOR U4592 ( .A(n4683), .B(n4262), .Z(n4686) );
  XNOR U4593 ( .A(p_input[428]), .B(n4687), .Z(n4262) );
  AND U4594 ( .A(n222), .B(n4688), .Z(n4687) );
  XOR U4595 ( .A(p_input[444]), .B(p_input[428]), .Z(n4688) );
  XNOR U4596 ( .A(n4259), .B(n4683), .Z(n4685) );
  XOR U4597 ( .A(n4689), .B(n4690), .Z(n4259) );
  AND U4598 ( .A(n219), .B(n4691), .Z(n4690) );
  XOR U4599 ( .A(p_input[412]), .B(p_input[396]), .Z(n4691) );
  XOR U4600 ( .A(n4692), .B(n4693), .Z(n4683) );
  AND U4601 ( .A(n4694), .B(n4695), .Z(n4693) );
  XOR U4602 ( .A(n4692), .B(n4274), .Z(n4695) );
  XNOR U4603 ( .A(p_input[427]), .B(n4696), .Z(n4274) );
  AND U4604 ( .A(n222), .B(n4697), .Z(n4696) );
  XOR U4605 ( .A(p_input[443]), .B(p_input[427]), .Z(n4697) );
  XNOR U4606 ( .A(n4271), .B(n4692), .Z(n4694) );
  XOR U4607 ( .A(n4698), .B(n4699), .Z(n4271) );
  AND U4608 ( .A(n219), .B(n4700), .Z(n4699) );
  XOR U4609 ( .A(p_input[411]), .B(p_input[395]), .Z(n4700) );
  XOR U4610 ( .A(n4701), .B(n4702), .Z(n4692) );
  AND U4611 ( .A(n4703), .B(n4704), .Z(n4702) );
  XOR U4612 ( .A(n4701), .B(n4286), .Z(n4704) );
  XNOR U4613 ( .A(p_input[426]), .B(n4705), .Z(n4286) );
  AND U4614 ( .A(n222), .B(n4706), .Z(n4705) );
  XOR U4615 ( .A(p_input[442]), .B(p_input[426]), .Z(n4706) );
  XNOR U4616 ( .A(n4283), .B(n4701), .Z(n4703) );
  XOR U4617 ( .A(n4707), .B(n4708), .Z(n4283) );
  AND U4618 ( .A(n219), .B(n4709), .Z(n4708) );
  XOR U4619 ( .A(p_input[410]), .B(p_input[394]), .Z(n4709) );
  XOR U4620 ( .A(n4710), .B(n4711), .Z(n4701) );
  AND U4621 ( .A(n4712), .B(n4713), .Z(n4711) );
  XOR U4622 ( .A(n4710), .B(n4298), .Z(n4713) );
  XNOR U4623 ( .A(p_input[425]), .B(n4714), .Z(n4298) );
  AND U4624 ( .A(n222), .B(n4715), .Z(n4714) );
  XOR U4625 ( .A(p_input[441]), .B(p_input[425]), .Z(n4715) );
  XNOR U4626 ( .A(n4295), .B(n4710), .Z(n4712) );
  XOR U4627 ( .A(n4716), .B(n4717), .Z(n4295) );
  AND U4628 ( .A(n219), .B(n4718), .Z(n4717) );
  XOR U4629 ( .A(p_input[409]), .B(p_input[393]), .Z(n4718) );
  XOR U4630 ( .A(n4719), .B(n4720), .Z(n4710) );
  AND U4631 ( .A(n4721), .B(n4722), .Z(n4720) );
  XOR U4632 ( .A(n4719), .B(n4310), .Z(n4722) );
  XNOR U4633 ( .A(p_input[424]), .B(n4723), .Z(n4310) );
  AND U4634 ( .A(n222), .B(n4724), .Z(n4723) );
  XOR U4635 ( .A(p_input[440]), .B(p_input[424]), .Z(n4724) );
  XNOR U4636 ( .A(n4307), .B(n4719), .Z(n4721) );
  XOR U4637 ( .A(n4725), .B(n4726), .Z(n4307) );
  AND U4638 ( .A(n219), .B(n4727), .Z(n4726) );
  XOR U4639 ( .A(p_input[408]), .B(p_input[392]), .Z(n4727) );
  XOR U4640 ( .A(n4728), .B(n4729), .Z(n4719) );
  AND U4641 ( .A(n4730), .B(n4731), .Z(n4729) );
  XOR U4642 ( .A(n4728), .B(n4322), .Z(n4731) );
  XNOR U4643 ( .A(p_input[423]), .B(n4732), .Z(n4322) );
  AND U4644 ( .A(n222), .B(n4733), .Z(n4732) );
  XOR U4645 ( .A(p_input[439]), .B(p_input[423]), .Z(n4733) );
  XNOR U4646 ( .A(n4319), .B(n4728), .Z(n4730) );
  XOR U4647 ( .A(n4734), .B(n4735), .Z(n4319) );
  AND U4648 ( .A(n219), .B(n4736), .Z(n4735) );
  XOR U4649 ( .A(p_input[407]), .B(p_input[391]), .Z(n4736) );
  XOR U4650 ( .A(n4737), .B(n4738), .Z(n4728) );
  AND U4651 ( .A(n4739), .B(n4740), .Z(n4738) );
  XOR U4652 ( .A(n4737), .B(n4334), .Z(n4740) );
  XNOR U4653 ( .A(p_input[422]), .B(n4741), .Z(n4334) );
  AND U4654 ( .A(n222), .B(n4742), .Z(n4741) );
  XOR U4655 ( .A(p_input[438]), .B(p_input[422]), .Z(n4742) );
  XNOR U4656 ( .A(n4331), .B(n4737), .Z(n4739) );
  XOR U4657 ( .A(n4743), .B(n4744), .Z(n4331) );
  AND U4658 ( .A(n219), .B(n4745), .Z(n4744) );
  XOR U4659 ( .A(p_input[406]), .B(p_input[390]), .Z(n4745) );
  XOR U4660 ( .A(n4746), .B(n4747), .Z(n4737) );
  AND U4661 ( .A(n4748), .B(n4749), .Z(n4747) );
  XOR U4662 ( .A(n4746), .B(n4346), .Z(n4749) );
  XNOR U4663 ( .A(p_input[421]), .B(n4750), .Z(n4346) );
  AND U4664 ( .A(n222), .B(n4751), .Z(n4750) );
  XOR U4665 ( .A(p_input[437]), .B(p_input[421]), .Z(n4751) );
  XNOR U4666 ( .A(n4343), .B(n4746), .Z(n4748) );
  XOR U4667 ( .A(n4752), .B(n4753), .Z(n4343) );
  AND U4668 ( .A(n219), .B(n4754), .Z(n4753) );
  XOR U4669 ( .A(p_input[405]), .B(p_input[389]), .Z(n4754) );
  XOR U4670 ( .A(n4755), .B(n4756), .Z(n4746) );
  AND U4671 ( .A(n4757), .B(n4758), .Z(n4756) );
  XOR U4672 ( .A(n4755), .B(n4358), .Z(n4758) );
  XNOR U4673 ( .A(p_input[420]), .B(n4759), .Z(n4358) );
  AND U4674 ( .A(n222), .B(n4760), .Z(n4759) );
  XOR U4675 ( .A(p_input[436]), .B(p_input[420]), .Z(n4760) );
  XNOR U4676 ( .A(n4355), .B(n4755), .Z(n4757) );
  XOR U4677 ( .A(n4761), .B(n4762), .Z(n4355) );
  AND U4678 ( .A(n219), .B(n4763), .Z(n4762) );
  XOR U4679 ( .A(p_input[404]), .B(p_input[388]), .Z(n4763) );
  XOR U4680 ( .A(n4764), .B(n4765), .Z(n4755) );
  AND U4681 ( .A(n4766), .B(n4767), .Z(n4765) );
  XOR U4682 ( .A(n4370), .B(n4764), .Z(n4767) );
  XNOR U4683 ( .A(p_input[419]), .B(n4768), .Z(n4370) );
  AND U4684 ( .A(n222), .B(n4769), .Z(n4768) );
  XOR U4685 ( .A(p_input[435]), .B(p_input[419]), .Z(n4769) );
  XNOR U4686 ( .A(n4764), .B(n4367), .Z(n4766) );
  XOR U4687 ( .A(n4770), .B(n4771), .Z(n4367) );
  AND U4688 ( .A(n219), .B(n4772), .Z(n4771) );
  XOR U4689 ( .A(p_input[403]), .B(p_input[387]), .Z(n4772) );
  XOR U4690 ( .A(n4773), .B(n4774), .Z(n4764) );
  AND U4691 ( .A(n4775), .B(n4776), .Z(n4774) );
  XOR U4692 ( .A(n4773), .B(n4382), .Z(n4776) );
  XNOR U4693 ( .A(p_input[418]), .B(n4777), .Z(n4382) );
  AND U4694 ( .A(n222), .B(n4778), .Z(n4777) );
  XOR U4695 ( .A(p_input[434]), .B(p_input[418]), .Z(n4778) );
  XNOR U4696 ( .A(n4379), .B(n4773), .Z(n4775) );
  XOR U4697 ( .A(n4779), .B(n4780), .Z(n4379) );
  AND U4698 ( .A(n219), .B(n4781), .Z(n4780) );
  XOR U4699 ( .A(p_input[402]), .B(p_input[386]), .Z(n4781) );
  XOR U4700 ( .A(n4782), .B(n4783), .Z(n4773) );
  AND U4701 ( .A(n4784), .B(n4785), .Z(n4783) );
  XNOR U4702 ( .A(n4786), .B(n4395), .Z(n4785) );
  XNOR U4703 ( .A(p_input[417]), .B(n4787), .Z(n4395) );
  AND U4704 ( .A(n222), .B(n4788), .Z(n4787) );
  XNOR U4705 ( .A(p_input[433]), .B(n4789), .Z(n4788) );
  IV U4706 ( .A(p_input[417]), .Z(n4789) );
  XNOR U4707 ( .A(n4392), .B(n4782), .Z(n4784) );
  XNOR U4708 ( .A(p_input[385]), .B(n4790), .Z(n4392) );
  AND U4709 ( .A(n219), .B(n4791), .Z(n4790) );
  XOR U4710 ( .A(p_input[401]), .B(p_input[385]), .Z(n4791) );
  IV U4711 ( .A(n4786), .Z(n4782) );
  AND U4712 ( .A(n4657), .B(n4660), .Z(n4786) );
  XOR U4713 ( .A(p_input[416]), .B(n4792), .Z(n4660) );
  AND U4714 ( .A(n222), .B(n4793), .Z(n4792) );
  XOR U4715 ( .A(p_input[432]), .B(p_input[416]), .Z(n4793) );
  XOR U4716 ( .A(n4794), .B(n4795), .Z(n222) );
  AND U4717 ( .A(n4796), .B(n4797), .Z(n4795) );
  XNOR U4718 ( .A(p_input[447]), .B(n4794), .Z(n4797) );
  XOR U4719 ( .A(n4794), .B(p_input[431]), .Z(n4796) );
  XOR U4720 ( .A(n4798), .B(n4799), .Z(n4794) );
  AND U4721 ( .A(n4800), .B(n4801), .Z(n4799) );
  XNOR U4722 ( .A(p_input[446]), .B(n4798), .Z(n4801) );
  XOR U4723 ( .A(n4798), .B(p_input[430]), .Z(n4800) );
  XOR U4724 ( .A(n4802), .B(n4803), .Z(n4798) );
  AND U4725 ( .A(n4804), .B(n4805), .Z(n4803) );
  XNOR U4726 ( .A(p_input[445]), .B(n4802), .Z(n4805) );
  XOR U4727 ( .A(n4802), .B(p_input[429]), .Z(n4804) );
  XOR U4728 ( .A(n4806), .B(n4807), .Z(n4802) );
  AND U4729 ( .A(n4808), .B(n4809), .Z(n4807) );
  XNOR U4730 ( .A(p_input[444]), .B(n4806), .Z(n4809) );
  XOR U4731 ( .A(n4806), .B(p_input[428]), .Z(n4808) );
  XOR U4732 ( .A(n4810), .B(n4811), .Z(n4806) );
  AND U4733 ( .A(n4812), .B(n4813), .Z(n4811) );
  XNOR U4734 ( .A(p_input[443]), .B(n4810), .Z(n4813) );
  XOR U4735 ( .A(n4810), .B(p_input[427]), .Z(n4812) );
  XOR U4736 ( .A(n4814), .B(n4815), .Z(n4810) );
  AND U4737 ( .A(n4816), .B(n4817), .Z(n4815) );
  XNOR U4738 ( .A(p_input[442]), .B(n4814), .Z(n4817) );
  XOR U4739 ( .A(n4814), .B(p_input[426]), .Z(n4816) );
  XOR U4740 ( .A(n4818), .B(n4819), .Z(n4814) );
  AND U4741 ( .A(n4820), .B(n4821), .Z(n4819) );
  XNOR U4742 ( .A(p_input[441]), .B(n4818), .Z(n4821) );
  XOR U4743 ( .A(n4818), .B(p_input[425]), .Z(n4820) );
  XOR U4744 ( .A(n4822), .B(n4823), .Z(n4818) );
  AND U4745 ( .A(n4824), .B(n4825), .Z(n4823) );
  XNOR U4746 ( .A(p_input[440]), .B(n4822), .Z(n4825) );
  XOR U4747 ( .A(n4822), .B(p_input[424]), .Z(n4824) );
  XOR U4748 ( .A(n4826), .B(n4827), .Z(n4822) );
  AND U4749 ( .A(n4828), .B(n4829), .Z(n4827) );
  XNOR U4750 ( .A(p_input[439]), .B(n4826), .Z(n4829) );
  XOR U4751 ( .A(n4826), .B(p_input[423]), .Z(n4828) );
  XOR U4752 ( .A(n4830), .B(n4831), .Z(n4826) );
  AND U4753 ( .A(n4832), .B(n4833), .Z(n4831) );
  XNOR U4754 ( .A(p_input[438]), .B(n4830), .Z(n4833) );
  XOR U4755 ( .A(n4830), .B(p_input[422]), .Z(n4832) );
  XOR U4756 ( .A(n4834), .B(n4835), .Z(n4830) );
  AND U4757 ( .A(n4836), .B(n4837), .Z(n4835) );
  XNOR U4758 ( .A(p_input[437]), .B(n4834), .Z(n4837) );
  XOR U4759 ( .A(n4834), .B(p_input[421]), .Z(n4836) );
  XOR U4760 ( .A(n4838), .B(n4839), .Z(n4834) );
  AND U4761 ( .A(n4840), .B(n4841), .Z(n4839) );
  XNOR U4762 ( .A(p_input[436]), .B(n4838), .Z(n4841) );
  XOR U4763 ( .A(n4838), .B(p_input[420]), .Z(n4840) );
  XOR U4764 ( .A(n4842), .B(n4843), .Z(n4838) );
  AND U4765 ( .A(n4844), .B(n4845), .Z(n4843) );
  XNOR U4766 ( .A(p_input[435]), .B(n4842), .Z(n4845) );
  XOR U4767 ( .A(n4842), .B(p_input[419]), .Z(n4844) );
  XOR U4768 ( .A(n4846), .B(n4847), .Z(n4842) );
  AND U4769 ( .A(n4848), .B(n4849), .Z(n4847) );
  XNOR U4770 ( .A(p_input[434]), .B(n4846), .Z(n4849) );
  XOR U4771 ( .A(n4846), .B(p_input[418]), .Z(n4848) );
  XNOR U4772 ( .A(n4850), .B(n4851), .Z(n4846) );
  AND U4773 ( .A(n4852), .B(n4853), .Z(n4851) );
  XOR U4774 ( .A(p_input[433]), .B(n4850), .Z(n4853) );
  XNOR U4775 ( .A(p_input[417]), .B(n4850), .Z(n4852) );
  AND U4776 ( .A(p_input[432]), .B(n4854), .Z(n4850) );
  IV U4777 ( .A(p_input[416]), .Z(n4854) );
  XNOR U4778 ( .A(p_input[384]), .B(n4855), .Z(n4657) );
  AND U4779 ( .A(n219), .B(n4856), .Z(n4855) );
  XOR U4780 ( .A(p_input[400]), .B(p_input[384]), .Z(n4856) );
  XOR U4781 ( .A(n4857), .B(n4858), .Z(n219) );
  AND U4782 ( .A(n4859), .B(n4860), .Z(n4858) );
  XNOR U4783 ( .A(p_input[415]), .B(n4857), .Z(n4860) );
  XOR U4784 ( .A(n4857), .B(p_input[399]), .Z(n4859) );
  XOR U4785 ( .A(n4861), .B(n4862), .Z(n4857) );
  AND U4786 ( .A(n4863), .B(n4864), .Z(n4862) );
  XNOR U4787 ( .A(p_input[414]), .B(n4861), .Z(n4864) );
  XNOR U4788 ( .A(n4861), .B(n4671), .Z(n4863) );
  IV U4789 ( .A(p_input[398]), .Z(n4671) );
  XOR U4790 ( .A(n4865), .B(n4866), .Z(n4861) );
  AND U4791 ( .A(n4867), .B(n4868), .Z(n4866) );
  XNOR U4792 ( .A(p_input[413]), .B(n4865), .Z(n4868) );
  XNOR U4793 ( .A(n4865), .B(n4680), .Z(n4867) );
  IV U4794 ( .A(p_input[397]), .Z(n4680) );
  XOR U4795 ( .A(n4869), .B(n4870), .Z(n4865) );
  AND U4796 ( .A(n4871), .B(n4872), .Z(n4870) );
  XNOR U4797 ( .A(p_input[412]), .B(n4869), .Z(n4872) );
  XNOR U4798 ( .A(n4869), .B(n4689), .Z(n4871) );
  IV U4799 ( .A(p_input[396]), .Z(n4689) );
  XOR U4800 ( .A(n4873), .B(n4874), .Z(n4869) );
  AND U4801 ( .A(n4875), .B(n4876), .Z(n4874) );
  XNOR U4802 ( .A(p_input[411]), .B(n4873), .Z(n4876) );
  XNOR U4803 ( .A(n4873), .B(n4698), .Z(n4875) );
  IV U4804 ( .A(p_input[395]), .Z(n4698) );
  XOR U4805 ( .A(n4877), .B(n4878), .Z(n4873) );
  AND U4806 ( .A(n4879), .B(n4880), .Z(n4878) );
  XNOR U4807 ( .A(p_input[410]), .B(n4877), .Z(n4880) );
  XNOR U4808 ( .A(n4877), .B(n4707), .Z(n4879) );
  IV U4809 ( .A(p_input[394]), .Z(n4707) );
  XOR U4810 ( .A(n4881), .B(n4882), .Z(n4877) );
  AND U4811 ( .A(n4883), .B(n4884), .Z(n4882) );
  XNOR U4812 ( .A(p_input[409]), .B(n4881), .Z(n4884) );
  XNOR U4813 ( .A(n4881), .B(n4716), .Z(n4883) );
  IV U4814 ( .A(p_input[393]), .Z(n4716) );
  XOR U4815 ( .A(n4885), .B(n4886), .Z(n4881) );
  AND U4816 ( .A(n4887), .B(n4888), .Z(n4886) );
  XNOR U4817 ( .A(p_input[408]), .B(n4885), .Z(n4888) );
  XNOR U4818 ( .A(n4885), .B(n4725), .Z(n4887) );
  IV U4819 ( .A(p_input[392]), .Z(n4725) );
  XOR U4820 ( .A(n4889), .B(n4890), .Z(n4885) );
  AND U4821 ( .A(n4891), .B(n4892), .Z(n4890) );
  XNOR U4822 ( .A(p_input[407]), .B(n4889), .Z(n4892) );
  XNOR U4823 ( .A(n4889), .B(n4734), .Z(n4891) );
  IV U4824 ( .A(p_input[391]), .Z(n4734) );
  XOR U4825 ( .A(n4893), .B(n4894), .Z(n4889) );
  AND U4826 ( .A(n4895), .B(n4896), .Z(n4894) );
  XNOR U4827 ( .A(p_input[406]), .B(n4893), .Z(n4896) );
  XNOR U4828 ( .A(n4893), .B(n4743), .Z(n4895) );
  IV U4829 ( .A(p_input[390]), .Z(n4743) );
  XOR U4830 ( .A(n4897), .B(n4898), .Z(n4893) );
  AND U4831 ( .A(n4899), .B(n4900), .Z(n4898) );
  XNOR U4832 ( .A(p_input[405]), .B(n4897), .Z(n4900) );
  XNOR U4833 ( .A(n4897), .B(n4752), .Z(n4899) );
  IV U4834 ( .A(p_input[389]), .Z(n4752) );
  XOR U4835 ( .A(n4901), .B(n4902), .Z(n4897) );
  AND U4836 ( .A(n4903), .B(n4904), .Z(n4902) );
  XNOR U4837 ( .A(p_input[404]), .B(n4901), .Z(n4904) );
  XNOR U4838 ( .A(n4901), .B(n4761), .Z(n4903) );
  IV U4839 ( .A(p_input[388]), .Z(n4761) );
  XOR U4840 ( .A(n4905), .B(n4906), .Z(n4901) );
  AND U4841 ( .A(n4907), .B(n4908), .Z(n4906) );
  XNOR U4842 ( .A(p_input[403]), .B(n4905), .Z(n4908) );
  XNOR U4843 ( .A(n4905), .B(n4770), .Z(n4907) );
  IV U4844 ( .A(p_input[387]), .Z(n4770) );
  XOR U4845 ( .A(n4909), .B(n4910), .Z(n4905) );
  AND U4846 ( .A(n4911), .B(n4912), .Z(n4910) );
  XNOR U4847 ( .A(p_input[402]), .B(n4909), .Z(n4912) );
  XNOR U4848 ( .A(n4909), .B(n4779), .Z(n4911) );
  IV U4849 ( .A(p_input[386]), .Z(n4779) );
  XNOR U4850 ( .A(n4913), .B(n4914), .Z(n4909) );
  AND U4851 ( .A(n4915), .B(n4916), .Z(n4914) );
  XOR U4852 ( .A(p_input[401]), .B(n4913), .Z(n4916) );
  XNOR U4853 ( .A(p_input[385]), .B(n4913), .Z(n4915) );
  AND U4854 ( .A(p_input[400]), .B(n4917), .Z(n4913) );
  IV U4855 ( .A(p_input[384]), .Z(n4917) );
  XOR U4856 ( .A(n4918), .B(n4919), .Z(n4033) );
  AND U4857 ( .A(n256), .B(n4920), .Z(n4919) );
  XNOR U4858 ( .A(n4921), .B(n4918), .Z(n4920) );
  XOR U4859 ( .A(n4922), .B(n4923), .Z(n256) );
  AND U4860 ( .A(n4924), .B(n4925), .Z(n4923) );
  XNOR U4861 ( .A(n4045), .B(n4922), .Z(n4925) );
  AND U4862 ( .A(n4926), .B(n4927), .Z(n4045) );
  XOR U4863 ( .A(n4922), .B(n4044), .Z(n4924) );
  AND U4864 ( .A(n4928), .B(n4929), .Z(n4044) );
  XOR U4865 ( .A(n4930), .B(n4931), .Z(n4922) );
  AND U4866 ( .A(n4932), .B(n4933), .Z(n4931) );
  XOR U4867 ( .A(n4930), .B(n4057), .Z(n4933) );
  XOR U4868 ( .A(n4934), .B(n4935), .Z(n4057) );
  AND U4869 ( .A(n190), .B(n4936), .Z(n4935) );
  XOR U4870 ( .A(n4937), .B(n4934), .Z(n4936) );
  XNOR U4871 ( .A(n4054), .B(n4930), .Z(n4932) );
  XOR U4872 ( .A(n4938), .B(n4939), .Z(n4054) );
  AND U4873 ( .A(n187), .B(n4940), .Z(n4939) );
  XOR U4874 ( .A(n4941), .B(n4938), .Z(n4940) );
  XOR U4875 ( .A(n4942), .B(n4943), .Z(n4930) );
  AND U4876 ( .A(n4944), .B(n4945), .Z(n4943) );
  XOR U4877 ( .A(n4942), .B(n4069), .Z(n4945) );
  XOR U4878 ( .A(n4946), .B(n4947), .Z(n4069) );
  AND U4879 ( .A(n190), .B(n4948), .Z(n4947) );
  XOR U4880 ( .A(n4949), .B(n4946), .Z(n4948) );
  XNOR U4881 ( .A(n4066), .B(n4942), .Z(n4944) );
  XOR U4882 ( .A(n4950), .B(n4951), .Z(n4066) );
  AND U4883 ( .A(n187), .B(n4952), .Z(n4951) );
  XOR U4884 ( .A(n4953), .B(n4950), .Z(n4952) );
  XOR U4885 ( .A(n4954), .B(n4955), .Z(n4942) );
  AND U4886 ( .A(n4956), .B(n4957), .Z(n4955) );
  XOR U4887 ( .A(n4954), .B(n4081), .Z(n4957) );
  XOR U4888 ( .A(n4958), .B(n4959), .Z(n4081) );
  AND U4889 ( .A(n190), .B(n4960), .Z(n4959) );
  XOR U4890 ( .A(n4961), .B(n4958), .Z(n4960) );
  XNOR U4891 ( .A(n4078), .B(n4954), .Z(n4956) );
  XOR U4892 ( .A(n4962), .B(n4963), .Z(n4078) );
  AND U4893 ( .A(n187), .B(n4964), .Z(n4963) );
  XOR U4894 ( .A(n4965), .B(n4962), .Z(n4964) );
  XOR U4895 ( .A(n4966), .B(n4967), .Z(n4954) );
  AND U4896 ( .A(n4968), .B(n4969), .Z(n4967) );
  XOR U4897 ( .A(n4966), .B(n4093), .Z(n4969) );
  XOR U4898 ( .A(n4970), .B(n4971), .Z(n4093) );
  AND U4899 ( .A(n190), .B(n4972), .Z(n4971) );
  XOR U4900 ( .A(n4973), .B(n4970), .Z(n4972) );
  XNOR U4901 ( .A(n4090), .B(n4966), .Z(n4968) );
  XOR U4902 ( .A(n4974), .B(n4975), .Z(n4090) );
  AND U4903 ( .A(n187), .B(n4976), .Z(n4975) );
  XOR U4904 ( .A(n4977), .B(n4974), .Z(n4976) );
  XOR U4905 ( .A(n4978), .B(n4979), .Z(n4966) );
  AND U4906 ( .A(n4980), .B(n4981), .Z(n4979) );
  XOR U4907 ( .A(n4978), .B(n4105), .Z(n4981) );
  XOR U4908 ( .A(n4982), .B(n4983), .Z(n4105) );
  AND U4909 ( .A(n190), .B(n4984), .Z(n4983) );
  XOR U4910 ( .A(n4985), .B(n4982), .Z(n4984) );
  XNOR U4911 ( .A(n4102), .B(n4978), .Z(n4980) );
  XOR U4912 ( .A(n4986), .B(n4987), .Z(n4102) );
  AND U4913 ( .A(n187), .B(n4988), .Z(n4987) );
  XOR U4914 ( .A(n4989), .B(n4986), .Z(n4988) );
  XOR U4915 ( .A(n4990), .B(n4991), .Z(n4978) );
  AND U4916 ( .A(n4992), .B(n4993), .Z(n4991) );
  XOR U4917 ( .A(n4990), .B(n4117), .Z(n4993) );
  XOR U4918 ( .A(n4994), .B(n4995), .Z(n4117) );
  AND U4919 ( .A(n190), .B(n4996), .Z(n4995) );
  XOR U4920 ( .A(n4997), .B(n4994), .Z(n4996) );
  XNOR U4921 ( .A(n4114), .B(n4990), .Z(n4992) );
  XOR U4922 ( .A(n4998), .B(n4999), .Z(n4114) );
  AND U4923 ( .A(n187), .B(n5000), .Z(n4999) );
  XOR U4924 ( .A(n5001), .B(n4998), .Z(n5000) );
  XOR U4925 ( .A(n5002), .B(n5003), .Z(n4990) );
  AND U4926 ( .A(n5004), .B(n5005), .Z(n5003) );
  XOR U4927 ( .A(n5002), .B(n4129), .Z(n5005) );
  XOR U4928 ( .A(n5006), .B(n5007), .Z(n4129) );
  AND U4929 ( .A(n190), .B(n5008), .Z(n5007) );
  XOR U4930 ( .A(n5009), .B(n5006), .Z(n5008) );
  XNOR U4931 ( .A(n4126), .B(n5002), .Z(n5004) );
  XOR U4932 ( .A(n5010), .B(n5011), .Z(n4126) );
  AND U4933 ( .A(n187), .B(n5012), .Z(n5011) );
  XOR U4934 ( .A(n5013), .B(n5010), .Z(n5012) );
  XOR U4935 ( .A(n5014), .B(n5015), .Z(n5002) );
  AND U4936 ( .A(n5016), .B(n5017), .Z(n5015) );
  XOR U4937 ( .A(n5014), .B(n4141), .Z(n5017) );
  XOR U4938 ( .A(n5018), .B(n5019), .Z(n4141) );
  AND U4939 ( .A(n190), .B(n5020), .Z(n5019) );
  XOR U4940 ( .A(n5021), .B(n5018), .Z(n5020) );
  XNOR U4941 ( .A(n4138), .B(n5014), .Z(n5016) );
  XOR U4942 ( .A(n5022), .B(n5023), .Z(n4138) );
  AND U4943 ( .A(n187), .B(n5024), .Z(n5023) );
  XOR U4944 ( .A(n5025), .B(n5022), .Z(n5024) );
  XOR U4945 ( .A(n5026), .B(n5027), .Z(n5014) );
  AND U4946 ( .A(n5028), .B(n5029), .Z(n5027) );
  XOR U4947 ( .A(n5026), .B(n4153), .Z(n5029) );
  XOR U4948 ( .A(n5030), .B(n5031), .Z(n4153) );
  AND U4949 ( .A(n190), .B(n5032), .Z(n5031) );
  XOR U4950 ( .A(n5033), .B(n5030), .Z(n5032) );
  XNOR U4951 ( .A(n4150), .B(n5026), .Z(n5028) );
  XOR U4952 ( .A(n5034), .B(n5035), .Z(n4150) );
  AND U4953 ( .A(n187), .B(n5036), .Z(n5035) );
  XOR U4954 ( .A(n5037), .B(n5034), .Z(n5036) );
  XOR U4955 ( .A(n5038), .B(n5039), .Z(n5026) );
  AND U4956 ( .A(n5040), .B(n5041), .Z(n5039) );
  XOR U4957 ( .A(n5038), .B(n4165), .Z(n5041) );
  XOR U4958 ( .A(n5042), .B(n5043), .Z(n4165) );
  AND U4959 ( .A(n190), .B(n5044), .Z(n5043) );
  XOR U4960 ( .A(n5045), .B(n5042), .Z(n5044) );
  XNOR U4961 ( .A(n4162), .B(n5038), .Z(n5040) );
  XOR U4962 ( .A(n5046), .B(n5047), .Z(n4162) );
  AND U4963 ( .A(n187), .B(n5048), .Z(n5047) );
  XOR U4964 ( .A(n5049), .B(n5046), .Z(n5048) );
  XOR U4965 ( .A(n5050), .B(n5051), .Z(n5038) );
  AND U4966 ( .A(n5052), .B(n5053), .Z(n5051) );
  XOR U4967 ( .A(n5050), .B(n4177), .Z(n5053) );
  XOR U4968 ( .A(n5054), .B(n5055), .Z(n4177) );
  AND U4969 ( .A(n190), .B(n5056), .Z(n5055) );
  XOR U4970 ( .A(n5057), .B(n5054), .Z(n5056) );
  XNOR U4971 ( .A(n4174), .B(n5050), .Z(n5052) );
  XOR U4972 ( .A(n5058), .B(n5059), .Z(n4174) );
  AND U4973 ( .A(n187), .B(n5060), .Z(n5059) );
  XOR U4974 ( .A(n5061), .B(n5058), .Z(n5060) );
  XOR U4975 ( .A(n5062), .B(n5063), .Z(n5050) );
  AND U4976 ( .A(n5064), .B(n5065), .Z(n5063) );
  XOR U4977 ( .A(n4189), .B(n5062), .Z(n5065) );
  XOR U4978 ( .A(n5066), .B(n5067), .Z(n4189) );
  AND U4979 ( .A(n190), .B(n5068), .Z(n5067) );
  XOR U4980 ( .A(n5066), .B(n5069), .Z(n5068) );
  XNOR U4981 ( .A(n5062), .B(n4186), .Z(n5064) );
  XOR U4982 ( .A(n5070), .B(n5071), .Z(n4186) );
  AND U4983 ( .A(n187), .B(n5072), .Z(n5071) );
  XOR U4984 ( .A(n5070), .B(n5073), .Z(n5072) );
  XOR U4985 ( .A(n5074), .B(n5075), .Z(n5062) );
  AND U4986 ( .A(n5076), .B(n5077), .Z(n5075) );
  XOR U4987 ( .A(n5074), .B(n4201), .Z(n5077) );
  XOR U4988 ( .A(n5078), .B(n5079), .Z(n4201) );
  AND U4989 ( .A(n190), .B(n5080), .Z(n5079) );
  XOR U4990 ( .A(n5081), .B(n5078), .Z(n5080) );
  XNOR U4991 ( .A(n4198), .B(n5074), .Z(n5076) );
  XOR U4992 ( .A(n5082), .B(n5083), .Z(n4198) );
  AND U4993 ( .A(n187), .B(n5084), .Z(n5083) );
  XOR U4994 ( .A(n5085), .B(n5082), .Z(n5084) );
  XOR U4995 ( .A(n5086), .B(n5087), .Z(n5074) );
  AND U4996 ( .A(n5088), .B(n5089), .Z(n5087) );
  XNOR U4997 ( .A(n5090), .B(n4214), .Z(n5089) );
  XOR U4998 ( .A(n5091), .B(n5092), .Z(n4214) );
  AND U4999 ( .A(n190), .B(n5093), .Z(n5092) );
  XOR U5000 ( .A(n5094), .B(n5091), .Z(n5093) );
  XNOR U5001 ( .A(n4211), .B(n5086), .Z(n5088) );
  XOR U5002 ( .A(n5095), .B(n5096), .Z(n4211) );
  AND U5003 ( .A(n187), .B(n5097), .Z(n5096) );
  XOR U5004 ( .A(n5098), .B(n5095), .Z(n5097) );
  IV U5005 ( .A(n5090), .Z(n5086) );
  AND U5006 ( .A(n4918), .B(n4921), .Z(n5090) );
  XNOR U5007 ( .A(n5099), .B(n5100), .Z(n4921) );
  AND U5008 ( .A(n190), .B(n5101), .Z(n5100) );
  XNOR U5009 ( .A(n5102), .B(n5099), .Z(n5101) );
  XOR U5010 ( .A(n5103), .B(n5104), .Z(n190) );
  AND U5011 ( .A(n5105), .B(n5106), .Z(n5104) );
  XNOR U5012 ( .A(n4926), .B(n5103), .Z(n5106) );
  AND U5013 ( .A(p_input[383]), .B(p_input[367]), .Z(n4926) );
  XOR U5014 ( .A(n5103), .B(n4927), .Z(n5105) );
  AND U5015 ( .A(p_input[351]), .B(p_input[335]), .Z(n4927) );
  XOR U5016 ( .A(n5107), .B(n5108), .Z(n5103) );
  AND U5017 ( .A(n5109), .B(n5110), .Z(n5108) );
  XOR U5018 ( .A(n5107), .B(n4937), .Z(n5110) );
  XNOR U5019 ( .A(p_input[366]), .B(n5111), .Z(n4937) );
  AND U5020 ( .A(n230), .B(n5112), .Z(n5111) );
  XOR U5021 ( .A(p_input[382]), .B(p_input[366]), .Z(n5112) );
  XNOR U5022 ( .A(n4934), .B(n5107), .Z(n5109) );
  XOR U5023 ( .A(n5113), .B(n5114), .Z(n4934) );
  AND U5024 ( .A(n228), .B(n5115), .Z(n5114) );
  XOR U5025 ( .A(p_input[350]), .B(p_input[334]), .Z(n5115) );
  XOR U5026 ( .A(n5116), .B(n5117), .Z(n5107) );
  AND U5027 ( .A(n5118), .B(n5119), .Z(n5117) );
  XOR U5028 ( .A(n5116), .B(n4949), .Z(n5119) );
  XNOR U5029 ( .A(p_input[365]), .B(n5120), .Z(n4949) );
  AND U5030 ( .A(n230), .B(n5121), .Z(n5120) );
  XOR U5031 ( .A(p_input[381]), .B(p_input[365]), .Z(n5121) );
  XNOR U5032 ( .A(n4946), .B(n5116), .Z(n5118) );
  XOR U5033 ( .A(n5122), .B(n5123), .Z(n4946) );
  AND U5034 ( .A(n228), .B(n5124), .Z(n5123) );
  XOR U5035 ( .A(p_input[349]), .B(p_input[333]), .Z(n5124) );
  XOR U5036 ( .A(n5125), .B(n5126), .Z(n5116) );
  AND U5037 ( .A(n5127), .B(n5128), .Z(n5126) );
  XOR U5038 ( .A(n5125), .B(n4961), .Z(n5128) );
  XNOR U5039 ( .A(p_input[364]), .B(n5129), .Z(n4961) );
  AND U5040 ( .A(n230), .B(n5130), .Z(n5129) );
  XOR U5041 ( .A(p_input[380]), .B(p_input[364]), .Z(n5130) );
  XNOR U5042 ( .A(n4958), .B(n5125), .Z(n5127) );
  XOR U5043 ( .A(n5131), .B(n5132), .Z(n4958) );
  AND U5044 ( .A(n228), .B(n5133), .Z(n5132) );
  XOR U5045 ( .A(p_input[348]), .B(p_input[332]), .Z(n5133) );
  XOR U5046 ( .A(n5134), .B(n5135), .Z(n5125) );
  AND U5047 ( .A(n5136), .B(n5137), .Z(n5135) );
  XOR U5048 ( .A(n5134), .B(n4973), .Z(n5137) );
  XNOR U5049 ( .A(p_input[363]), .B(n5138), .Z(n4973) );
  AND U5050 ( .A(n230), .B(n5139), .Z(n5138) );
  XOR U5051 ( .A(p_input[379]), .B(p_input[363]), .Z(n5139) );
  XNOR U5052 ( .A(n4970), .B(n5134), .Z(n5136) );
  XOR U5053 ( .A(n5140), .B(n5141), .Z(n4970) );
  AND U5054 ( .A(n228), .B(n5142), .Z(n5141) );
  XOR U5055 ( .A(p_input[347]), .B(p_input[331]), .Z(n5142) );
  XOR U5056 ( .A(n5143), .B(n5144), .Z(n5134) );
  AND U5057 ( .A(n5145), .B(n5146), .Z(n5144) );
  XOR U5058 ( .A(n5143), .B(n4985), .Z(n5146) );
  XNOR U5059 ( .A(p_input[362]), .B(n5147), .Z(n4985) );
  AND U5060 ( .A(n230), .B(n5148), .Z(n5147) );
  XOR U5061 ( .A(p_input[378]), .B(p_input[362]), .Z(n5148) );
  XNOR U5062 ( .A(n4982), .B(n5143), .Z(n5145) );
  XOR U5063 ( .A(n5149), .B(n5150), .Z(n4982) );
  AND U5064 ( .A(n228), .B(n5151), .Z(n5150) );
  XOR U5065 ( .A(p_input[346]), .B(p_input[330]), .Z(n5151) );
  XOR U5066 ( .A(n5152), .B(n5153), .Z(n5143) );
  AND U5067 ( .A(n5154), .B(n5155), .Z(n5153) );
  XOR U5068 ( .A(n5152), .B(n4997), .Z(n5155) );
  XNOR U5069 ( .A(p_input[361]), .B(n5156), .Z(n4997) );
  AND U5070 ( .A(n230), .B(n5157), .Z(n5156) );
  XOR U5071 ( .A(p_input[377]), .B(p_input[361]), .Z(n5157) );
  XNOR U5072 ( .A(n4994), .B(n5152), .Z(n5154) );
  XOR U5073 ( .A(n5158), .B(n5159), .Z(n4994) );
  AND U5074 ( .A(n228), .B(n5160), .Z(n5159) );
  XOR U5075 ( .A(p_input[345]), .B(p_input[329]), .Z(n5160) );
  XOR U5076 ( .A(n5161), .B(n5162), .Z(n5152) );
  AND U5077 ( .A(n5163), .B(n5164), .Z(n5162) );
  XOR U5078 ( .A(n5161), .B(n5009), .Z(n5164) );
  XNOR U5079 ( .A(p_input[360]), .B(n5165), .Z(n5009) );
  AND U5080 ( .A(n230), .B(n5166), .Z(n5165) );
  XOR U5081 ( .A(p_input[376]), .B(p_input[360]), .Z(n5166) );
  XNOR U5082 ( .A(n5006), .B(n5161), .Z(n5163) );
  XOR U5083 ( .A(n5167), .B(n5168), .Z(n5006) );
  AND U5084 ( .A(n228), .B(n5169), .Z(n5168) );
  XOR U5085 ( .A(p_input[344]), .B(p_input[328]), .Z(n5169) );
  XOR U5086 ( .A(n5170), .B(n5171), .Z(n5161) );
  AND U5087 ( .A(n5172), .B(n5173), .Z(n5171) );
  XOR U5088 ( .A(n5170), .B(n5021), .Z(n5173) );
  XNOR U5089 ( .A(p_input[359]), .B(n5174), .Z(n5021) );
  AND U5090 ( .A(n230), .B(n5175), .Z(n5174) );
  XOR U5091 ( .A(p_input[375]), .B(p_input[359]), .Z(n5175) );
  XNOR U5092 ( .A(n5018), .B(n5170), .Z(n5172) );
  XOR U5093 ( .A(n5176), .B(n5177), .Z(n5018) );
  AND U5094 ( .A(n228), .B(n5178), .Z(n5177) );
  XOR U5095 ( .A(p_input[343]), .B(p_input[327]), .Z(n5178) );
  XOR U5096 ( .A(n5179), .B(n5180), .Z(n5170) );
  AND U5097 ( .A(n5181), .B(n5182), .Z(n5180) );
  XOR U5098 ( .A(n5179), .B(n5033), .Z(n5182) );
  XNOR U5099 ( .A(p_input[358]), .B(n5183), .Z(n5033) );
  AND U5100 ( .A(n230), .B(n5184), .Z(n5183) );
  XOR U5101 ( .A(p_input[374]), .B(p_input[358]), .Z(n5184) );
  XNOR U5102 ( .A(n5030), .B(n5179), .Z(n5181) );
  XOR U5103 ( .A(n5185), .B(n5186), .Z(n5030) );
  AND U5104 ( .A(n228), .B(n5187), .Z(n5186) );
  XOR U5105 ( .A(p_input[342]), .B(p_input[326]), .Z(n5187) );
  XOR U5106 ( .A(n5188), .B(n5189), .Z(n5179) );
  AND U5107 ( .A(n5190), .B(n5191), .Z(n5189) );
  XOR U5108 ( .A(n5188), .B(n5045), .Z(n5191) );
  XNOR U5109 ( .A(p_input[357]), .B(n5192), .Z(n5045) );
  AND U5110 ( .A(n230), .B(n5193), .Z(n5192) );
  XOR U5111 ( .A(p_input[373]), .B(p_input[357]), .Z(n5193) );
  XNOR U5112 ( .A(n5042), .B(n5188), .Z(n5190) );
  XOR U5113 ( .A(n5194), .B(n5195), .Z(n5042) );
  AND U5114 ( .A(n228), .B(n5196), .Z(n5195) );
  XOR U5115 ( .A(p_input[341]), .B(p_input[325]), .Z(n5196) );
  XOR U5116 ( .A(n5197), .B(n5198), .Z(n5188) );
  AND U5117 ( .A(n5199), .B(n5200), .Z(n5198) );
  XOR U5118 ( .A(n5197), .B(n5057), .Z(n5200) );
  XNOR U5119 ( .A(p_input[356]), .B(n5201), .Z(n5057) );
  AND U5120 ( .A(n230), .B(n5202), .Z(n5201) );
  XOR U5121 ( .A(p_input[372]), .B(p_input[356]), .Z(n5202) );
  XNOR U5122 ( .A(n5054), .B(n5197), .Z(n5199) );
  XOR U5123 ( .A(n5203), .B(n5204), .Z(n5054) );
  AND U5124 ( .A(n228), .B(n5205), .Z(n5204) );
  XOR U5125 ( .A(p_input[340]), .B(p_input[324]), .Z(n5205) );
  XOR U5126 ( .A(n5206), .B(n5207), .Z(n5197) );
  AND U5127 ( .A(n5208), .B(n5209), .Z(n5207) );
  XOR U5128 ( .A(n5069), .B(n5206), .Z(n5209) );
  XNOR U5129 ( .A(p_input[355]), .B(n5210), .Z(n5069) );
  AND U5130 ( .A(n230), .B(n5211), .Z(n5210) );
  XOR U5131 ( .A(p_input[371]), .B(p_input[355]), .Z(n5211) );
  XNOR U5132 ( .A(n5206), .B(n5066), .Z(n5208) );
  XOR U5133 ( .A(n5212), .B(n5213), .Z(n5066) );
  AND U5134 ( .A(n228), .B(n5214), .Z(n5213) );
  XOR U5135 ( .A(p_input[339]), .B(p_input[323]), .Z(n5214) );
  XOR U5136 ( .A(n5215), .B(n5216), .Z(n5206) );
  AND U5137 ( .A(n5217), .B(n5218), .Z(n5216) );
  XOR U5138 ( .A(n5215), .B(n5081), .Z(n5218) );
  XNOR U5139 ( .A(p_input[354]), .B(n5219), .Z(n5081) );
  AND U5140 ( .A(n230), .B(n5220), .Z(n5219) );
  XOR U5141 ( .A(p_input[370]), .B(p_input[354]), .Z(n5220) );
  XNOR U5142 ( .A(n5078), .B(n5215), .Z(n5217) );
  XOR U5143 ( .A(n5221), .B(n5222), .Z(n5078) );
  AND U5144 ( .A(n228), .B(n5223), .Z(n5222) );
  XOR U5145 ( .A(p_input[338]), .B(p_input[322]), .Z(n5223) );
  XOR U5146 ( .A(n5224), .B(n5225), .Z(n5215) );
  AND U5147 ( .A(n5226), .B(n5227), .Z(n5225) );
  XNOR U5148 ( .A(n5228), .B(n5094), .Z(n5227) );
  XNOR U5149 ( .A(p_input[353]), .B(n5229), .Z(n5094) );
  AND U5150 ( .A(n230), .B(n5230), .Z(n5229) );
  XNOR U5151 ( .A(p_input[369]), .B(n5231), .Z(n5230) );
  IV U5152 ( .A(p_input[353]), .Z(n5231) );
  XNOR U5153 ( .A(n5091), .B(n5224), .Z(n5226) );
  XNOR U5154 ( .A(p_input[321]), .B(n5232), .Z(n5091) );
  AND U5155 ( .A(n228), .B(n5233), .Z(n5232) );
  XOR U5156 ( .A(p_input[337]), .B(p_input[321]), .Z(n5233) );
  IV U5157 ( .A(n5228), .Z(n5224) );
  AND U5158 ( .A(n5099), .B(n5102), .Z(n5228) );
  XOR U5159 ( .A(p_input[352]), .B(n5234), .Z(n5102) );
  AND U5160 ( .A(n230), .B(n5235), .Z(n5234) );
  XOR U5161 ( .A(p_input[368]), .B(p_input[352]), .Z(n5235) );
  XOR U5162 ( .A(n5236), .B(n5237), .Z(n230) );
  AND U5163 ( .A(n5238), .B(n5239), .Z(n5237) );
  XNOR U5164 ( .A(p_input[383]), .B(n5236), .Z(n5239) );
  XOR U5165 ( .A(n5236), .B(p_input[367]), .Z(n5238) );
  XOR U5166 ( .A(n5240), .B(n5241), .Z(n5236) );
  AND U5167 ( .A(n5242), .B(n5243), .Z(n5241) );
  XNOR U5168 ( .A(p_input[382]), .B(n5240), .Z(n5243) );
  XOR U5169 ( .A(n5240), .B(p_input[366]), .Z(n5242) );
  XOR U5170 ( .A(n5244), .B(n5245), .Z(n5240) );
  AND U5171 ( .A(n5246), .B(n5247), .Z(n5245) );
  XNOR U5172 ( .A(p_input[381]), .B(n5244), .Z(n5247) );
  XOR U5173 ( .A(n5244), .B(p_input[365]), .Z(n5246) );
  XOR U5174 ( .A(n5248), .B(n5249), .Z(n5244) );
  AND U5175 ( .A(n5250), .B(n5251), .Z(n5249) );
  XNOR U5176 ( .A(p_input[380]), .B(n5248), .Z(n5251) );
  XOR U5177 ( .A(n5248), .B(p_input[364]), .Z(n5250) );
  XOR U5178 ( .A(n5252), .B(n5253), .Z(n5248) );
  AND U5179 ( .A(n5254), .B(n5255), .Z(n5253) );
  XNOR U5180 ( .A(p_input[379]), .B(n5252), .Z(n5255) );
  XOR U5181 ( .A(n5252), .B(p_input[363]), .Z(n5254) );
  XOR U5182 ( .A(n5256), .B(n5257), .Z(n5252) );
  AND U5183 ( .A(n5258), .B(n5259), .Z(n5257) );
  XNOR U5184 ( .A(p_input[378]), .B(n5256), .Z(n5259) );
  XOR U5185 ( .A(n5256), .B(p_input[362]), .Z(n5258) );
  XOR U5186 ( .A(n5260), .B(n5261), .Z(n5256) );
  AND U5187 ( .A(n5262), .B(n5263), .Z(n5261) );
  XNOR U5188 ( .A(p_input[377]), .B(n5260), .Z(n5263) );
  XOR U5189 ( .A(n5260), .B(p_input[361]), .Z(n5262) );
  XOR U5190 ( .A(n5264), .B(n5265), .Z(n5260) );
  AND U5191 ( .A(n5266), .B(n5267), .Z(n5265) );
  XNOR U5192 ( .A(p_input[376]), .B(n5264), .Z(n5267) );
  XOR U5193 ( .A(n5264), .B(p_input[360]), .Z(n5266) );
  XOR U5194 ( .A(n5268), .B(n5269), .Z(n5264) );
  AND U5195 ( .A(n5270), .B(n5271), .Z(n5269) );
  XNOR U5196 ( .A(p_input[375]), .B(n5268), .Z(n5271) );
  XOR U5197 ( .A(n5268), .B(p_input[359]), .Z(n5270) );
  XOR U5198 ( .A(n5272), .B(n5273), .Z(n5268) );
  AND U5199 ( .A(n5274), .B(n5275), .Z(n5273) );
  XNOR U5200 ( .A(p_input[374]), .B(n5272), .Z(n5275) );
  XOR U5201 ( .A(n5272), .B(p_input[358]), .Z(n5274) );
  XOR U5202 ( .A(n5276), .B(n5277), .Z(n5272) );
  AND U5203 ( .A(n5278), .B(n5279), .Z(n5277) );
  XNOR U5204 ( .A(p_input[373]), .B(n5276), .Z(n5279) );
  XOR U5205 ( .A(n5276), .B(p_input[357]), .Z(n5278) );
  XOR U5206 ( .A(n5280), .B(n5281), .Z(n5276) );
  AND U5207 ( .A(n5282), .B(n5283), .Z(n5281) );
  XNOR U5208 ( .A(p_input[372]), .B(n5280), .Z(n5283) );
  XOR U5209 ( .A(n5280), .B(p_input[356]), .Z(n5282) );
  XOR U5210 ( .A(n5284), .B(n5285), .Z(n5280) );
  AND U5211 ( .A(n5286), .B(n5287), .Z(n5285) );
  XNOR U5212 ( .A(p_input[371]), .B(n5284), .Z(n5287) );
  XOR U5213 ( .A(n5284), .B(p_input[355]), .Z(n5286) );
  XOR U5214 ( .A(n5288), .B(n5289), .Z(n5284) );
  AND U5215 ( .A(n5290), .B(n5291), .Z(n5289) );
  XNOR U5216 ( .A(p_input[370]), .B(n5288), .Z(n5291) );
  XOR U5217 ( .A(n5288), .B(p_input[354]), .Z(n5290) );
  XNOR U5218 ( .A(n5292), .B(n5293), .Z(n5288) );
  AND U5219 ( .A(n5294), .B(n5295), .Z(n5293) );
  XOR U5220 ( .A(p_input[369]), .B(n5292), .Z(n5295) );
  XNOR U5221 ( .A(p_input[353]), .B(n5292), .Z(n5294) );
  AND U5222 ( .A(p_input[368]), .B(n5296), .Z(n5292) );
  IV U5223 ( .A(p_input[352]), .Z(n5296) );
  XNOR U5224 ( .A(p_input[320]), .B(n5297), .Z(n5099) );
  AND U5225 ( .A(n228), .B(n5298), .Z(n5297) );
  XOR U5226 ( .A(p_input[336]), .B(p_input[320]), .Z(n5298) );
  XOR U5227 ( .A(n5299), .B(n5300), .Z(n228) );
  AND U5228 ( .A(n5301), .B(n5302), .Z(n5300) );
  XNOR U5229 ( .A(p_input[351]), .B(n5299), .Z(n5302) );
  XOR U5230 ( .A(n5299), .B(p_input[335]), .Z(n5301) );
  XOR U5231 ( .A(n5303), .B(n5304), .Z(n5299) );
  AND U5232 ( .A(n5305), .B(n5306), .Z(n5304) );
  XNOR U5233 ( .A(p_input[350]), .B(n5303), .Z(n5306) );
  XNOR U5234 ( .A(n5303), .B(n5113), .Z(n5305) );
  IV U5235 ( .A(p_input[334]), .Z(n5113) );
  XOR U5236 ( .A(n5307), .B(n5308), .Z(n5303) );
  AND U5237 ( .A(n5309), .B(n5310), .Z(n5308) );
  XNOR U5238 ( .A(p_input[349]), .B(n5307), .Z(n5310) );
  XNOR U5239 ( .A(n5307), .B(n5122), .Z(n5309) );
  IV U5240 ( .A(p_input[333]), .Z(n5122) );
  XOR U5241 ( .A(n5311), .B(n5312), .Z(n5307) );
  AND U5242 ( .A(n5313), .B(n5314), .Z(n5312) );
  XNOR U5243 ( .A(p_input[348]), .B(n5311), .Z(n5314) );
  XNOR U5244 ( .A(n5311), .B(n5131), .Z(n5313) );
  IV U5245 ( .A(p_input[332]), .Z(n5131) );
  XOR U5246 ( .A(n5315), .B(n5316), .Z(n5311) );
  AND U5247 ( .A(n5317), .B(n5318), .Z(n5316) );
  XNOR U5248 ( .A(p_input[347]), .B(n5315), .Z(n5318) );
  XNOR U5249 ( .A(n5315), .B(n5140), .Z(n5317) );
  IV U5250 ( .A(p_input[331]), .Z(n5140) );
  XOR U5251 ( .A(n5319), .B(n5320), .Z(n5315) );
  AND U5252 ( .A(n5321), .B(n5322), .Z(n5320) );
  XNOR U5253 ( .A(p_input[346]), .B(n5319), .Z(n5322) );
  XNOR U5254 ( .A(n5319), .B(n5149), .Z(n5321) );
  IV U5255 ( .A(p_input[330]), .Z(n5149) );
  XOR U5256 ( .A(n5323), .B(n5324), .Z(n5319) );
  AND U5257 ( .A(n5325), .B(n5326), .Z(n5324) );
  XNOR U5258 ( .A(p_input[345]), .B(n5323), .Z(n5326) );
  XNOR U5259 ( .A(n5323), .B(n5158), .Z(n5325) );
  IV U5260 ( .A(p_input[329]), .Z(n5158) );
  XOR U5261 ( .A(n5327), .B(n5328), .Z(n5323) );
  AND U5262 ( .A(n5329), .B(n5330), .Z(n5328) );
  XNOR U5263 ( .A(p_input[344]), .B(n5327), .Z(n5330) );
  XNOR U5264 ( .A(n5327), .B(n5167), .Z(n5329) );
  IV U5265 ( .A(p_input[328]), .Z(n5167) );
  XOR U5266 ( .A(n5331), .B(n5332), .Z(n5327) );
  AND U5267 ( .A(n5333), .B(n5334), .Z(n5332) );
  XNOR U5268 ( .A(p_input[343]), .B(n5331), .Z(n5334) );
  XNOR U5269 ( .A(n5331), .B(n5176), .Z(n5333) );
  IV U5270 ( .A(p_input[327]), .Z(n5176) );
  XOR U5271 ( .A(n5335), .B(n5336), .Z(n5331) );
  AND U5272 ( .A(n5337), .B(n5338), .Z(n5336) );
  XNOR U5273 ( .A(p_input[342]), .B(n5335), .Z(n5338) );
  XNOR U5274 ( .A(n5335), .B(n5185), .Z(n5337) );
  IV U5275 ( .A(p_input[326]), .Z(n5185) );
  XOR U5276 ( .A(n5339), .B(n5340), .Z(n5335) );
  AND U5277 ( .A(n5341), .B(n5342), .Z(n5340) );
  XNOR U5278 ( .A(p_input[341]), .B(n5339), .Z(n5342) );
  XNOR U5279 ( .A(n5339), .B(n5194), .Z(n5341) );
  IV U5280 ( .A(p_input[325]), .Z(n5194) );
  XOR U5281 ( .A(n5343), .B(n5344), .Z(n5339) );
  AND U5282 ( .A(n5345), .B(n5346), .Z(n5344) );
  XNOR U5283 ( .A(p_input[340]), .B(n5343), .Z(n5346) );
  XNOR U5284 ( .A(n5343), .B(n5203), .Z(n5345) );
  IV U5285 ( .A(p_input[324]), .Z(n5203) );
  XOR U5286 ( .A(n5347), .B(n5348), .Z(n5343) );
  AND U5287 ( .A(n5349), .B(n5350), .Z(n5348) );
  XNOR U5288 ( .A(p_input[339]), .B(n5347), .Z(n5350) );
  XNOR U5289 ( .A(n5347), .B(n5212), .Z(n5349) );
  IV U5290 ( .A(p_input[323]), .Z(n5212) );
  XOR U5291 ( .A(n5351), .B(n5352), .Z(n5347) );
  AND U5292 ( .A(n5353), .B(n5354), .Z(n5352) );
  XNOR U5293 ( .A(p_input[338]), .B(n5351), .Z(n5354) );
  XNOR U5294 ( .A(n5351), .B(n5221), .Z(n5353) );
  IV U5295 ( .A(p_input[322]), .Z(n5221) );
  XNOR U5296 ( .A(n5355), .B(n5356), .Z(n5351) );
  AND U5297 ( .A(n5357), .B(n5358), .Z(n5356) );
  XOR U5298 ( .A(p_input[337]), .B(n5355), .Z(n5358) );
  XNOR U5299 ( .A(p_input[321]), .B(n5355), .Z(n5357) );
  AND U5300 ( .A(p_input[336]), .B(n5359), .Z(n5355) );
  IV U5301 ( .A(p_input[320]), .Z(n5359) );
  XOR U5302 ( .A(n5360), .B(n5361), .Z(n4918) );
  AND U5303 ( .A(n187), .B(n5362), .Z(n5361) );
  XNOR U5304 ( .A(n5363), .B(n5360), .Z(n5362) );
  XOR U5305 ( .A(n5364), .B(n5365), .Z(n187) );
  AND U5306 ( .A(n5366), .B(n5367), .Z(n5365) );
  XNOR U5307 ( .A(n4929), .B(n5364), .Z(n5367) );
  AND U5308 ( .A(p_input[319]), .B(p_input[303]), .Z(n4929) );
  XOR U5309 ( .A(n5364), .B(n4928), .Z(n5366) );
  AND U5310 ( .A(p_input[271]), .B(p_input[287]), .Z(n4928) );
  XOR U5311 ( .A(n5368), .B(n5369), .Z(n5364) );
  AND U5312 ( .A(n5370), .B(n5371), .Z(n5369) );
  XOR U5313 ( .A(n5368), .B(n4941), .Z(n5371) );
  XNOR U5314 ( .A(p_input[302]), .B(n5372), .Z(n4941) );
  AND U5315 ( .A(n234), .B(n5373), .Z(n5372) );
  XOR U5316 ( .A(p_input[318]), .B(p_input[302]), .Z(n5373) );
  XNOR U5317 ( .A(n4938), .B(n5368), .Z(n5370) );
  XOR U5318 ( .A(n5374), .B(n5375), .Z(n4938) );
  AND U5319 ( .A(n231), .B(n5376), .Z(n5375) );
  XOR U5320 ( .A(p_input[286]), .B(p_input[270]), .Z(n5376) );
  XOR U5321 ( .A(n5377), .B(n5378), .Z(n5368) );
  AND U5322 ( .A(n5379), .B(n5380), .Z(n5378) );
  XOR U5323 ( .A(n5377), .B(n4953), .Z(n5380) );
  XNOR U5324 ( .A(p_input[301]), .B(n5381), .Z(n4953) );
  AND U5325 ( .A(n234), .B(n5382), .Z(n5381) );
  XOR U5326 ( .A(p_input[317]), .B(p_input[301]), .Z(n5382) );
  XNOR U5327 ( .A(n4950), .B(n5377), .Z(n5379) );
  XOR U5328 ( .A(n5383), .B(n5384), .Z(n4950) );
  AND U5329 ( .A(n231), .B(n5385), .Z(n5384) );
  XOR U5330 ( .A(p_input[285]), .B(p_input[269]), .Z(n5385) );
  XOR U5331 ( .A(n5386), .B(n5387), .Z(n5377) );
  AND U5332 ( .A(n5388), .B(n5389), .Z(n5387) );
  XOR U5333 ( .A(n5386), .B(n4965), .Z(n5389) );
  XNOR U5334 ( .A(p_input[300]), .B(n5390), .Z(n4965) );
  AND U5335 ( .A(n234), .B(n5391), .Z(n5390) );
  XOR U5336 ( .A(p_input[316]), .B(p_input[300]), .Z(n5391) );
  XNOR U5337 ( .A(n4962), .B(n5386), .Z(n5388) );
  XOR U5338 ( .A(n5392), .B(n5393), .Z(n4962) );
  AND U5339 ( .A(n231), .B(n5394), .Z(n5393) );
  XOR U5340 ( .A(p_input[284]), .B(p_input[268]), .Z(n5394) );
  XOR U5341 ( .A(n5395), .B(n5396), .Z(n5386) );
  AND U5342 ( .A(n5397), .B(n5398), .Z(n5396) );
  XOR U5343 ( .A(n5395), .B(n4977), .Z(n5398) );
  XNOR U5344 ( .A(p_input[299]), .B(n5399), .Z(n4977) );
  AND U5345 ( .A(n234), .B(n5400), .Z(n5399) );
  XOR U5346 ( .A(p_input[315]), .B(p_input[299]), .Z(n5400) );
  XNOR U5347 ( .A(n4974), .B(n5395), .Z(n5397) );
  XOR U5348 ( .A(n5401), .B(n5402), .Z(n4974) );
  AND U5349 ( .A(n231), .B(n5403), .Z(n5402) );
  XOR U5350 ( .A(p_input[283]), .B(p_input[267]), .Z(n5403) );
  XOR U5351 ( .A(n5404), .B(n5405), .Z(n5395) );
  AND U5352 ( .A(n5406), .B(n5407), .Z(n5405) );
  XOR U5353 ( .A(n5404), .B(n4989), .Z(n5407) );
  XNOR U5354 ( .A(p_input[298]), .B(n5408), .Z(n4989) );
  AND U5355 ( .A(n234), .B(n5409), .Z(n5408) );
  XOR U5356 ( .A(p_input[314]), .B(p_input[298]), .Z(n5409) );
  XNOR U5357 ( .A(n4986), .B(n5404), .Z(n5406) );
  XOR U5358 ( .A(n5410), .B(n5411), .Z(n4986) );
  AND U5359 ( .A(n231), .B(n5412), .Z(n5411) );
  XOR U5360 ( .A(p_input[282]), .B(p_input[266]), .Z(n5412) );
  XOR U5361 ( .A(n5413), .B(n5414), .Z(n5404) );
  AND U5362 ( .A(n5415), .B(n5416), .Z(n5414) );
  XOR U5363 ( .A(n5413), .B(n5001), .Z(n5416) );
  XNOR U5364 ( .A(p_input[297]), .B(n5417), .Z(n5001) );
  AND U5365 ( .A(n234), .B(n5418), .Z(n5417) );
  XOR U5366 ( .A(p_input[313]), .B(p_input[297]), .Z(n5418) );
  XNOR U5367 ( .A(n4998), .B(n5413), .Z(n5415) );
  XOR U5368 ( .A(n5419), .B(n5420), .Z(n4998) );
  AND U5369 ( .A(n231), .B(n5421), .Z(n5420) );
  XOR U5370 ( .A(p_input[281]), .B(p_input[265]), .Z(n5421) );
  XOR U5371 ( .A(n5422), .B(n5423), .Z(n5413) );
  AND U5372 ( .A(n5424), .B(n5425), .Z(n5423) );
  XOR U5373 ( .A(n5422), .B(n5013), .Z(n5425) );
  XNOR U5374 ( .A(p_input[296]), .B(n5426), .Z(n5013) );
  AND U5375 ( .A(n234), .B(n5427), .Z(n5426) );
  XOR U5376 ( .A(p_input[312]), .B(p_input[296]), .Z(n5427) );
  XNOR U5377 ( .A(n5010), .B(n5422), .Z(n5424) );
  XOR U5378 ( .A(n5428), .B(n5429), .Z(n5010) );
  AND U5379 ( .A(n231), .B(n5430), .Z(n5429) );
  XOR U5380 ( .A(p_input[280]), .B(p_input[264]), .Z(n5430) );
  XOR U5381 ( .A(n5431), .B(n5432), .Z(n5422) );
  AND U5382 ( .A(n5433), .B(n5434), .Z(n5432) );
  XOR U5383 ( .A(n5431), .B(n5025), .Z(n5434) );
  XNOR U5384 ( .A(p_input[295]), .B(n5435), .Z(n5025) );
  AND U5385 ( .A(n234), .B(n5436), .Z(n5435) );
  XOR U5386 ( .A(p_input[311]), .B(p_input[295]), .Z(n5436) );
  XNOR U5387 ( .A(n5022), .B(n5431), .Z(n5433) );
  XOR U5388 ( .A(n5437), .B(n5438), .Z(n5022) );
  AND U5389 ( .A(n231), .B(n5439), .Z(n5438) );
  XOR U5390 ( .A(p_input[279]), .B(p_input[263]), .Z(n5439) );
  XOR U5391 ( .A(n5440), .B(n5441), .Z(n5431) );
  AND U5392 ( .A(n5442), .B(n5443), .Z(n5441) );
  XOR U5393 ( .A(n5440), .B(n5037), .Z(n5443) );
  XNOR U5394 ( .A(p_input[294]), .B(n5444), .Z(n5037) );
  AND U5395 ( .A(n234), .B(n5445), .Z(n5444) );
  XOR U5396 ( .A(p_input[310]), .B(p_input[294]), .Z(n5445) );
  XNOR U5397 ( .A(n5034), .B(n5440), .Z(n5442) );
  XOR U5398 ( .A(n5446), .B(n5447), .Z(n5034) );
  AND U5399 ( .A(n231), .B(n5448), .Z(n5447) );
  XOR U5400 ( .A(p_input[278]), .B(p_input[262]), .Z(n5448) );
  XOR U5401 ( .A(n5449), .B(n5450), .Z(n5440) );
  AND U5402 ( .A(n5451), .B(n5452), .Z(n5450) );
  XOR U5403 ( .A(n5449), .B(n5049), .Z(n5452) );
  XNOR U5404 ( .A(p_input[293]), .B(n5453), .Z(n5049) );
  AND U5405 ( .A(n234), .B(n5454), .Z(n5453) );
  XOR U5406 ( .A(p_input[309]), .B(p_input[293]), .Z(n5454) );
  XNOR U5407 ( .A(n5046), .B(n5449), .Z(n5451) );
  XOR U5408 ( .A(n5455), .B(n5456), .Z(n5046) );
  AND U5409 ( .A(n231), .B(n5457), .Z(n5456) );
  XOR U5410 ( .A(p_input[277]), .B(p_input[261]), .Z(n5457) );
  XOR U5411 ( .A(n5458), .B(n5459), .Z(n5449) );
  AND U5412 ( .A(n5460), .B(n5461), .Z(n5459) );
  XOR U5413 ( .A(n5458), .B(n5061), .Z(n5461) );
  XNOR U5414 ( .A(p_input[292]), .B(n5462), .Z(n5061) );
  AND U5415 ( .A(n234), .B(n5463), .Z(n5462) );
  XOR U5416 ( .A(p_input[308]), .B(p_input[292]), .Z(n5463) );
  XNOR U5417 ( .A(n5058), .B(n5458), .Z(n5460) );
  XOR U5418 ( .A(n5464), .B(n5465), .Z(n5058) );
  AND U5419 ( .A(n231), .B(n5466), .Z(n5465) );
  XOR U5420 ( .A(p_input[276]), .B(p_input[260]), .Z(n5466) );
  XOR U5421 ( .A(n5467), .B(n5468), .Z(n5458) );
  AND U5422 ( .A(n5469), .B(n5470), .Z(n5468) );
  XOR U5423 ( .A(n5073), .B(n5467), .Z(n5470) );
  XNOR U5424 ( .A(p_input[291]), .B(n5471), .Z(n5073) );
  AND U5425 ( .A(n234), .B(n5472), .Z(n5471) );
  XOR U5426 ( .A(p_input[307]), .B(p_input[291]), .Z(n5472) );
  XNOR U5427 ( .A(n5467), .B(n5070), .Z(n5469) );
  XOR U5428 ( .A(n5473), .B(n5474), .Z(n5070) );
  AND U5429 ( .A(n231), .B(n5475), .Z(n5474) );
  XOR U5430 ( .A(p_input[275]), .B(p_input[259]), .Z(n5475) );
  XOR U5431 ( .A(n5476), .B(n5477), .Z(n5467) );
  AND U5432 ( .A(n5478), .B(n5479), .Z(n5477) );
  XOR U5433 ( .A(n5476), .B(n5085), .Z(n5479) );
  XNOR U5434 ( .A(p_input[290]), .B(n5480), .Z(n5085) );
  AND U5435 ( .A(n234), .B(n5481), .Z(n5480) );
  XOR U5436 ( .A(p_input[306]), .B(p_input[290]), .Z(n5481) );
  XNOR U5437 ( .A(n5082), .B(n5476), .Z(n5478) );
  XOR U5438 ( .A(n5482), .B(n5483), .Z(n5082) );
  AND U5439 ( .A(n231), .B(n5484), .Z(n5483) );
  XOR U5440 ( .A(p_input[274]), .B(p_input[258]), .Z(n5484) );
  XOR U5441 ( .A(n5485), .B(n5486), .Z(n5476) );
  AND U5442 ( .A(n5487), .B(n5488), .Z(n5486) );
  XNOR U5443 ( .A(n5489), .B(n5098), .Z(n5488) );
  XNOR U5444 ( .A(p_input[289]), .B(n5490), .Z(n5098) );
  AND U5445 ( .A(n234), .B(n5491), .Z(n5490) );
  XNOR U5446 ( .A(p_input[305]), .B(n5492), .Z(n5491) );
  IV U5447 ( .A(p_input[289]), .Z(n5492) );
  XNOR U5448 ( .A(n5095), .B(n5485), .Z(n5487) );
  XNOR U5449 ( .A(p_input[257]), .B(n5493), .Z(n5095) );
  AND U5450 ( .A(n231), .B(n5494), .Z(n5493) );
  XOR U5451 ( .A(p_input[273]), .B(p_input[257]), .Z(n5494) );
  IV U5452 ( .A(n5489), .Z(n5485) );
  AND U5453 ( .A(n5360), .B(n5363), .Z(n5489) );
  XOR U5454 ( .A(p_input[288]), .B(n5495), .Z(n5363) );
  AND U5455 ( .A(n234), .B(n5496), .Z(n5495) );
  XOR U5456 ( .A(p_input[304]), .B(p_input[288]), .Z(n5496) );
  XOR U5457 ( .A(n5497), .B(n5498), .Z(n234) );
  AND U5458 ( .A(n5499), .B(n5500), .Z(n5498) );
  XNOR U5459 ( .A(p_input[319]), .B(n5497), .Z(n5500) );
  XOR U5460 ( .A(n5497), .B(p_input[303]), .Z(n5499) );
  XOR U5461 ( .A(n5501), .B(n5502), .Z(n5497) );
  AND U5462 ( .A(n5503), .B(n5504), .Z(n5502) );
  XNOR U5463 ( .A(p_input[318]), .B(n5501), .Z(n5504) );
  XOR U5464 ( .A(n5501), .B(p_input[302]), .Z(n5503) );
  XOR U5465 ( .A(n5505), .B(n5506), .Z(n5501) );
  AND U5466 ( .A(n5507), .B(n5508), .Z(n5506) );
  XNOR U5467 ( .A(p_input[317]), .B(n5505), .Z(n5508) );
  XOR U5468 ( .A(n5505), .B(p_input[301]), .Z(n5507) );
  XOR U5469 ( .A(n5509), .B(n5510), .Z(n5505) );
  AND U5470 ( .A(n5511), .B(n5512), .Z(n5510) );
  XNOR U5471 ( .A(p_input[316]), .B(n5509), .Z(n5512) );
  XOR U5472 ( .A(n5509), .B(p_input[300]), .Z(n5511) );
  XOR U5473 ( .A(n5513), .B(n5514), .Z(n5509) );
  AND U5474 ( .A(n5515), .B(n5516), .Z(n5514) );
  XNOR U5475 ( .A(p_input[315]), .B(n5513), .Z(n5516) );
  XOR U5476 ( .A(n5513), .B(p_input[299]), .Z(n5515) );
  XOR U5477 ( .A(n5517), .B(n5518), .Z(n5513) );
  AND U5478 ( .A(n5519), .B(n5520), .Z(n5518) );
  XNOR U5479 ( .A(p_input[314]), .B(n5517), .Z(n5520) );
  XOR U5480 ( .A(n5517), .B(p_input[298]), .Z(n5519) );
  XOR U5481 ( .A(n5521), .B(n5522), .Z(n5517) );
  AND U5482 ( .A(n5523), .B(n5524), .Z(n5522) );
  XNOR U5483 ( .A(p_input[313]), .B(n5521), .Z(n5524) );
  XOR U5484 ( .A(n5521), .B(p_input[297]), .Z(n5523) );
  XOR U5485 ( .A(n5525), .B(n5526), .Z(n5521) );
  AND U5486 ( .A(n5527), .B(n5528), .Z(n5526) );
  XNOR U5487 ( .A(p_input[312]), .B(n5525), .Z(n5528) );
  XOR U5488 ( .A(n5525), .B(p_input[296]), .Z(n5527) );
  XOR U5489 ( .A(n5529), .B(n5530), .Z(n5525) );
  AND U5490 ( .A(n5531), .B(n5532), .Z(n5530) );
  XNOR U5491 ( .A(p_input[311]), .B(n5529), .Z(n5532) );
  XOR U5492 ( .A(n5529), .B(p_input[295]), .Z(n5531) );
  XOR U5493 ( .A(n5533), .B(n5534), .Z(n5529) );
  AND U5494 ( .A(n5535), .B(n5536), .Z(n5534) );
  XNOR U5495 ( .A(p_input[310]), .B(n5533), .Z(n5536) );
  XOR U5496 ( .A(n5533), .B(p_input[294]), .Z(n5535) );
  XOR U5497 ( .A(n5537), .B(n5538), .Z(n5533) );
  AND U5498 ( .A(n5539), .B(n5540), .Z(n5538) );
  XNOR U5499 ( .A(p_input[309]), .B(n5537), .Z(n5540) );
  XOR U5500 ( .A(n5537), .B(p_input[293]), .Z(n5539) );
  XOR U5501 ( .A(n5541), .B(n5542), .Z(n5537) );
  AND U5502 ( .A(n5543), .B(n5544), .Z(n5542) );
  XNOR U5503 ( .A(p_input[308]), .B(n5541), .Z(n5544) );
  XOR U5504 ( .A(n5541), .B(p_input[292]), .Z(n5543) );
  XOR U5505 ( .A(n5545), .B(n5546), .Z(n5541) );
  AND U5506 ( .A(n5547), .B(n5548), .Z(n5546) );
  XNOR U5507 ( .A(p_input[307]), .B(n5545), .Z(n5548) );
  XOR U5508 ( .A(n5545), .B(p_input[291]), .Z(n5547) );
  XOR U5509 ( .A(n5549), .B(n5550), .Z(n5545) );
  AND U5510 ( .A(n5551), .B(n5552), .Z(n5550) );
  XNOR U5511 ( .A(p_input[306]), .B(n5549), .Z(n5552) );
  XOR U5512 ( .A(n5549), .B(p_input[290]), .Z(n5551) );
  XNOR U5513 ( .A(n5553), .B(n5554), .Z(n5549) );
  AND U5514 ( .A(n5555), .B(n5556), .Z(n5554) );
  XOR U5515 ( .A(p_input[305]), .B(n5553), .Z(n5556) );
  XNOR U5516 ( .A(p_input[289]), .B(n5553), .Z(n5555) );
  AND U5517 ( .A(p_input[304]), .B(n5557), .Z(n5553) );
  IV U5518 ( .A(p_input[288]), .Z(n5557) );
  XNOR U5519 ( .A(p_input[256]), .B(n5558), .Z(n5360) );
  AND U5520 ( .A(n231), .B(n5559), .Z(n5558) );
  XOR U5521 ( .A(p_input[272]), .B(p_input[256]), .Z(n5559) );
  XOR U5522 ( .A(n5560), .B(n5561), .Z(n231) );
  AND U5523 ( .A(n5562), .B(n5563), .Z(n5561) );
  XNOR U5524 ( .A(p_input[287]), .B(n5560), .Z(n5563) );
  XOR U5525 ( .A(n5560), .B(p_input[271]), .Z(n5562) );
  XOR U5526 ( .A(n5564), .B(n5565), .Z(n5560) );
  AND U5527 ( .A(n5566), .B(n5567), .Z(n5565) );
  XNOR U5528 ( .A(p_input[286]), .B(n5564), .Z(n5567) );
  XNOR U5529 ( .A(n5564), .B(n5374), .Z(n5566) );
  IV U5530 ( .A(p_input[270]), .Z(n5374) );
  XOR U5531 ( .A(n5568), .B(n5569), .Z(n5564) );
  AND U5532 ( .A(n5570), .B(n5571), .Z(n5569) );
  XNOR U5533 ( .A(p_input[285]), .B(n5568), .Z(n5571) );
  XNOR U5534 ( .A(n5568), .B(n5383), .Z(n5570) );
  IV U5535 ( .A(p_input[269]), .Z(n5383) );
  XOR U5536 ( .A(n5572), .B(n5573), .Z(n5568) );
  AND U5537 ( .A(n5574), .B(n5575), .Z(n5573) );
  XNOR U5538 ( .A(p_input[284]), .B(n5572), .Z(n5575) );
  XNOR U5539 ( .A(n5572), .B(n5392), .Z(n5574) );
  IV U5540 ( .A(p_input[268]), .Z(n5392) );
  XOR U5541 ( .A(n5576), .B(n5577), .Z(n5572) );
  AND U5542 ( .A(n5578), .B(n5579), .Z(n5577) );
  XNOR U5543 ( .A(p_input[283]), .B(n5576), .Z(n5579) );
  XNOR U5544 ( .A(n5576), .B(n5401), .Z(n5578) );
  IV U5545 ( .A(p_input[267]), .Z(n5401) );
  XOR U5546 ( .A(n5580), .B(n5581), .Z(n5576) );
  AND U5547 ( .A(n5582), .B(n5583), .Z(n5581) );
  XNOR U5548 ( .A(p_input[282]), .B(n5580), .Z(n5583) );
  XNOR U5549 ( .A(n5580), .B(n5410), .Z(n5582) );
  IV U5550 ( .A(p_input[266]), .Z(n5410) );
  XOR U5551 ( .A(n5584), .B(n5585), .Z(n5580) );
  AND U5552 ( .A(n5586), .B(n5587), .Z(n5585) );
  XNOR U5553 ( .A(p_input[281]), .B(n5584), .Z(n5587) );
  XNOR U5554 ( .A(n5584), .B(n5419), .Z(n5586) );
  IV U5555 ( .A(p_input[265]), .Z(n5419) );
  XOR U5556 ( .A(n5588), .B(n5589), .Z(n5584) );
  AND U5557 ( .A(n5590), .B(n5591), .Z(n5589) );
  XNOR U5558 ( .A(p_input[280]), .B(n5588), .Z(n5591) );
  XNOR U5559 ( .A(n5588), .B(n5428), .Z(n5590) );
  IV U5560 ( .A(p_input[264]), .Z(n5428) );
  XOR U5561 ( .A(n5592), .B(n5593), .Z(n5588) );
  AND U5562 ( .A(n5594), .B(n5595), .Z(n5593) );
  XNOR U5563 ( .A(p_input[279]), .B(n5592), .Z(n5595) );
  XNOR U5564 ( .A(n5592), .B(n5437), .Z(n5594) );
  IV U5565 ( .A(p_input[263]), .Z(n5437) );
  XOR U5566 ( .A(n5596), .B(n5597), .Z(n5592) );
  AND U5567 ( .A(n5598), .B(n5599), .Z(n5597) );
  XNOR U5568 ( .A(p_input[278]), .B(n5596), .Z(n5599) );
  XNOR U5569 ( .A(n5596), .B(n5446), .Z(n5598) );
  IV U5570 ( .A(p_input[262]), .Z(n5446) );
  XOR U5571 ( .A(n5600), .B(n5601), .Z(n5596) );
  AND U5572 ( .A(n5602), .B(n5603), .Z(n5601) );
  XNOR U5573 ( .A(p_input[277]), .B(n5600), .Z(n5603) );
  XNOR U5574 ( .A(n5600), .B(n5455), .Z(n5602) );
  IV U5575 ( .A(p_input[261]), .Z(n5455) );
  XOR U5576 ( .A(n5604), .B(n5605), .Z(n5600) );
  AND U5577 ( .A(n5606), .B(n5607), .Z(n5605) );
  XNOR U5578 ( .A(p_input[276]), .B(n5604), .Z(n5607) );
  XNOR U5579 ( .A(n5604), .B(n5464), .Z(n5606) );
  IV U5580 ( .A(p_input[260]), .Z(n5464) );
  XOR U5581 ( .A(n5608), .B(n5609), .Z(n5604) );
  AND U5582 ( .A(n5610), .B(n5611), .Z(n5609) );
  XNOR U5583 ( .A(p_input[275]), .B(n5608), .Z(n5611) );
  XNOR U5584 ( .A(n5608), .B(n5473), .Z(n5610) );
  IV U5585 ( .A(p_input[259]), .Z(n5473) );
  XOR U5586 ( .A(n5612), .B(n5613), .Z(n5608) );
  AND U5587 ( .A(n5614), .B(n5615), .Z(n5613) );
  XNOR U5588 ( .A(p_input[274]), .B(n5612), .Z(n5615) );
  XNOR U5589 ( .A(n5612), .B(n5482), .Z(n5614) );
  IV U5590 ( .A(p_input[258]), .Z(n5482) );
  XNOR U5591 ( .A(n5616), .B(n5617), .Z(n5612) );
  AND U5592 ( .A(n5618), .B(n5619), .Z(n5617) );
  XOR U5593 ( .A(p_input[273]), .B(n5616), .Z(n5619) );
  XNOR U5594 ( .A(p_input[257]), .B(n5616), .Z(n5618) );
  AND U5595 ( .A(p_input[272]), .B(n5620), .Z(n5616) );
  IV U5596 ( .A(p_input[256]), .Z(n5620) );
  XOR U5597 ( .A(n5621), .B(n5622), .Z(n3848) );
  AND U5598 ( .A(n287), .B(n5623), .Z(n5622) );
  XNOR U5599 ( .A(n5624), .B(n5621), .Z(n5623) );
  XOR U5600 ( .A(n5625), .B(n5626), .Z(n287) );
  AND U5601 ( .A(n5627), .B(n5628), .Z(n5626) );
  XNOR U5602 ( .A(n3863), .B(n5625), .Z(n5628) );
  AND U5603 ( .A(n5629), .B(n5630), .Z(n3863) );
  XNOR U5604 ( .A(n5625), .B(n3860), .Z(n5627) );
  IV U5605 ( .A(n5631), .Z(n3860) );
  AND U5606 ( .A(n5632), .B(n5633), .Z(n5631) );
  XOR U5607 ( .A(n5634), .B(n5635), .Z(n5625) );
  AND U5608 ( .A(n5636), .B(n5637), .Z(n5635) );
  XOR U5609 ( .A(n5634), .B(n3875), .Z(n5637) );
  XOR U5610 ( .A(n5638), .B(n5639), .Z(n3875) );
  AND U5611 ( .A(n262), .B(n5640), .Z(n5639) );
  XOR U5612 ( .A(n5641), .B(n5638), .Z(n5640) );
  XNOR U5613 ( .A(n3872), .B(n5634), .Z(n5636) );
  XOR U5614 ( .A(n5642), .B(n5643), .Z(n3872) );
  AND U5615 ( .A(n259), .B(n5644), .Z(n5643) );
  XOR U5616 ( .A(n5645), .B(n5642), .Z(n5644) );
  XOR U5617 ( .A(n5646), .B(n5647), .Z(n5634) );
  AND U5618 ( .A(n5648), .B(n5649), .Z(n5647) );
  XOR U5619 ( .A(n5646), .B(n3887), .Z(n5649) );
  XOR U5620 ( .A(n5650), .B(n5651), .Z(n3887) );
  AND U5621 ( .A(n262), .B(n5652), .Z(n5651) );
  XOR U5622 ( .A(n5653), .B(n5650), .Z(n5652) );
  XNOR U5623 ( .A(n3884), .B(n5646), .Z(n5648) );
  XOR U5624 ( .A(n5654), .B(n5655), .Z(n3884) );
  AND U5625 ( .A(n259), .B(n5656), .Z(n5655) );
  XOR U5626 ( .A(n5657), .B(n5654), .Z(n5656) );
  XOR U5627 ( .A(n5658), .B(n5659), .Z(n5646) );
  AND U5628 ( .A(n5660), .B(n5661), .Z(n5659) );
  XOR U5629 ( .A(n5658), .B(n3899), .Z(n5661) );
  XOR U5630 ( .A(n5662), .B(n5663), .Z(n3899) );
  AND U5631 ( .A(n262), .B(n5664), .Z(n5663) );
  XOR U5632 ( .A(n5665), .B(n5662), .Z(n5664) );
  XNOR U5633 ( .A(n3896), .B(n5658), .Z(n5660) );
  XOR U5634 ( .A(n5666), .B(n5667), .Z(n3896) );
  AND U5635 ( .A(n259), .B(n5668), .Z(n5667) );
  XOR U5636 ( .A(n5669), .B(n5666), .Z(n5668) );
  XOR U5637 ( .A(n5670), .B(n5671), .Z(n5658) );
  AND U5638 ( .A(n5672), .B(n5673), .Z(n5671) );
  XOR U5639 ( .A(n5670), .B(n3911), .Z(n5673) );
  XOR U5640 ( .A(n5674), .B(n5675), .Z(n3911) );
  AND U5641 ( .A(n262), .B(n5676), .Z(n5675) );
  XOR U5642 ( .A(n5677), .B(n5674), .Z(n5676) );
  XNOR U5643 ( .A(n3908), .B(n5670), .Z(n5672) );
  XOR U5644 ( .A(n5678), .B(n5679), .Z(n3908) );
  AND U5645 ( .A(n259), .B(n5680), .Z(n5679) );
  XOR U5646 ( .A(n5681), .B(n5678), .Z(n5680) );
  XOR U5647 ( .A(n5682), .B(n5683), .Z(n5670) );
  AND U5648 ( .A(n5684), .B(n5685), .Z(n5683) );
  XOR U5649 ( .A(n5682), .B(n3923), .Z(n5685) );
  XOR U5650 ( .A(n5686), .B(n5687), .Z(n3923) );
  AND U5651 ( .A(n262), .B(n5688), .Z(n5687) );
  XOR U5652 ( .A(n5689), .B(n5686), .Z(n5688) );
  XNOR U5653 ( .A(n3920), .B(n5682), .Z(n5684) );
  XOR U5654 ( .A(n5690), .B(n5691), .Z(n3920) );
  AND U5655 ( .A(n259), .B(n5692), .Z(n5691) );
  XOR U5656 ( .A(n5693), .B(n5690), .Z(n5692) );
  XOR U5657 ( .A(n5694), .B(n5695), .Z(n5682) );
  AND U5658 ( .A(n5696), .B(n5697), .Z(n5695) );
  XOR U5659 ( .A(n5694), .B(n3935), .Z(n5697) );
  XOR U5660 ( .A(n5698), .B(n5699), .Z(n3935) );
  AND U5661 ( .A(n262), .B(n5700), .Z(n5699) );
  XOR U5662 ( .A(n5701), .B(n5698), .Z(n5700) );
  XNOR U5663 ( .A(n3932), .B(n5694), .Z(n5696) );
  XOR U5664 ( .A(n5702), .B(n5703), .Z(n3932) );
  AND U5665 ( .A(n259), .B(n5704), .Z(n5703) );
  XOR U5666 ( .A(n5705), .B(n5702), .Z(n5704) );
  XOR U5667 ( .A(n5706), .B(n5707), .Z(n5694) );
  AND U5668 ( .A(n5708), .B(n5709), .Z(n5707) );
  XOR U5669 ( .A(n5706), .B(n3947), .Z(n5709) );
  XOR U5670 ( .A(n5710), .B(n5711), .Z(n3947) );
  AND U5671 ( .A(n262), .B(n5712), .Z(n5711) );
  XOR U5672 ( .A(n5713), .B(n5710), .Z(n5712) );
  XNOR U5673 ( .A(n3944), .B(n5706), .Z(n5708) );
  XOR U5674 ( .A(n5714), .B(n5715), .Z(n3944) );
  AND U5675 ( .A(n259), .B(n5716), .Z(n5715) );
  XOR U5676 ( .A(n5717), .B(n5714), .Z(n5716) );
  XOR U5677 ( .A(n5718), .B(n5719), .Z(n5706) );
  AND U5678 ( .A(n5720), .B(n5721), .Z(n5719) );
  XOR U5679 ( .A(n5718), .B(n3959), .Z(n5721) );
  XOR U5680 ( .A(n5722), .B(n5723), .Z(n3959) );
  AND U5681 ( .A(n262), .B(n5724), .Z(n5723) );
  XOR U5682 ( .A(n5725), .B(n5722), .Z(n5724) );
  XNOR U5683 ( .A(n3956), .B(n5718), .Z(n5720) );
  XOR U5684 ( .A(n5726), .B(n5727), .Z(n3956) );
  AND U5685 ( .A(n259), .B(n5728), .Z(n5727) );
  XOR U5686 ( .A(n5729), .B(n5726), .Z(n5728) );
  XOR U5687 ( .A(n5730), .B(n5731), .Z(n5718) );
  AND U5688 ( .A(n5732), .B(n5733), .Z(n5731) );
  XOR U5689 ( .A(n5730), .B(n3971), .Z(n5733) );
  XOR U5690 ( .A(n5734), .B(n5735), .Z(n3971) );
  AND U5691 ( .A(n262), .B(n5736), .Z(n5735) );
  XOR U5692 ( .A(n5737), .B(n5734), .Z(n5736) );
  XNOR U5693 ( .A(n3968), .B(n5730), .Z(n5732) );
  XOR U5694 ( .A(n5738), .B(n5739), .Z(n3968) );
  AND U5695 ( .A(n259), .B(n5740), .Z(n5739) );
  XOR U5696 ( .A(n5741), .B(n5738), .Z(n5740) );
  XOR U5697 ( .A(n5742), .B(n5743), .Z(n5730) );
  AND U5698 ( .A(n5744), .B(n5745), .Z(n5743) );
  XOR U5699 ( .A(n5742), .B(n3983), .Z(n5745) );
  XOR U5700 ( .A(n5746), .B(n5747), .Z(n3983) );
  AND U5701 ( .A(n262), .B(n5748), .Z(n5747) );
  XOR U5702 ( .A(n5749), .B(n5746), .Z(n5748) );
  XNOR U5703 ( .A(n3980), .B(n5742), .Z(n5744) );
  XOR U5704 ( .A(n5750), .B(n5751), .Z(n3980) );
  AND U5705 ( .A(n259), .B(n5752), .Z(n5751) );
  XOR U5706 ( .A(n5753), .B(n5750), .Z(n5752) );
  XOR U5707 ( .A(n5754), .B(n5755), .Z(n5742) );
  AND U5708 ( .A(n5756), .B(n5757), .Z(n5755) );
  XOR U5709 ( .A(n5754), .B(n3995), .Z(n5757) );
  XOR U5710 ( .A(n5758), .B(n5759), .Z(n3995) );
  AND U5711 ( .A(n262), .B(n5760), .Z(n5759) );
  XOR U5712 ( .A(n5761), .B(n5758), .Z(n5760) );
  XNOR U5713 ( .A(n3992), .B(n5754), .Z(n5756) );
  XOR U5714 ( .A(n5762), .B(n5763), .Z(n3992) );
  AND U5715 ( .A(n259), .B(n5764), .Z(n5763) );
  XOR U5716 ( .A(n5765), .B(n5762), .Z(n5764) );
  XOR U5717 ( .A(n5766), .B(n5767), .Z(n5754) );
  AND U5718 ( .A(n5768), .B(n5769), .Z(n5767) );
  XOR U5719 ( .A(n4007), .B(n5766), .Z(n5769) );
  XOR U5720 ( .A(n5770), .B(n5771), .Z(n4007) );
  AND U5721 ( .A(n262), .B(n5772), .Z(n5771) );
  XOR U5722 ( .A(n5770), .B(n5773), .Z(n5772) );
  XNOR U5723 ( .A(n5766), .B(n4004), .Z(n5768) );
  XOR U5724 ( .A(n5774), .B(n5775), .Z(n4004) );
  AND U5725 ( .A(n259), .B(n5776), .Z(n5775) );
  XOR U5726 ( .A(n5774), .B(n5777), .Z(n5776) );
  XOR U5727 ( .A(n5778), .B(n5779), .Z(n5766) );
  AND U5728 ( .A(n5780), .B(n5781), .Z(n5779) );
  XOR U5729 ( .A(n5778), .B(n4019), .Z(n5781) );
  XOR U5730 ( .A(n5782), .B(n5783), .Z(n4019) );
  AND U5731 ( .A(n262), .B(n5784), .Z(n5783) );
  XOR U5732 ( .A(n5785), .B(n5782), .Z(n5784) );
  XNOR U5733 ( .A(n4016), .B(n5778), .Z(n5780) );
  XOR U5734 ( .A(n5786), .B(n5787), .Z(n4016) );
  AND U5735 ( .A(n259), .B(n5788), .Z(n5787) );
  XOR U5736 ( .A(n5789), .B(n5786), .Z(n5788) );
  XOR U5737 ( .A(n5790), .B(n5791), .Z(n5778) );
  AND U5738 ( .A(n5792), .B(n5793), .Z(n5791) );
  XNOR U5739 ( .A(n5794), .B(n4032), .Z(n5793) );
  XOR U5740 ( .A(n5795), .B(n5796), .Z(n4032) );
  AND U5741 ( .A(n262), .B(n5797), .Z(n5796) );
  XOR U5742 ( .A(n5798), .B(n5795), .Z(n5797) );
  XNOR U5743 ( .A(n4029), .B(n5790), .Z(n5792) );
  XOR U5744 ( .A(n5799), .B(n5800), .Z(n4029) );
  AND U5745 ( .A(n259), .B(n5801), .Z(n5800) );
  XOR U5746 ( .A(n5802), .B(n5799), .Z(n5801) );
  IV U5747 ( .A(n5794), .Z(n5790) );
  AND U5748 ( .A(n5621), .B(n5624), .Z(n5794) );
  XNOR U5749 ( .A(n5803), .B(n5804), .Z(n5624) );
  AND U5750 ( .A(n262), .B(n5805), .Z(n5804) );
  XNOR U5751 ( .A(n5806), .B(n5803), .Z(n5805) );
  XOR U5752 ( .A(n5807), .B(n5808), .Z(n262) );
  AND U5753 ( .A(n5809), .B(n5810), .Z(n5808) );
  XNOR U5754 ( .A(n5629), .B(n5807), .Z(n5810) );
  AND U5755 ( .A(n5811), .B(n5812), .Z(n5629) );
  XOR U5756 ( .A(n5807), .B(n5630), .Z(n5809) );
  AND U5757 ( .A(n5813), .B(n5814), .Z(n5630) );
  XOR U5758 ( .A(n5815), .B(n5816), .Z(n5807) );
  AND U5759 ( .A(n5817), .B(n5818), .Z(n5816) );
  XOR U5760 ( .A(n5815), .B(n5641), .Z(n5818) );
  XOR U5761 ( .A(n5819), .B(n5820), .Z(n5641) );
  AND U5762 ( .A(n198), .B(n5821), .Z(n5820) );
  XOR U5763 ( .A(n5822), .B(n5819), .Z(n5821) );
  XNOR U5764 ( .A(n5638), .B(n5815), .Z(n5817) );
  XOR U5765 ( .A(n5823), .B(n5824), .Z(n5638) );
  AND U5766 ( .A(n196), .B(n5825), .Z(n5824) );
  XOR U5767 ( .A(n5826), .B(n5823), .Z(n5825) );
  XOR U5768 ( .A(n5827), .B(n5828), .Z(n5815) );
  AND U5769 ( .A(n5829), .B(n5830), .Z(n5828) );
  XOR U5770 ( .A(n5827), .B(n5653), .Z(n5830) );
  XOR U5771 ( .A(n5831), .B(n5832), .Z(n5653) );
  AND U5772 ( .A(n198), .B(n5833), .Z(n5832) );
  XOR U5773 ( .A(n5834), .B(n5831), .Z(n5833) );
  XNOR U5774 ( .A(n5650), .B(n5827), .Z(n5829) );
  XOR U5775 ( .A(n5835), .B(n5836), .Z(n5650) );
  AND U5776 ( .A(n196), .B(n5837), .Z(n5836) );
  XOR U5777 ( .A(n5838), .B(n5835), .Z(n5837) );
  XOR U5778 ( .A(n5839), .B(n5840), .Z(n5827) );
  AND U5779 ( .A(n5841), .B(n5842), .Z(n5840) );
  XOR U5780 ( .A(n5839), .B(n5665), .Z(n5842) );
  XOR U5781 ( .A(n5843), .B(n5844), .Z(n5665) );
  AND U5782 ( .A(n198), .B(n5845), .Z(n5844) );
  XOR U5783 ( .A(n5846), .B(n5843), .Z(n5845) );
  XNOR U5784 ( .A(n5662), .B(n5839), .Z(n5841) );
  XOR U5785 ( .A(n5847), .B(n5848), .Z(n5662) );
  AND U5786 ( .A(n196), .B(n5849), .Z(n5848) );
  XOR U5787 ( .A(n5850), .B(n5847), .Z(n5849) );
  XOR U5788 ( .A(n5851), .B(n5852), .Z(n5839) );
  AND U5789 ( .A(n5853), .B(n5854), .Z(n5852) );
  XOR U5790 ( .A(n5851), .B(n5677), .Z(n5854) );
  XOR U5791 ( .A(n5855), .B(n5856), .Z(n5677) );
  AND U5792 ( .A(n198), .B(n5857), .Z(n5856) );
  XOR U5793 ( .A(n5858), .B(n5855), .Z(n5857) );
  XNOR U5794 ( .A(n5674), .B(n5851), .Z(n5853) );
  XOR U5795 ( .A(n5859), .B(n5860), .Z(n5674) );
  AND U5796 ( .A(n196), .B(n5861), .Z(n5860) );
  XOR U5797 ( .A(n5862), .B(n5859), .Z(n5861) );
  XOR U5798 ( .A(n5863), .B(n5864), .Z(n5851) );
  AND U5799 ( .A(n5865), .B(n5866), .Z(n5864) );
  XOR U5800 ( .A(n5863), .B(n5689), .Z(n5866) );
  XOR U5801 ( .A(n5867), .B(n5868), .Z(n5689) );
  AND U5802 ( .A(n198), .B(n5869), .Z(n5868) );
  XOR U5803 ( .A(n5870), .B(n5867), .Z(n5869) );
  XNOR U5804 ( .A(n5686), .B(n5863), .Z(n5865) );
  XOR U5805 ( .A(n5871), .B(n5872), .Z(n5686) );
  AND U5806 ( .A(n196), .B(n5873), .Z(n5872) );
  XOR U5807 ( .A(n5874), .B(n5871), .Z(n5873) );
  XOR U5808 ( .A(n5875), .B(n5876), .Z(n5863) );
  AND U5809 ( .A(n5877), .B(n5878), .Z(n5876) );
  XOR U5810 ( .A(n5875), .B(n5701), .Z(n5878) );
  XOR U5811 ( .A(n5879), .B(n5880), .Z(n5701) );
  AND U5812 ( .A(n198), .B(n5881), .Z(n5880) );
  XOR U5813 ( .A(n5882), .B(n5879), .Z(n5881) );
  XNOR U5814 ( .A(n5698), .B(n5875), .Z(n5877) );
  XOR U5815 ( .A(n5883), .B(n5884), .Z(n5698) );
  AND U5816 ( .A(n196), .B(n5885), .Z(n5884) );
  XOR U5817 ( .A(n5886), .B(n5883), .Z(n5885) );
  XOR U5818 ( .A(n5887), .B(n5888), .Z(n5875) );
  AND U5819 ( .A(n5889), .B(n5890), .Z(n5888) );
  XOR U5820 ( .A(n5887), .B(n5713), .Z(n5890) );
  XOR U5821 ( .A(n5891), .B(n5892), .Z(n5713) );
  AND U5822 ( .A(n198), .B(n5893), .Z(n5892) );
  XOR U5823 ( .A(n5894), .B(n5891), .Z(n5893) );
  XNOR U5824 ( .A(n5710), .B(n5887), .Z(n5889) );
  XOR U5825 ( .A(n5895), .B(n5896), .Z(n5710) );
  AND U5826 ( .A(n196), .B(n5897), .Z(n5896) );
  XOR U5827 ( .A(n5898), .B(n5895), .Z(n5897) );
  XOR U5828 ( .A(n5899), .B(n5900), .Z(n5887) );
  AND U5829 ( .A(n5901), .B(n5902), .Z(n5900) );
  XOR U5830 ( .A(n5899), .B(n5725), .Z(n5902) );
  XOR U5831 ( .A(n5903), .B(n5904), .Z(n5725) );
  AND U5832 ( .A(n198), .B(n5905), .Z(n5904) );
  XOR U5833 ( .A(n5906), .B(n5903), .Z(n5905) );
  XNOR U5834 ( .A(n5722), .B(n5899), .Z(n5901) );
  XOR U5835 ( .A(n5907), .B(n5908), .Z(n5722) );
  AND U5836 ( .A(n196), .B(n5909), .Z(n5908) );
  XOR U5837 ( .A(n5910), .B(n5907), .Z(n5909) );
  XOR U5838 ( .A(n5911), .B(n5912), .Z(n5899) );
  AND U5839 ( .A(n5913), .B(n5914), .Z(n5912) );
  XOR U5840 ( .A(n5911), .B(n5737), .Z(n5914) );
  XOR U5841 ( .A(n5915), .B(n5916), .Z(n5737) );
  AND U5842 ( .A(n198), .B(n5917), .Z(n5916) );
  XOR U5843 ( .A(n5918), .B(n5915), .Z(n5917) );
  XNOR U5844 ( .A(n5734), .B(n5911), .Z(n5913) );
  XOR U5845 ( .A(n5919), .B(n5920), .Z(n5734) );
  AND U5846 ( .A(n196), .B(n5921), .Z(n5920) );
  XOR U5847 ( .A(n5922), .B(n5919), .Z(n5921) );
  XOR U5848 ( .A(n5923), .B(n5924), .Z(n5911) );
  AND U5849 ( .A(n5925), .B(n5926), .Z(n5924) );
  XOR U5850 ( .A(n5923), .B(n5749), .Z(n5926) );
  XOR U5851 ( .A(n5927), .B(n5928), .Z(n5749) );
  AND U5852 ( .A(n198), .B(n5929), .Z(n5928) );
  XOR U5853 ( .A(n5930), .B(n5927), .Z(n5929) );
  XNOR U5854 ( .A(n5746), .B(n5923), .Z(n5925) );
  XOR U5855 ( .A(n5931), .B(n5932), .Z(n5746) );
  AND U5856 ( .A(n196), .B(n5933), .Z(n5932) );
  XOR U5857 ( .A(n5934), .B(n5931), .Z(n5933) );
  XOR U5858 ( .A(n5935), .B(n5936), .Z(n5923) );
  AND U5859 ( .A(n5937), .B(n5938), .Z(n5936) );
  XOR U5860 ( .A(n5935), .B(n5761), .Z(n5938) );
  XOR U5861 ( .A(n5939), .B(n5940), .Z(n5761) );
  AND U5862 ( .A(n198), .B(n5941), .Z(n5940) );
  XOR U5863 ( .A(n5942), .B(n5939), .Z(n5941) );
  XNOR U5864 ( .A(n5758), .B(n5935), .Z(n5937) );
  XOR U5865 ( .A(n5943), .B(n5944), .Z(n5758) );
  AND U5866 ( .A(n196), .B(n5945), .Z(n5944) );
  XOR U5867 ( .A(n5946), .B(n5943), .Z(n5945) );
  XOR U5868 ( .A(n5947), .B(n5948), .Z(n5935) );
  AND U5869 ( .A(n5949), .B(n5950), .Z(n5948) );
  XOR U5870 ( .A(n5773), .B(n5947), .Z(n5950) );
  XOR U5871 ( .A(n5951), .B(n5952), .Z(n5773) );
  AND U5872 ( .A(n198), .B(n5953), .Z(n5952) );
  XOR U5873 ( .A(n5951), .B(n5954), .Z(n5953) );
  XNOR U5874 ( .A(n5947), .B(n5770), .Z(n5949) );
  XOR U5875 ( .A(n5955), .B(n5956), .Z(n5770) );
  AND U5876 ( .A(n196), .B(n5957), .Z(n5956) );
  XOR U5877 ( .A(n5955), .B(n5958), .Z(n5957) );
  XOR U5878 ( .A(n5959), .B(n5960), .Z(n5947) );
  AND U5879 ( .A(n5961), .B(n5962), .Z(n5960) );
  XOR U5880 ( .A(n5959), .B(n5785), .Z(n5962) );
  XOR U5881 ( .A(n5963), .B(n5964), .Z(n5785) );
  AND U5882 ( .A(n198), .B(n5965), .Z(n5964) );
  XOR U5883 ( .A(n5966), .B(n5963), .Z(n5965) );
  XNOR U5884 ( .A(n5782), .B(n5959), .Z(n5961) );
  XOR U5885 ( .A(n5967), .B(n5968), .Z(n5782) );
  AND U5886 ( .A(n196), .B(n5969), .Z(n5968) );
  XOR U5887 ( .A(n5970), .B(n5967), .Z(n5969) );
  XOR U5888 ( .A(n5971), .B(n5972), .Z(n5959) );
  AND U5889 ( .A(n5973), .B(n5974), .Z(n5972) );
  XNOR U5890 ( .A(n5975), .B(n5798), .Z(n5974) );
  XOR U5891 ( .A(n5976), .B(n5977), .Z(n5798) );
  AND U5892 ( .A(n198), .B(n5978), .Z(n5977) );
  XOR U5893 ( .A(n5979), .B(n5976), .Z(n5978) );
  XNOR U5894 ( .A(n5795), .B(n5971), .Z(n5973) );
  XOR U5895 ( .A(n5980), .B(n5981), .Z(n5795) );
  AND U5896 ( .A(n196), .B(n5982), .Z(n5981) );
  XOR U5897 ( .A(n5983), .B(n5980), .Z(n5982) );
  IV U5898 ( .A(n5975), .Z(n5971) );
  AND U5899 ( .A(n5803), .B(n5806), .Z(n5975) );
  XNOR U5900 ( .A(n5984), .B(n5985), .Z(n5806) );
  AND U5901 ( .A(n198), .B(n5986), .Z(n5985) );
  XNOR U5902 ( .A(n5987), .B(n5984), .Z(n5986) );
  XOR U5903 ( .A(n5988), .B(n5989), .Z(n198) );
  AND U5904 ( .A(n5990), .B(n5991), .Z(n5989) );
  XNOR U5905 ( .A(n5811), .B(n5988), .Z(n5991) );
  AND U5906 ( .A(p_input[255]), .B(p_input[239]), .Z(n5811) );
  XOR U5907 ( .A(n5988), .B(n5812), .Z(n5990) );
  AND U5908 ( .A(p_input[223]), .B(p_input[207]), .Z(n5812) );
  XOR U5909 ( .A(n5992), .B(n5993), .Z(n5988) );
  AND U5910 ( .A(n5994), .B(n5995), .Z(n5993) );
  XOR U5911 ( .A(n5992), .B(n5822), .Z(n5995) );
  XNOR U5912 ( .A(p_input[238]), .B(n5996), .Z(n5822) );
  AND U5913 ( .A(n274), .B(n5997), .Z(n5996) );
  XOR U5914 ( .A(p_input[254]), .B(p_input[238]), .Z(n5997) );
  XNOR U5915 ( .A(n5819), .B(n5992), .Z(n5994) );
  XOR U5916 ( .A(n5998), .B(n5999), .Z(n5819) );
  AND U5917 ( .A(n272), .B(n6000), .Z(n5999) );
  XOR U5918 ( .A(p_input[222]), .B(p_input[206]), .Z(n6000) );
  XOR U5919 ( .A(n6001), .B(n6002), .Z(n5992) );
  AND U5920 ( .A(n6003), .B(n6004), .Z(n6002) );
  XOR U5921 ( .A(n6001), .B(n5834), .Z(n6004) );
  XNOR U5922 ( .A(p_input[237]), .B(n6005), .Z(n5834) );
  AND U5923 ( .A(n274), .B(n6006), .Z(n6005) );
  XOR U5924 ( .A(p_input[253]), .B(p_input[237]), .Z(n6006) );
  XNOR U5925 ( .A(n5831), .B(n6001), .Z(n6003) );
  XOR U5926 ( .A(n6007), .B(n6008), .Z(n5831) );
  AND U5927 ( .A(n272), .B(n6009), .Z(n6008) );
  XOR U5928 ( .A(p_input[221]), .B(p_input[205]), .Z(n6009) );
  XOR U5929 ( .A(n6010), .B(n6011), .Z(n6001) );
  AND U5930 ( .A(n6012), .B(n6013), .Z(n6011) );
  XOR U5931 ( .A(n6010), .B(n5846), .Z(n6013) );
  XNOR U5932 ( .A(p_input[236]), .B(n6014), .Z(n5846) );
  AND U5933 ( .A(n274), .B(n6015), .Z(n6014) );
  XOR U5934 ( .A(p_input[252]), .B(p_input[236]), .Z(n6015) );
  XNOR U5935 ( .A(n5843), .B(n6010), .Z(n6012) );
  XOR U5936 ( .A(n6016), .B(n6017), .Z(n5843) );
  AND U5937 ( .A(n272), .B(n6018), .Z(n6017) );
  XOR U5938 ( .A(p_input[220]), .B(p_input[204]), .Z(n6018) );
  XOR U5939 ( .A(n6019), .B(n6020), .Z(n6010) );
  AND U5940 ( .A(n6021), .B(n6022), .Z(n6020) );
  XOR U5941 ( .A(n6019), .B(n5858), .Z(n6022) );
  XNOR U5942 ( .A(p_input[235]), .B(n6023), .Z(n5858) );
  AND U5943 ( .A(n274), .B(n6024), .Z(n6023) );
  XOR U5944 ( .A(p_input[251]), .B(p_input[235]), .Z(n6024) );
  XNOR U5945 ( .A(n5855), .B(n6019), .Z(n6021) );
  XOR U5946 ( .A(n6025), .B(n6026), .Z(n5855) );
  AND U5947 ( .A(n272), .B(n6027), .Z(n6026) );
  XOR U5948 ( .A(p_input[219]), .B(p_input[203]), .Z(n6027) );
  XOR U5949 ( .A(n6028), .B(n6029), .Z(n6019) );
  AND U5950 ( .A(n6030), .B(n6031), .Z(n6029) );
  XOR U5951 ( .A(n6028), .B(n5870), .Z(n6031) );
  XNOR U5952 ( .A(p_input[234]), .B(n6032), .Z(n5870) );
  AND U5953 ( .A(n274), .B(n6033), .Z(n6032) );
  XOR U5954 ( .A(p_input[250]), .B(p_input[234]), .Z(n6033) );
  XNOR U5955 ( .A(n5867), .B(n6028), .Z(n6030) );
  XOR U5956 ( .A(n6034), .B(n6035), .Z(n5867) );
  AND U5957 ( .A(n272), .B(n6036), .Z(n6035) );
  XOR U5958 ( .A(p_input[218]), .B(p_input[202]), .Z(n6036) );
  XOR U5959 ( .A(n6037), .B(n6038), .Z(n6028) );
  AND U5960 ( .A(n6039), .B(n6040), .Z(n6038) );
  XOR U5961 ( .A(n6037), .B(n5882), .Z(n6040) );
  XNOR U5962 ( .A(p_input[233]), .B(n6041), .Z(n5882) );
  AND U5963 ( .A(n274), .B(n6042), .Z(n6041) );
  XOR U5964 ( .A(p_input[249]), .B(p_input[233]), .Z(n6042) );
  XNOR U5965 ( .A(n5879), .B(n6037), .Z(n6039) );
  XOR U5966 ( .A(n6043), .B(n6044), .Z(n5879) );
  AND U5967 ( .A(n272), .B(n6045), .Z(n6044) );
  XOR U5968 ( .A(p_input[217]), .B(p_input[201]), .Z(n6045) );
  XOR U5969 ( .A(n6046), .B(n6047), .Z(n6037) );
  AND U5970 ( .A(n6048), .B(n6049), .Z(n6047) );
  XOR U5971 ( .A(n6046), .B(n5894), .Z(n6049) );
  XNOR U5972 ( .A(p_input[232]), .B(n6050), .Z(n5894) );
  AND U5973 ( .A(n274), .B(n6051), .Z(n6050) );
  XOR U5974 ( .A(p_input[248]), .B(p_input[232]), .Z(n6051) );
  XNOR U5975 ( .A(n5891), .B(n6046), .Z(n6048) );
  XOR U5976 ( .A(n6052), .B(n6053), .Z(n5891) );
  AND U5977 ( .A(n272), .B(n6054), .Z(n6053) );
  XOR U5978 ( .A(p_input[216]), .B(p_input[200]), .Z(n6054) );
  XOR U5979 ( .A(n6055), .B(n6056), .Z(n6046) );
  AND U5980 ( .A(n6057), .B(n6058), .Z(n6056) );
  XOR U5981 ( .A(n6055), .B(n5906), .Z(n6058) );
  XNOR U5982 ( .A(p_input[231]), .B(n6059), .Z(n5906) );
  AND U5983 ( .A(n274), .B(n6060), .Z(n6059) );
  XOR U5984 ( .A(p_input[247]), .B(p_input[231]), .Z(n6060) );
  XNOR U5985 ( .A(n5903), .B(n6055), .Z(n6057) );
  XOR U5986 ( .A(n6061), .B(n6062), .Z(n5903) );
  AND U5987 ( .A(n272), .B(n6063), .Z(n6062) );
  XOR U5988 ( .A(p_input[215]), .B(p_input[199]), .Z(n6063) );
  XOR U5989 ( .A(n6064), .B(n6065), .Z(n6055) );
  AND U5990 ( .A(n6066), .B(n6067), .Z(n6065) );
  XOR U5991 ( .A(n6064), .B(n5918), .Z(n6067) );
  XNOR U5992 ( .A(p_input[230]), .B(n6068), .Z(n5918) );
  AND U5993 ( .A(n274), .B(n6069), .Z(n6068) );
  XOR U5994 ( .A(p_input[246]), .B(p_input[230]), .Z(n6069) );
  XNOR U5995 ( .A(n5915), .B(n6064), .Z(n6066) );
  XOR U5996 ( .A(n6070), .B(n6071), .Z(n5915) );
  AND U5997 ( .A(n272), .B(n6072), .Z(n6071) );
  XOR U5998 ( .A(p_input[214]), .B(p_input[198]), .Z(n6072) );
  XOR U5999 ( .A(n6073), .B(n6074), .Z(n6064) );
  AND U6000 ( .A(n6075), .B(n6076), .Z(n6074) );
  XOR U6001 ( .A(n6073), .B(n5930), .Z(n6076) );
  XNOR U6002 ( .A(p_input[229]), .B(n6077), .Z(n5930) );
  AND U6003 ( .A(n274), .B(n6078), .Z(n6077) );
  XOR U6004 ( .A(p_input[245]), .B(p_input[229]), .Z(n6078) );
  XNOR U6005 ( .A(n5927), .B(n6073), .Z(n6075) );
  XOR U6006 ( .A(n6079), .B(n6080), .Z(n5927) );
  AND U6007 ( .A(n272), .B(n6081), .Z(n6080) );
  XOR U6008 ( .A(p_input[213]), .B(p_input[197]), .Z(n6081) );
  XOR U6009 ( .A(n6082), .B(n6083), .Z(n6073) );
  AND U6010 ( .A(n6084), .B(n6085), .Z(n6083) );
  XOR U6011 ( .A(n6082), .B(n5942), .Z(n6085) );
  XNOR U6012 ( .A(p_input[228]), .B(n6086), .Z(n5942) );
  AND U6013 ( .A(n274), .B(n6087), .Z(n6086) );
  XOR U6014 ( .A(p_input[244]), .B(p_input[228]), .Z(n6087) );
  XNOR U6015 ( .A(n5939), .B(n6082), .Z(n6084) );
  XOR U6016 ( .A(n6088), .B(n6089), .Z(n5939) );
  AND U6017 ( .A(n272), .B(n6090), .Z(n6089) );
  XOR U6018 ( .A(p_input[212]), .B(p_input[196]), .Z(n6090) );
  XOR U6019 ( .A(n6091), .B(n6092), .Z(n6082) );
  AND U6020 ( .A(n6093), .B(n6094), .Z(n6092) );
  XOR U6021 ( .A(n5954), .B(n6091), .Z(n6094) );
  XNOR U6022 ( .A(p_input[227]), .B(n6095), .Z(n5954) );
  AND U6023 ( .A(n274), .B(n6096), .Z(n6095) );
  XOR U6024 ( .A(p_input[243]), .B(p_input[227]), .Z(n6096) );
  XNOR U6025 ( .A(n6091), .B(n5951), .Z(n6093) );
  XOR U6026 ( .A(n6097), .B(n6098), .Z(n5951) );
  AND U6027 ( .A(n272), .B(n6099), .Z(n6098) );
  XOR U6028 ( .A(p_input[211]), .B(p_input[195]), .Z(n6099) );
  XOR U6029 ( .A(n6100), .B(n6101), .Z(n6091) );
  AND U6030 ( .A(n6102), .B(n6103), .Z(n6101) );
  XOR U6031 ( .A(n6100), .B(n5966), .Z(n6103) );
  XNOR U6032 ( .A(p_input[226]), .B(n6104), .Z(n5966) );
  AND U6033 ( .A(n274), .B(n6105), .Z(n6104) );
  XOR U6034 ( .A(p_input[242]), .B(p_input[226]), .Z(n6105) );
  XNOR U6035 ( .A(n5963), .B(n6100), .Z(n6102) );
  XOR U6036 ( .A(n6106), .B(n6107), .Z(n5963) );
  AND U6037 ( .A(n272), .B(n6108), .Z(n6107) );
  XOR U6038 ( .A(p_input[210]), .B(p_input[194]), .Z(n6108) );
  XOR U6039 ( .A(n6109), .B(n6110), .Z(n6100) );
  AND U6040 ( .A(n6111), .B(n6112), .Z(n6110) );
  XNOR U6041 ( .A(n6113), .B(n5979), .Z(n6112) );
  XNOR U6042 ( .A(p_input[225]), .B(n6114), .Z(n5979) );
  AND U6043 ( .A(n274), .B(n6115), .Z(n6114) );
  XNOR U6044 ( .A(p_input[241]), .B(n6116), .Z(n6115) );
  IV U6045 ( .A(p_input[225]), .Z(n6116) );
  XNOR U6046 ( .A(n5976), .B(n6109), .Z(n6111) );
  XNOR U6047 ( .A(p_input[193]), .B(n6117), .Z(n5976) );
  AND U6048 ( .A(n272), .B(n6118), .Z(n6117) );
  XOR U6049 ( .A(p_input[209]), .B(p_input[193]), .Z(n6118) );
  IV U6050 ( .A(n6113), .Z(n6109) );
  AND U6051 ( .A(n5984), .B(n5987), .Z(n6113) );
  XOR U6052 ( .A(p_input[224]), .B(n6119), .Z(n5987) );
  AND U6053 ( .A(n274), .B(n6120), .Z(n6119) );
  XOR U6054 ( .A(p_input[240]), .B(p_input[224]), .Z(n6120) );
  XOR U6055 ( .A(n6121), .B(n6122), .Z(n274) );
  AND U6056 ( .A(n6123), .B(n6124), .Z(n6122) );
  XNOR U6057 ( .A(p_input[255]), .B(n6121), .Z(n6124) );
  XOR U6058 ( .A(n6121), .B(p_input[239]), .Z(n6123) );
  XOR U6059 ( .A(n6125), .B(n6126), .Z(n6121) );
  AND U6060 ( .A(n6127), .B(n6128), .Z(n6126) );
  XNOR U6061 ( .A(p_input[254]), .B(n6125), .Z(n6128) );
  XOR U6062 ( .A(n6125), .B(p_input[238]), .Z(n6127) );
  XOR U6063 ( .A(n6129), .B(n6130), .Z(n6125) );
  AND U6064 ( .A(n6131), .B(n6132), .Z(n6130) );
  XNOR U6065 ( .A(p_input[253]), .B(n6129), .Z(n6132) );
  XOR U6066 ( .A(n6129), .B(p_input[237]), .Z(n6131) );
  XOR U6067 ( .A(n6133), .B(n6134), .Z(n6129) );
  AND U6068 ( .A(n6135), .B(n6136), .Z(n6134) );
  XNOR U6069 ( .A(p_input[252]), .B(n6133), .Z(n6136) );
  XOR U6070 ( .A(n6133), .B(p_input[236]), .Z(n6135) );
  XOR U6071 ( .A(n6137), .B(n6138), .Z(n6133) );
  AND U6072 ( .A(n6139), .B(n6140), .Z(n6138) );
  XNOR U6073 ( .A(p_input[251]), .B(n6137), .Z(n6140) );
  XOR U6074 ( .A(n6137), .B(p_input[235]), .Z(n6139) );
  XOR U6075 ( .A(n6141), .B(n6142), .Z(n6137) );
  AND U6076 ( .A(n6143), .B(n6144), .Z(n6142) );
  XNOR U6077 ( .A(p_input[250]), .B(n6141), .Z(n6144) );
  XOR U6078 ( .A(n6141), .B(p_input[234]), .Z(n6143) );
  XOR U6079 ( .A(n6145), .B(n6146), .Z(n6141) );
  AND U6080 ( .A(n6147), .B(n6148), .Z(n6146) );
  XNOR U6081 ( .A(p_input[249]), .B(n6145), .Z(n6148) );
  XOR U6082 ( .A(n6145), .B(p_input[233]), .Z(n6147) );
  XOR U6083 ( .A(n6149), .B(n6150), .Z(n6145) );
  AND U6084 ( .A(n6151), .B(n6152), .Z(n6150) );
  XNOR U6085 ( .A(p_input[248]), .B(n6149), .Z(n6152) );
  XOR U6086 ( .A(n6149), .B(p_input[232]), .Z(n6151) );
  XOR U6087 ( .A(n6153), .B(n6154), .Z(n6149) );
  AND U6088 ( .A(n6155), .B(n6156), .Z(n6154) );
  XNOR U6089 ( .A(p_input[247]), .B(n6153), .Z(n6156) );
  XOR U6090 ( .A(n6153), .B(p_input[231]), .Z(n6155) );
  XOR U6091 ( .A(n6157), .B(n6158), .Z(n6153) );
  AND U6092 ( .A(n6159), .B(n6160), .Z(n6158) );
  XNOR U6093 ( .A(p_input[246]), .B(n6157), .Z(n6160) );
  XOR U6094 ( .A(n6157), .B(p_input[230]), .Z(n6159) );
  XOR U6095 ( .A(n6161), .B(n6162), .Z(n6157) );
  AND U6096 ( .A(n6163), .B(n6164), .Z(n6162) );
  XNOR U6097 ( .A(p_input[245]), .B(n6161), .Z(n6164) );
  XOR U6098 ( .A(n6161), .B(p_input[229]), .Z(n6163) );
  XOR U6099 ( .A(n6165), .B(n6166), .Z(n6161) );
  AND U6100 ( .A(n6167), .B(n6168), .Z(n6166) );
  XNOR U6101 ( .A(p_input[244]), .B(n6165), .Z(n6168) );
  XOR U6102 ( .A(n6165), .B(p_input[228]), .Z(n6167) );
  XOR U6103 ( .A(n6169), .B(n6170), .Z(n6165) );
  AND U6104 ( .A(n6171), .B(n6172), .Z(n6170) );
  XNOR U6105 ( .A(p_input[243]), .B(n6169), .Z(n6172) );
  XOR U6106 ( .A(n6169), .B(p_input[227]), .Z(n6171) );
  XOR U6107 ( .A(n6173), .B(n6174), .Z(n6169) );
  AND U6108 ( .A(n6175), .B(n6176), .Z(n6174) );
  XNOR U6109 ( .A(p_input[242]), .B(n6173), .Z(n6176) );
  XOR U6110 ( .A(n6173), .B(p_input[226]), .Z(n6175) );
  XNOR U6111 ( .A(n6177), .B(n6178), .Z(n6173) );
  AND U6112 ( .A(n6179), .B(n6180), .Z(n6178) );
  XOR U6113 ( .A(p_input[241]), .B(n6177), .Z(n6180) );
  XNOR U6114 ( .A(p_input[225]), .B(n6177), .Z(n6179) );
  AND U6115 ( .A(p_input[240]), .B(n6181), .Z(n6177) );
  IV U6116 ( .A(p_input[224]), .Z(n6181) );
  XNOR U6117 ( .A(p_input[192]), .B(n6182), .Z(n5984) );
  AND U6118 ( .A(n272), .B(n6183), .Z(n6182) );
  XOR U6119 ( .A(p_input[208]), .B(p_input[192]), .Z(n6183) );
  XOR U6120 ( .A(n6184), .B(n6185), .Z(n272) );
  AND U6121 ( .A(n6186), .B(n6187), .Z(n6185) );
  XNOR U6122 ( .A(p_input[223]), .B(n6184), .Z(n6187) );
  XOR U6123 ( .A(n6184), .B(p_input[207]), .Z(n6186) );
  XOR U6124 ( .A(n6188), .B(n6189), .Z(n6184) );
  AND U6125 ( .A(n6190), .B(n6191), .Z(n6189) );
  XNOR U6126 ( .A(p_input[222]), .B(n6188), .Z(n6191) );
  XNOR U6127 ( .A(n6188), .B(n5998), .Z(n6190) );
  IV U6128 ( .A(p_input[206]), .Z(n5998) );
  XOR U6129 ( .A(n6192), .B(n6193), .Z(n6188) );
  AND U6130 ( .A(n6194), .B(n6195), .Z(n6193) );
  XNOR U6131 ( .A(p_input[221]), .B(n6192), .Z(n6195) );
  XNOR U6132 ( .A(n6192), .B(n6007), .Z(n6194) );
  IV U6133 ( .A(p_input[205]), .Z(n6007) );
  XOR U6134 ( .A(n6196), .B(n6197), .Z(n6192) );
  AND U6135 ( .A(n6198), .B(n6199), .Z(n6197) );
  XNOR U6136 ( .A(p_input[220]), .B(n6196), .Z(n6199) );
  XNOR U6137 ( .A(n6196), .B(n6016), .Z(n6198) );
  IV U6138 ( .A(p_input[204]), .Z(n6016) );
  XOR U6139 ( .A(n6200), .B(n6201), .Z(n6196) );
  AND U6140 ( .A(n6202), .B(n6203), .Z(n6201) );
  XNOR U6141 ( .A(p_input[219]), .B(n6200), .Z(n6203) );
  XNOR U6142 ( .A(n6200), .B(n6025), .Z(n6202) );
  IV U6143 ( .A(p_input[203]), .Z(n6025) );
  XOR U6144 ( .A(n6204), .B(n6205), .Z(n6200) );
  AND U6145 ( .A(n6206), .B(n6207), .Z(n6205) );
  XNOR U6146 ( .A(p_input[218]), .B(n6204), .Z(n6207) );
  XNOR U6147 ( .A(n6204), .B(n6034), .Z(n6206) );
  IV U6148 ( .A(p_input[202]), .Z(n6034) );
  XOR U6149 ( .A(n6208), .B(n6209), .Z(n6204) );
  AND U6150 ( .A(n6210), .B(n6211), .Z(n6209) );
  XNOR U6151 ( .A(p_input[217]), .B(n6208), .Z(n6211) );
  XNOR U6152 ( .A(n6208), .B(n6043), .Z(n6210) );
  IV U6153 ( .A(p_input[201]), .Z(n6043) );
  XOR U6154 ( .A(n6212), .B(n6213), .Z(n6208) );
  AND U6155 ( .A(n6214), .B(n6215), .Z(n6213) );
  XNOR U6156 ( .A(p_input[216]), .B(n6212), .Z(n6215) );
  XNOR U6157 ( .A(n6212), .B(n6052), .Z(n6214) );
  IV U6158 ( .A(p_input[200]), .Z(n6052) );
  XOR U6159 ( .A(n6216), .B(n6217), .Z(n6212) );
  AND U6160 ( .A(n6218), .B(n6219), .Z(n6217) );
  XNOR U6161 ( .A(p_input[215]), .B(n6216), .Z(n6219) );
  XNOR U6162 ( .A(n6216), .B(n6061), .Z(n6218) );
  IV U6163 ( .A(p_input[199]), .Z(n6061) );
  XOR U6164 ( .A(n6220), .B(n6221), .Z(n6216) );
  AND U6165 ( .A(n6222), .B(n6223), .Z(n6221) );
  XNOR U6166 ( .A(p_input[214]), .B(n6220), .Z(n6223) );
  XNOR U6167 ( .A(n6220), .B(n6070), .Z(n6222) );
  IV U6168 ( .A(p_input[198]), .Z(n6070) );
  XOR U6169 ( .A(n6224), .B(n6225), .Z(n6220) );
  AND U6170 ( .A(n6226), .B(n6227), .Z(n6225) );
  XNOR U6171 ( .A(p_input[213]), .B(n6224), .Z(n6227) );
  XNOR U6172 ( .A(n6224), .B(n6079), .Z(n6226) );
  IV U6173 ( .A(p_input[197]), .Z(n6079) );
  XOR U6174 ( .A(n6228), .B(n6229), .Z(n6224) );
  AND U6175 ( .A(n6230), .B(n6231), .Z(n6229) );
  XNOR U6176 ( .A(p_input[212]), .B(n6228), .Z(n6231) );
  XNOR U6177 ( .A(n6228), .B(n6088), .Z(n6230) );
  IV U6178 ( .A(p_input[196]), .Z(n6088) );
  XOR U6179 ( .A(n6232), .B(n6233), .Z(n6228) );
  AND U6180 ( .A(n6234), .B(n6235), .Z(n6233) );
  XNOR U6181 ( .A(p_input[211]), .B(n6232), .Z(n6235) );
  XNOR U6182 ( .A(n6232), .B(n6097), .Z(n6234) );
  IV U6183 ( .A(p_input[195]), .Z(n6097) );
  XOR U6184 ( .A(n6236), .B(n6237), .Z(n6232) );
  AND U6185 ( .A(n6238), .B(n6239), .Z(n6237) );
  XNOR U6186 ( .A(p_input[210]), .B(n6236), .Z(n6239) );
  XNOR U6187 ( .A(n6236), .B(n6106), .Z(n6238) );
  IV U6188 ( .A(p_input[194]), .Z(n6106) );
  XNOR U6189 ( .A(n6240), .B(n6241), .Z(n6236) );
  AND U6190 ( .A(n6242), .B(n6243), .Z(n6241) );
  XOR U6191 ( .A(p_input[209]), .B(n6240), .Z(n6243) );
  XNOR U6192 ( .A(p_input[193]), .B(n6240), .Z(n6242) );
  AND U6193 ( .A(p_input[208]), .B(n6244), .Z(n6240) );
  IV U6194 ( .A(p_input[192]), .Z(n6244) );
  XOR U6195 ( .A(n6245), .B(n6246), .Z(n5803) );
  AND U6196 ( .A(n196), .B(n6247), .Z(n6246) );
  XNOR U6197 ( .A(n6248), .B(n6245), .Z(n6247) );
  XOR U6198 ( .A(n6249), .B(n6250), .Z(n196) );
  AND U6199 ( .A(n6251), .B(n6252), .Z(n6250) );
  XNOR U6200 ( .A(n5813), .B(n6249), .Z(n6252) );
  AND U6201 ( .A(p_input[191]), .B(p_input[175]), .Z(n5813) );
  XOR U6202 ( .A(n6249), .B(n5814), .Z(n6251) );
  AND U6203 ( .A(p_input[159]), .B(p_input[143]), .Z(n5814) );
  XOR U6204 ( .A(n6253), .B(n6254), .Z(n6249) );
  AND U6205 ( .A(n6255), .B(n6256), .Z(n6254) );
  XOR U6206 ( .A(n6253), .B(n5826), .Z(n6256) );
  XNOR U6207 ( .A(p_input[174]), .B(n6257), .Z(n5826) );
  AND U6208 ( .A(n278), .B(n6258), .Z(n6257) );
  XOR U6209 ( .A(p_input[190]), .B(p_input[174]), .Z(n6258) );
  XNOR U6210 ( .A(n5823), .B(n6253), .Z(n6255) );
  XOR U6211 ( .A(n6259), .B(n6260), .Z(n5823) );
  AND U6212 ( .A(n275), .B(n6261), .Z(n6260) );
  XOR U6213 ( .A(p_input[158]), .B(p_input[142]), .Z(n6261) );
  XOR U6214 ( .A(n6262), .B(n6263), .Z(n6253) );
  AND U6215 ( .A(n6264), .B(n6265), .Z(n6263) );
  XOR U6216 ( .A(n6262), .B(n5838), .Z(n6265) );
  XNOR U6217 ( .A(p_input[173]), .B(n6266), .Z(n5838) );
  AND U6218 ( .A(n278), .B(n6267), .Z(n6266) );
  XOR U6219 ( .A(p_input[189]), .B(p_input[173]), .Z(n6267) );
  XNOR U6220 ( .A(n5835), .B(n6262), .Z(n6264) );
  XOR U6221 ( .A(n6268), .B(n6269), .Z(n5835) );
  AND U6222 ( .A(n275), .B(n6270), .Z(n6269) );
  XOR U6223 ( .A(p_input[157]), .B(p_input[141]), .Z(n6270) );
  XOR U6224 ( .A(n6271), .B(n6272), .Z(n6262) );
  AND U6225 ( .A(n6273), .B(n6274), .Z(n6272) );
  XOR U6226 ( .A(n6271), .B(n5850), .Z(n6274) );
  XNOR U6227 ( .A(p_input[172]), .B(n6275), .Z(n5850) );
  AND U6228 ( .A(n278), .B(n6276), .Z(n6275) );
  XOR U6229 ( .A(p_input[188]), .B(p_input[172]), .Z(n6276) );
  XNOR U6230 ( .A(n5847), .B(n6271), .Z(n6273) );
  XOR U6231 ( .A(n6277), .B(n6278), .Z(n5847) );
  AND U6232 ( .A(n275), .B(n6279), .Z(n6278) );
  XOR U6233 ( .A(p_input[156]), .B(p_input[140]), .Z(n6279) );
  XOR U6234 ( .A(n6280), .B(n6281), .Z(n6271) );
  AND U6235 ( .A(n6282), .B(n6283), .Z(n6281) );
  XOR U6236 ( .A(n6280), .B(n5862), .Z(n6283) );
  XNOR U6237 ( .A(p_input[171]), .B(n6284), .Z(n5862) );
  AND U6238 ( .A(n278), .B(n6285), .Z(n6284) );
  XOR U6239 ( .A(p_input[187]), .B(p_input[171]), .Z(n6285) );
  XNOR U6240 ( .A(n5859), .B(n6280), .Z(n6282) );
  XOR U6241 ( .A(n6286), .B(n6287), .Z(n5859) );
  AND U6242 ( .A(n275), .B(n6288), .Z(n6287) );
  XOR U6243 ( .A(p_input[155]), .B(p_input[139]), .Z(n6288) );
  XOR U6244 ( .A(n6289), .B(n6290), .Z(n6280) );
  AND U6245 ( .A(n6291), .B(n6292), .Z(n6290) );
  XOR U6246 ( .A(n6289), .B(n5874), .Z(n6292) );
  XNOR U6247 ( .A(p_input[170]), .B(n6293), .Z(n5874) );
  AND U6248 ( .A(n278), .B(n6294), .Z(n6293) );
  XOR U6249 ( .A(p_input[186]), .B(p_input[170]), .Z(n6294) );
  XNOR U6250 ( .A(n5871), .B(n6289), .Z(n6291) );
  XOR U6251 ( .A(n6295), .B(n6296), .Z(n5871) );
  AND U6252 ( .A(n275), .B(n6297), .Z(n6296) );
  XOR U6253 ( .A(p_input[154]), .B(p_input[138]), .Z(n6297) );
  XOR U6254 ( .A(n6298), .B(n6299), .Z(n6289) );
  AND U6255 ( .A(n6300), .B(n6301), .Z(n6299) );
  XOR U6256 ( .A(n6298), .B(n5886), .Z(n6301) );
  XNOR U6257 ( .A(p_input[169]), .B(n6302), .Z(n5886) );
  AND U6258 ( .A(n278), .B(n6303), .Z(n6302) );
  XOR U6259 ( .A(p_input[185]), .B(p_input[169]), .Z(n6303) );
  XNOR U6260 ( .A(n5883), .B(n6298), .Z(n6300) );
  XOR U6261 ( .A(n6304), .B(n6305), .Z(n5883) );
  AND U6262 ( .A(n275), .B(n6306), .Z(n6305) );
  XOR U6263 ( .A(p_input[153]), .B(p_input[137]), .Z(n6306) );
  XOR U6264 ( .A(n6307), .B(n6308), .Z(n6298) );
  AND U6265 ( .A(n6309), .B(n6310), .Z(n6308) );
  XOR U6266 ( .A(n6307), .B(n5898), .Z(n6310) );
  XNOR U6267 ( .A(p_input[168]), .B(n6311), .Z(n5898) );
  AND U6268 ( .A(n278), .B(n6312), .Z(n6311) );
  XOR U6269 ( .A(p_input[184]), .B(p_input[168]), .Z(n6312) );
  XNOR U6270 ( .A(n5895), .B(n6307), .Z(n6309) );
  XOR U6271 ( .A(n6313), .B(n6314), .Z(n5895) );
  AND U6272 ( .A(n275), .B(n6315), .Z(n6314) );
  XOR U6273 ( .A(p_input[152]), .B(p_input[136]), .Z(n6315) );
  XOR U6274 ( .A(n6316), .B(n6317), .Z(n6307) );
  AND U6275 ( .A(n6318), .B(n6319), .Z(n6317) );
  XOR U6276 ( .A(n6316), .B(n5910), .Z(n6319) );
  XNOR U6277 ( .A(p_input[167]), .B(n6320), .Z(n5910) );
  AND U6278 ( .A(n278), .B(n6321), .Z(n6320) );
  XOR U6279 ( .A(p_input[183]), .B(p_input[167]), .Z(n6321) );
  XNOR U6280 ( .A(n5907), .B(n6316), .Z(n6318) );
  XOR U6281 ( .A(n6322), .B(n6323), .Z(n5907) );
  AND U6282 ( .A(n275), .B(n6324), .Z(n6323) );
  XOR U6283 ( .A(p_input[151]), .B(p_input[135]), .Z(n6324) );
  XOR U6284 ( .A(n6325), .B(n6326), .Z(n6316) );
  AND U6285 ( .A(n6327), .B(n6328), .Z(n6326) );
  XOR U6286 ( .A(n6325), .B(n5922), .Z(n6328) );
  XNOR U6287 ( .A(p_input[166]), .B(n6329), .Z(n5922) );
  AND U6288 ( .A(n278), .B(n6330), .Z(n6329) );
  XOR U6289 ( .A(p_input[182]), .B(p_input[166]), .Z(n6330) );
  XNOR U6290 ( .A(n5919), .B(n6325), .Z(n6327) );
  XOR U6291 ( .A(n6331), .B(n6332), .Z(n5919) );
  AND U6292 ( .A(n275), .B(n6333), .Z(n6332) );
  XOR U6293 ( .A(p_input[150]), .B(p_input[134]), .Z(n6333) );
  XOR U6294 ( .A(n6334), .B(n6335), .Z(n6325) );
  AND U6295 ( .A(n6336), .B(n6337), .Z(n6335) );
  XOR U6296 ( .A(n6334), .B(n5934), .Z(n6337) );
  XNOR U6297 ( .A(p_input[165]), .B(n6338), .Z(n5934) );
  AND U6298 ( .A(n278), .B(n6339), .Z(n6338) );
  XOR U6299 ( .A(p_input[181]), .B(p_input[165]), .Z(n6339) );
  XNOR U6300 ( .A(n5931), .B(n6334), .Z(n6336) );
  XOR U6301 ( .A(n6340), .B(n6341), .Z(n5931) );
  AND U6302 ( .A(n275), .B(n6342), .Z(n6341) );
  XOR U6303 ( .A(p_input[149]), .B(p_input[133]), .Z(n6342) );
  XOR U6304 ( .A(n6343), .B(n6344), .Z(n6334) );
  AND U6305 ( .A(n6345), .B(n6346), .Z(n6344) );
  XOR U6306 ( .A(n6343), .B(n5946), .Z(n6346) );
  XNOR U6307 ( .A(p_input[164]), .B(n6347), .Z(n5946) );
  AND U6308 ( .A(n278), .B(n6348), .Z(n6347) );
  XOR U6309 ( .A(p_input[180]), .B(p_input[164]), .Z(n6348) );
  XNOR U6310 ( .A(n5943), .B(n6343), .Z(n6345) );
  XOR U6311 ( .A(n6349), .B(n6350), .Z(n5943) );
  AND U6312 ( .A(n275), .B(n6351), .Z(n6350) );
  XOR U6313 ( .A(p_input[148]), .B(p_input[132]), .Z(n6351) );
  XOR U6314 ( .A(n6352), .B(n6353), .Z(n6343) );
  AND U6315 ( .A(n6354), .B(n6355), .Z(n6353) );
  XOR U6316 ( .A(n5958), .B(n6352), .Z(n6355) );
  XNOR U6317 ( .A(p_input[163]), .B(n6356), .Z(n5958) );
  AND U6318 ( .A(n278), .B(n6357), .Z(n6356) );
  XOR U6319 ( .A(p_input[179]), .B(p_input[163]), .Z(n6357) );
  XNOR U6320 ( .A(n6352), .B(n5955), .Z(n6354) );
  XOR U6321 ( .A(n6358), .B(n6359), .Z(n5955) );
  AND U6322 ( .A(n275), .B(n6360), .Z(n6359) );
  XOR U6323 ( .A(p_input[147]), .B(p_input[131]), .Z(n6360) );
  XOR U6324 ( .A(n6361), .B(n6362), .Z(n6352) );
  AND U6325 ( .A(n6363), .B(n6364), .Z(n6362) );
  XOR U6326 ( .A(n6361), .B(n5970), .Z(n6364) );
  XNOR U6327 ( .A(p_input[162]), .B(n6365), .Z(n5970) );
  AND U6328 ( .A(n278), .B(n6366), .Z(n6365) );
  XOR U6329 ( .A(p_input[178]), .B(p_input[162]), .Z(n6366) );
  XNOR U6330 ( .A(n5967), .B(n6361), .Z(n6363) );
  XOR U6331 ( .A(n6367), .B(n6368), .Z(n5967) );
  AND U6332 ( .A(n275), .B(n6369), .Z(n6368) );
  XOR U6333 ( .A(p_input[146]), .B(p_input[130]), .Z(n6369) );
  XOR U6334 ( .A(n6370), .B(n6371), .Z(n6361) );
  AND U6335 ( .A(n6372), .B(n6373), .Z(n6371) );
  XNOR U6336 ( .A(n6374), .B(n5983), .Z(n6373) );
  XNOR U6337 ( .A(p_input[161]), .B(n6375), .Z(n5983) );
  AND U6338 ( .A(n278), .B(n6376), .Z(n6375) );
  XNOR U6339 ( .A(p_input[177]), .B(n6377), .Z(n6376) );
  IV U6340 ( .A(p_input[161]), .Z(n6377) );
  XNOR U6341 ( .A(n5980), .B(n6370), .Z(n6372) );
  XNOR U6342 ( .A(p_input[129]), .B(n6378), .Z(n5980) );
  AND U6343 ( .A(n275), .B(n6379), .Z(n6378) );
  XOR U6344 ( .A(p_input[145]), .B(p_input[129]), .Z(n6379) );
  IV U6345 ( .A(n6374), .Z(n6370) );
  AND U6346 ( .A(n6245), .B(n6248), .Z(n6374) );
  XOR U6347 ( .A(p_input[160]), .B(n6380), .Z(n6248) );
  AND U6348 ( .A(n278), .B(n6381), .Z(n6380) );
  XOR U6349 ( .A(p_input[176]), .B(p_input[160]), .Z(n6381) );
  XOR U6350 ( .A(n6382), .B(n6383), .Z(n278) );
  AND U6351 ( .A(n6384), .B(n6385), .Z(n6383) );
  XNOR U6352 ( .A(p_input[191]), .B(n6382), .Z(n6385) );
  XOR U6353 ( .A(n6382), .B(p_input[175]), .Z(n6384) );
  XOR U6354 ( .A(n6386), .B(n6387), .Z(n6382) );
  AND U6355 ( .A(n6388), .B(n6389), .Z(n6387) );
  XNOR U6356 ( .A(p_input[190]), .B(n6386), .Z(n6389) );
  XOR U6357 ( .A(n6386), .B(p_input[174]), .Z(n6388) );
  XOR U6358 ( .A(n6390), .B(n6391), .Z(n6386) );
  AND U6359 ( .A(n6392), .B(n6393), .Z(n6391) );
  XNOR U6360 ( .A(p_input[189]), .B(n6390), .Z(n6393) );
  XOR U6361 ( .A(n6390), .B(p_input[173]), .Z(n6392) );
  XOR U6362 ( .A(n6394), .B(n6395), .Z(n6390) );
  AND U6363 ( .A(n6396), .B(n6397), .Z(n6395) );
  XNOR U6364 ( .A(p_input[188]), .B(n6394), .Z(n6397) );
  XOR U6365 ( .A(n6394), .B(p_input[172]), .Z(n6396) );
  XOR U6366 ( .A(n6398), .B(n6399), .Z(n6394) );
  AND U6367 ( .A(n6400), .B(n6401), .Z(n6399) );
  XNOR U6368 ( .A(p_input[187]), .B(n6398), .Z(n6401) );
  XOR U6369 ( .A(n6398), .B(p_input[171]), .Z(n6400) );
  XOR U6370 ( .A(n6402), .B(n6403), .Z(n6398) );
  AND U6371 ( .A(n6404), .B(n6405), .Z(n6403) );
  XNOR U6372 ( .A(p_input[186]), .B(n6402), .Z(n6405) );
  XOR U6373 ( .A(n6402), .B(p_input[170]), .Z(n6404) );
  XOR U6374 ( .A(n6406), .B(n6407), .Z(n6402) );
  AND U6375 ( .A(n6408), .B(n6409), .Z(n6407) );
  XNOR U6376 ( .A(p_input[185]), .B(n6406), .Z(n6409) );
  XOR U6377 ( .A(n6406), .B(p_input[169]), .Z(n6408) );
  XOR U6378 ( .A(n6410), .B(n6411), .Z(n6406) );
  AND U6379 ( .A(n6412), .B(n6413), .Z(n6411) );
  XNOR U6380 ( .A(p_input[184]), .B(n6410), .Z(n6413) );
  XOR U6381 ( .A(n6410), .B(p_input[168]), .Z(n6412) );
  XOR U6382 ( .A(n6414), .B(n6415), .Z(n6410) );
  AND U6383 ( .A(n6416), .B(n6417), .Z(n6415) );
  XNOR U6384 ( .A(p_input[183]), .B(n6414), .Z(n6417) );
  XOR U6385 ( .A(n6414), .B(p_input[167]), .Z(n6416) );
  XOR U6386 ( .A(n6418), .B(n6419), .Z(n6414) );
  AND U6387 ( .A(n6420), .B(n6421), .Z(n6419) );
  XNOR U6388 ( .A(p_input[182]), .B(n6418), .Z(n6421) );
  XOR U6389 ( .A(n6418), .B(p_input[166]), .Z(n6420) );
  XOR U6390 ( .A(n6422), .B(n6423), .Z(n6418) );
  AND U6391 ( .A(n6424), .B(n6425), .Z(n6423) );
  XNOR U6392 ( .A(p_input[181]), .B(n6422), .Z(n6425) );
  XOR U6393 ( .A(n6422), .B(p_input[165]), .Z(n6424) );
  XOR U6394 ( .A(n6426), .B(n6427), .Z(n6422) );
  AND U6395 ( .A(n6428), .B(n6429), .Z(n6427) );
  XNOR U6396 ( .A(p_input[180]), .B(n6426), .Z(n6429) );
  XOR U6397 ( .A(n6426), .B(p_input[164]), .Z(n6428) );
  XOR U6398 ( .A(n6430), .B(n6431), .Z(n6426) );
  AND U6399 ( .A(n6432), .B(n6433), .Z(n6431) );
  XNOR U6400 ( .A(p_input[179]), .B(n6430), .Z(n6433) );
  XOR U6401 ( .A(n6430), .B(p_input[163]), .Z(n6432) );
  XOR U6402 ( .A(n6434), .B(n6435), .Z(n6430) );
  AND U6403 ( .A(n6436), .B(n6437), .Z(n6435) );
  XNOR U6404 ( .A(p_input[178]), .B(n6434), .Z(n6437) );
  XOR U6405 ( .A(n6434), .B(p_input[162]), .Z(n6436) );
  XNOR U6406 ( .A(n6438), .B(n6439), .Z(n6434) );
  AND U6407 ( .A(n6440), .B(n6441), .Z(n6439) );
  XOR U6408 ( .A(p_input[177]), .B(n6438), .Z(n6441) );
  XNOR U6409 ( .A(p_input[161]), .B(n6438), .Z(n6440) );
  AND U6410 ( .A(p_input[176]), .B(n6442), .Z(n6438) );
  IV U6411 ( .A(p_input[160]), .Z(n6442) );
  XNOR U6412 ( .A(p_input[128]), .B(n6443), .Z(n6245) );
  AND U6413 ( .A(n275), .B(n6444), .Z(n6443) );
  XOR U6414 ( .A(p_input[144]), .B(p_input[128]), .Z(n6444) );
  XOR U6415 ( .A(n6445), .B(n6446), .Z(n275) );
  AND U6416 ( .A(n6447), .B(n6448), .Z(n6446) );
  XNOR U6417 ( .A(p_input[159]), .B(n6445), .Z(n6448) );
  XOR U6418 ( .A(n6445), .B(p_input[143]), .Z(n6447) );
  XOR U6419 ( .A(n6449), .B(n6450), .Z(n6445) );
  AND U6420 ( .A(n6451), .B(n6452), .Z(n6450) );
  XNOR U6421 ( .A(p_input[158]), .B(n6449), .Z(n6452) );
  XNOR U6422 ( .A(n6449), .B(n6259), .Z(n6451) );
  IV U6423 ( .A(p_input[142]), .Z(n6259) );
  XOR U6424 ( .A(n6453), .B(n6454), .Z(n6449) );
  AND U6425 ( .A(n6455), .B(n6456), .Z(n6454) );
  XNOR U6426 ( .A(p_input[157]), .B(n6453), .Z(n6456) );
  XNOR U6427 ( .A(n6453), .B(n6268), .Z(n6455) );
  IV U6428 ( .A(p_input[141]), .Z(n6268) );
  XOR U6429 ( .A(n6457), .B(n6458), .Z(n6453) );
  AND U6430 ( .A(n6459), .B(n6460), .Z(n6458) );
  XNOR U6431 ( .A(p_input[156]), .B(n6457), .Z(n6460) );
  XNOR U6432 ( .A(n6457), .B(n6277), .Z(n6459) );
  IV U6433 ( .A(p_input[140]), .Z(n6277) );
  XOR U6434 ( .A(n6461), .B(n6462), .Z(n6457) );
  AND U6435 ( .A(n6463), .B(n6464), .Z(n6462) );
  XNOR U6436 ( .A(p_input[155]), .B(n6461), .Z(n6464) );
  XNOR U6437 ( .A(n6461), .B(n6286), .Z(n6463) );
  IV U6438 ( .A(p_input[139]), .Z(n6286) );
  XOR U6439 ( .A(n6465), .B(n6466), .Z(n6461) );
  AND U6440 ( .A(n6467), .B(n6468), .Z(n6466) );
  XNOR U6441 ( .A(p_input[154]), .B(n6465), .Z(n6468) );
  XNOR U6442 ( .A(n6465), .B(n6295), .Z(n6467) );
  IV U6443 ( .A(p_input[138]), .Z(n6295) );
  XOR U6444 ( .A(n6469), .B(n6470), .Z(n6465) );
  AND U6445 ( .A(n6471), .B(n6472), .Z(n6470) );
  XNOR U6446 ( .A(p_input[153]), .B(n6469), .Z(n6472) );
  XNOR U6447 ( .A(n6469), .B(n6304), .Z(n6471) );
  IV U6448 ( .A(p_input[137]), .Z(n6304) );
  XOR U6449 ( .A(n6473), .B(n6474), .Z(n6469) );
  AND U6450 ( .A(n6475), .B(n6476), .Z(n6474) );
  XNOR U6451 ( .A(p_input[152]), .B(n6473), .Z(n6476) );
  XNOR U6452 ( .A(n6473), .B(n6313), .Z(n6475) );
  IV U6453 ( .A(p_input[136]), .Z(n6313) );
  XOR U6454 ( .A(n6477), .B(n6478), .Z(n6473) );
  AND U6455 ( .A(n6479), .B(n6480), .Z(n6478) );
  XNOR U6456 ( .A(p_input[151]), .B(n6477), .Z(n6480) );
  XNOR U6457 ( .A(n6477), .B(n6322), .Z(n6479) );
  IV U6458 ( .A(p_input[135]), .Z(n6322) );
  XOR U6459 ( .A(n6481), .B(n6482), .Z(n6477) );
  AND U6460 ( .A(n6483), .B(n6484), .Z(n6482) );
  XNOR U6461 ( .A(p_input[150]), .B(n6481), .Z(n6484) );
  XNOR U6462 ( .A(n6481), .B(n6331), .Z(n6483) );
  IV U6463 ( .A(p_input[134]), .Z(n6331) );
  XOR U6464 ( .A(n6485), .B(n6486), .Z(n6481) );
  AND U6465 ( .A(n6487), .B(n6488), .Z(n6486) );
  XNOR U6466 ( .A(p_input[149]), .B(n6485), .Z(n6488) );
  XNOR U6467 ( .A(n6485), .B(n6340), .Z(n6487) );
  IV U6468 ( .A(p_input[133]), .Z(n6340) );
  XOR U6469 ( .A(n6489), .B(n6490), .Z(n6485) );
  AND U6470 ( .A(n6491), .B(n6492), .Z(n6490) );
  XNOR U6471 ( .A(p_input[148]), .B(n6489), .Z(n6492) );
  XNOR U6472 ( .A(n6489), .B(n6349), .Z(n6491) );
  IV U6473 ( .A(p_input[132]), .Z(n6349) );
  XOR U6474 ( .A(n6493), .B(n6494), .Z(n6489) );
  AND U6475 ( .A(n6495), .B(n6496), .Z(n6494) );
  XNOR U6476 ( .A(p_input[147]), .B(n6493), .Z(n6496) );
  XNOR U6477 ( .A(n6493), .B(n6358), .Z(n6495) );
  IV U6478 ( .A(p_input[131]), .Z(n6358) );
  XOR U6479 ( .A(n6497), .B(n6498), .Z(n6493) );
  AND U6480 ( .A(n6499), .B(n6500), .Z(n6498) );
  XNOR U6481 ( .A(p_input[146]), .B(n6497), .Z(n6500) );
  XNOR U6482 ( .A(n6497), .B(n6367), .Z(n6499) );
  IV U6483 ( .A(p_input[130]), .Z(n6367) );
  XNOR U6484 ( .A(n6501), .B(n6502), .Z(n6497) );
  AND U6485 ( .A(n6503), .B(n6504), .Z(n6502) );
  XOR U6486 ( .A(p_input[145]), .B(n6501), .Z(n6504) );
  XNOR U6487 ( .A(p_input[129]), .B(n6501), .Z(n6503) );
  AND U6488 ( .A(p_input[144]), .B(n6505), .Z(n6501) );
  IV U6489 ( .A(p_input[128]), .Z(n6505) );
  XOR U6490 ( .A(n6506), .B(n6507), .Z(n5621) );
  AND U6491 ( .A(n259), .B(n6508), .Z(n6507) );
  XNOR U6492 ( .A(n6509), .B(n6506), .Z(n6508) );
  XOR U6493 ( .A(n6510), .B(n6511), .Z(n259) );
  AND U6494 ( .A(n6512), .B(n6513), .Z(n6511) );
  XNOR U6495 ( .A(n5633), .B(n6510), .Z(n6513) );
  AND U6496 ( .A(n6514), .B(n6515), .Z(n5633) );
  XOR U6497 ( .A(n6510), .B(n5632), .Z(n6512) );
  AND U6498 ( .A(n6516), .B(n6517), .Z(n5632) );
  XOR U6499 ( .A(n6518), .B(n6519), .Z(n6510) );
  AND U6500 ( .A(n6520), .B(n6521), .Z(n6519) );
  XOR U6501 ( .A(n6518), .B(n5645), .Z(n6521) );
  XOR U6502 ( .A(n6522), .B(n6523), .Z(n5645) );
  AND U6503 ( .A(n202), .B(n6524), .Z(n6523) );
  XOR U6504 ( .A(n6525), .B(n6522), .Z(n6524) );
  XNOR U6505 ( .A(n5642), .B(n6518), .Z(n6520) );
  XOR U6506 ( .A(n6526), .B(n6527), .Z(n5642) );
  AND U6507 ( .A(n199), .B(n6528), .Z(n6527) );
  XOR U6508 ( .A(n6529), .B(n6526), .Z(n6528) );
  XOR U6509 ( .A(n6530), .B(n6531), .Z(n6518) );
  AND U6510 ( .A(n6532), .B(n6533), .Z(n6531) );
  XOR U6511 ( .A(n6530), .B(n5657), .Z(n6533) );
  XOR U6512 ( .A(n6534), .B(n6535), .Z(n5657) );
  AND U6513 ( .A(n202), .B(n6536), .Z(n6535) );
  XOR U6514 ( .A(n6537), .B(n6534), .Z(n6536) );
  XNOR U6515 ( .A(n5654), .B(n6530), .Z(n6532) );
  XOR U6516 ( .A(n6538), .B(n6539), .Z(n5654) );
  AND U6517 ( .A(n199), .B(n6540), .Z(n6539) );
  XOR U6518 ( .A(n6541), .B(n6538), .Z(n6540) );
  XOR U6519 ( .A(n6542), .B(n6543), .Z(n6530) );
  AND U6520 ( .A(n6544), .B(n6545), .Z(n6543) );
  XOR U6521 ( .A(n6542), .B(n5669), .Z(n6545) );
  XOR U6522 ( .A(n6546), .B(n6547), .Z(n5669) );
  AND U6523 ( .A(n202), .B(n6548), .Z(n6547) );
  XOR U6524 ( .A(n6549), .B(n6546), .Z(n6548) );
  XNOR U6525 ( .A(n5666), .B(n6542), .Z(n6544) );
  XOR U6526 ( .A(n6550), .B(n6551), .Z(n5666) );
  AND U6527 ( .A(n199), .B(n6552), .Z(n6551) );
  XOR U6528 ( .A(n6553), .B(n6550), .Z(n6552) );
  XOR U6529 ( .A(n6554), .B(n6555), .Z(n6542) );
  AND U6530 ( .A(n6556), .B(n6557), .Z(n6555) );
  XOR U6531 ( .A(n6554), .B(n5681), .Z(n6557) );
  XOR U6532 ( .A(n6558), .B(n6559), .Z(n5681) );
  AND U6533 ( .A(n202), .B(n6560), .Z(n6559) );
  XOR U6534 ( .A(n6561), .B(n6558), .Z(n6560) );
  XNOR U6535 ( .A(n5678), .B(n6554), .Z(n6556) );
  XOR U6536 ( .A(n6562), .B(n6563), .Z(n5678) );
  AND U6537 ( .A(n199), .B(n6564), .Z(n6563) );
  XOR U6538 ( .A(n6565), .B(n6562), .Z(n6564) );
  XOR U6539 ( .A(n6566), .B(n6567), .Z(n6554) );
  AND U6540 ( .A(n6568), .B(n6569), .Z(n6567) );
  XOR U6541 ( .A(n6566), .B(n5693), .Z(n6569) );
  XOR U6542 ( .A(n6570), .B(n6571), .Z(n5693) );
  AND U6543 ( .A(n202), .B(n6572), .Z(n6571) );
  XOR U6544 ( .A(n6573), .B(n6570), .Z(n6572) );
  XNOR U6545 ( .A(n5690), .B(n6566), .Z(n6568) );
  XOR U6546 ( .A(n6574), .B(n6575), .Z(n5690) );
  AND U6547 ( .A(n199), .B(n6576), .Z(n6575) );
  XOR U6548 ( .A(n6577), .B(n6574), .Z(n6576) );
  XOR U6549 ( .A(n6578), .B(n6579), .Z(n6566) );
  AND U6550 ( .A(n6580), .B(n6581), .Z(n6579) );
  XOR U6551 ( .A(n6578), .B(n5705), .Z(n6581) );
  XOR U6552 ( .A(n6582), .B(n6583), .Z(n5705) );
  AND U6553 ( .A(n202), .B(n6584), .Z(n6583) );
  XOR U6554 ( .A(n6585), .B(n6582), .Z(n6584) );
  XNOR U6555 ( .A(n5702), .B(n6578), .Z(n6580) );
  XOR U6556 ( .A(n6586), .B(n6587), .Z(n5702) );
  AND U6557 ( .A(n199), .B(n6588), .Z(n6587) );
  XOR U6558 ( .A(n6589), .B(n6586), .Z(n6588) );
  XOR U6559 ( .A(n6590), .B(n6591), .Z(n6578) );
  AND U6560 ( .A(n6592), .B(n6593), .Z(n6591) );
  XOR U6561 ( .A(n6590), .B(n5717), .Z(n6593) );
  XOR U6562 ( .A(n6594), .B(n6595), .Z(n5717) );
  AND U6563 ( .A(n202), .B(n6596), .Z(n6595) );
  XOR U6564 ( .A(n6597), .B(n6594), .Z(n6596) );
  XNOR U6565 ( .A(n5714), .B(n6590), .Z(n6592) );
  XOR U6566 ( .A(n6598), .B(n6599), .Z(n5714) );
  AND U6567 ( .A(n199), .B(n6600), .Z(n6599) );
  XOR U6568 ( .A(n6601), .B(n6598), .Z(n6600) );
  XOR U6569 ( .A(n6602), .B(n6603), .Z(n6590) );
  AND U6570 ( .A(n6604), .B(n6605), .Z(n6603) );
  XOR U6571 ( .A(n6602), .B(n5729), .Z(n6605) );
  XOR U6572 ( .A(n6606), .B(n6607), .Z(n5729) );
  AND U6573 ( .A(n202), .B(n6608), .Z(n6607) );
  XOR U6574 ( .A(n6609), .B(n6606), .Z(n6608) );
  XNOR U6575 ( .A(n5726), .B(n6602), .Z(n6604) );
  XOR U6576 ( .A(n6610), .B(n6611), .Z(n5726) );
  AND U6577 ( .A(n199), .B(n6612), .Z(n6611) );
  XOR U6578 ( .A(n6613), .B(n6610), .Z(n6612) );
  XOR U6579 ( .A(n6614), .B(n6615), .Z(n6602) );
  AND U6580 ( .A(n6616), .B(n6617), .Z(n6615) );
  XOR U6581 ( .A(n6614), .B(n5741), .Z(n6617) );
  XOR U6582 ( .A(n6618), .B(n6619), .Z(n5741) );
  AND U6583 ( .A(n202), .B(n6620), .Z(n6619) );
  XOR U6584 ( .A(n6621), .B(n6618), .Z(n6620) );
  XNOR U6585 ( .A(n5738), .B(n6614), .Z(n6616) );
  XOR U6586 ( .A(n6622), .B(n6623), .Z(n5738) );
  AND U6587 ( .A(n199), .B(n6624), .Z(n6623) );
  XOR U6588 ( .A(n6625), .B(n6622), .Z(n6624) );
  XOR U6589 ( .A(n6626), .B(n6627), .Z(n6614) );
  AND U6590 ( .A(n6628), .B(n6629), .Z(n6627) );
  XOR U6591 ( .A(n6626), .B(n5753), .Z(n6629) );
  XOR U6592 ( .A(n6630), .B(n6631), .Z(n5753) );
  AND U6593 ( .A(n202), .B(n6632), .Z(n6631) );
  XOR U6594 ( .A(n6633), .B(n6630), .Z(n6632) );
  XNOR U6595 ( .A(n5750), .B(n6626), .Z(n6628) );
  XOR U6596 ( .A(n6634), .B(n6635), .Z(n5750) );
  AND U6597 ( .A(n199), .B(n6636), .Z(n6635) );
  XOR U6598 ( .A(n6637), .B(n6634), .Z(n6636) );
  XOR U6599 ( .A(n6638), .B(n6639), .Z(n6626) );
  AND U6600 ( .A(n6640), .B(n6641), .Z(n6639) );
  XOR U6601 ( .A(n6638), .B(n5765), .Z(n6641) );
  XOR U6602 ( .A(n6642), .B(n6643), .Z(n5765) );
  AND U6603 ( .A(n202), .B(n6644), .Z(n6643) );
  XOR U6604 ( .A(n6645), .B(n6642), .Z(n6644) );
  XNOR U6605 ( .A(n5762), .B(n6638), .Z(n6640) );
  XOR U6606 ( .A(n6646), .B(n6647), .Z(n5762) );
  AND U6607 ( .A(n199), .B(n6648), .Z(n6647) );
  XOR U6608 ( .A(n6649), .B(n6646), .Z(n6648) );
  XOR U6609 ( .A(n6650), .B(n6651), .Z(n6638) );
  AND U6610 ( .A(n6652), .B(n6653), .Z(n6651) );
  XOR U6611 ( .A(n5777), .B(n6650), .Z(n6653) );
  XOR U6612 ( .A(n6654), .B(n6655), .Z(n5777) );
  AND U6613 ( .A(n202), .B(n6656), .Z(n6655) );
  XOR U6614 ( .A(n6654), .B(n6657), .Z(n6656) );
  XNOR U6615 ( .A(n6650), .B(n5774), .Z(n6652) );
  XOR U6616 ( .A(n6658), .B(n6659), .Z(n5774) );
  AND U6617 ( .A(n199), .B(n6660), .Z(n6659) );
  XOR U6618 ( .A(n6658), .B(n6661), .Z(n6660) );
  XOR U6619 ( .A(n6662), .B(n6663), .Z(n6650) );
  AND U6620 ( .A(n6664), .B(n6665), .Z(n6663) );
  XOR U6621 ( .A(n6662), .B(n5789), .Z(n6665) );
  XOR U6622 ( .A(n6666), .B(n6667), .Z(n5789) );
  AND U6623 ( .A(n202), .B(n6668), .Z(n6667) );
  XOR U6624 ( .A(n6669), .B(n6666), .Z(n6668) );
  XNOR U6625 ( .A(n5786), .B(n6662), .Z(n6664) );
  XOR U6626 ( .A(n6670), .B(n6671), .Z(n5786) );
  AND U6627 ( .A(n199), .B(n6672), .Z(n6671) );
  XOR U6628 ( .A(n6673), .B(n6670), .Z(n6672) );
  XOR U6629 ( .A(n6674), .B(n6675), .Z(n6662) );
  AND U6630 ( .A(n6676), .B(n6677), .Z(n6675) );
  XNOR U6631 ( .A(n6678), .B(n5802), .Z(n6677) );
  XOR U6632 ( .A(n6679), .B(n6680), .Z(n5802) );
  AND U6633 ( .A(n202), .B(n6681), .Z(n6680) );
  XOR U6634 ( .A(n6682), .B(n6679), .Z(n6681) );
  XNOR U6635 ( .A(n5799), .B(n6674), .Z(n6676) );
  XOR U6636 ( .A(n6683), .B(n6684), .Z(n5799) );
  AND U6637 ( .A(n199), .B(n6685), .Z(n6684) );
  XOR U6638 ( .A(n6686), .B(n6683), .Z(n6685) );
  IV U6639 ( .A(n6678), .Z(n6674) );
  AND U6640 ( .A(n6506), .B(n6509), .Z(n6678) );
  XNOR U6641 ( .A(n6687), .B(n6688), .Z(n6509) );
  AND U6642 ( .A(n202), .B(n6689), .Z(n6688) );
  XNOR U6643 ( .A(n6690), .B(n6687), .Z(n6689) );
  XOR U6644 ( .A(n6691), .B(n6692), .Z(n202) );
  AND U6645 ( .A(n6693), .B(n6694), .Z(n6692) );
  XNOR U6646 ( .A(n6514), .B(n6691), .Z(n6694) );
  AND U6647 ( .A(p_input[127]), .B(p_input[111]), .Z(n6514) );
  XOR U6648 ( .A(n6691), .B(n6515), .Z(n6693) );
  AND U6649 ( .A(p_input[95]), .B(p_input[79]), .Z(n6515) );
  XOR U6650 ( .A(n6695), .B(n6696), .Z(n6691) );
  AND U6651 ( .A(n6697), .B(n6698), .Z(n6696) );
  XOR U6652 ( .A(n6695), .B(n6525), .Z(n6698) );
  XNOR U6653 ( .A(p_input[110]), .B(n6699), .Z(n6525) );
  AND U6654 ( .A(n298), .B(n6700), .Z(n6699) );
  XOR U6655 ( .A(p_input[126]), .B(p_input[110]), .Z(n6700) );
  XNOR U6656 ( .A(n6522), .B(n6695), .Z(n6697) );
  XOR U6657 ( .A(n6701), .B(n6702), .Z(n6522) );
  AND U6658 ( .A(n296), .B(n6703), .Z(n6702) );
  XOR U6659 ( .A(p_input[94]), .B(p_input[78]), .Z(n6703) );
  XOR U6660 ( .A(n6704), .B(n6705), .Z(n6695) );
  AND U6661 ( .A(n6706), .B(n6707), .Z(n6705) );
  XOR U6662 ( .A(n6704), .B(n6537), .Z(n6707) );
  XNOR U6663 ( .A(p_input[109]), .B(n6708), .Z(n6537) );
  AND U6664 ( .A(n298), .B(n6709), .Z(n6708) );
  XOR U6665 ( .A(p_input[125]), .B(p_input[109]), .Z(n6709) );
  XNOR U6666 ( .A(n6534), .B(n6704), .Z(n6706) );
  XOR U6667 ( .A(n6710), .B(n6711), .Z(n6534) );
  AND U6668 ( .A(n296), .B(n6712), .Z(n6711) );
  XOR U6669 ( .A(p_input[93]), .B(p_input[77]), .Z(n6712) );
  XOR U6670 ( .A(n6713), .B(n6714), .Z(n6704) );
  AND U6671 ( .A(n6715), .B(n6716), .Z(n6714) );
  XOR U6672 ( .A(n6713), .B(n6549), .Z(n6716) );
  XNOR U6673 ( .A(p_input[108]), .B(n6717), .Z(n6549) );
  AND U6674 ( .A(n298), .B(n6718), .Z(n6717) );
  XOR U6675 ( .A(p_input[124]), .B(p_input[108]), .Z(n6718) );
  XNOR U6676 ( .A(n6546), .B(n6713), .Z(n6715) );
  XOR U6677 ( .A(n6719), .B(n6720), .Z(n6546) );
  AND U6678 ( .A(n296), .B(n6721), .Z(n6720) );
  XOR U6679 ( .A(p_input[92]), .B(p_input[76]), .Z(n6721) );
  XOR U6680 ( .A(n6722), .B(n6723), .Z(n6713) );
  AND U6681 ( .A(n6724), .B(n6725), .Z(n6723) );
  XOR U6682 ( .A(n6722), .B(n6561), .Z(n6725) );
  XNOR U6683 ( .A(p_input[107]), .B(n6726), .Z(n6561) );
  AND U6684 ( .A(n298), .B(n6727), .Z(n6726) );
  XOR U6685 ( .A(p_input[123]), .B(p_input[107]), .Z(n6727) );
  XNOR U6686 ( .A(n6558), .B(n6722), .Z(n6724) );
  XOR U6687 ( .A(n6728), .B(n6729), .Z(n6558) );
  AND U6688 ( .A(n296), .B(n6730), .Z(n6729) );
  XOR U6689 ( .A(p_input[91]), .B(p_input[75]), .Z(n6730) );
  XOR U6690 ( .A(n6731), .B(n6732), .Z(n6722) );
  AND U6691 ( .A(n6733), .B(n6734), .Z(n6732) );
  XOR U6692 ( .A(n6731), .B(n6573), .Z(n6734) );
  XNOR U6693 ( .A(p_input[106]), .B(n6735), .Z(n6573) );
  AND U6694 ( .A(n298), .B(n6736), .Z(n6735) );
  XOR U6695 ( .A(p_input[122]), .B(p_input[106]), .Z(n6736) );
  XNOR U6696 ( .A(n6570), .B(n6731), .Z(n6733) );
  XOR U6697 ( .A(n6737), .B(n6738), .Z(n6570) );
  AND U6698 ( .A(n296), .B(n6739), .Z(n6738) );
  XOR U6699 ( .A(p_input[90]), .B(p_input[74]), .Z(n6739) );
  XOR U6700 ( .A(n6740), .B(n6741), .Z(n6731) );
  AND U6701 ( .A(n6742), .B(n6743), .Z(n6741) );
  XOR U6702 ( .A(n6740), .B(n6585), .Z(n6743) );
  XNOR U6703 ( .A(p_input[105]), .B(n6744), .Z(n6585) );
  AND U6704 ( .A(n298), .B(n6745), .Z(n6744) );
  XOR U6705 ( .A(p_input[121]), .B(p_input[105]), .Z(n6745) );
  XNOR U6706 ( .A(n6582), .B(n6740), .Z(n6742) );
  XOR U6707 ( .A(n6746), .B(n6747), .Z(n6582) );
  AND U6708 ( .A(n296), .B(n6748), .Z(n6747) );
  XOR U6709 ( .A(p_input[89]), .B(p_input[73]), .Z(n6748) );
  XOR U6710 ( .A(n6749), .B(n6750), .Z(n6740) );
  AND U6711 ( .A(n6751), .B(n6752), .Z(n6750) );
  XOR U6712 ( .A(n6749), .B(n6597), .Z(n6752) );
  XNOR U6713 ( .A(p_input[104]), .B(n6753), .Z(n6597) );
  AND U6714 ( .A(n298), .B(n6754), .Z(n6753) );
  XOR U6715 ( .A(p_input[120]), .B(p_input[104]), .Z(n6754) );
  XNOR U6716 ( .A(n6594), .B(n6749), .Z(n6751) );
  XOR U6717 ( .A(n6755), .B(n6756), .Z(n6594) );
  AND U6718 ( .A(n296), .B(n6757), .Z(n6756) );
  XOR U6719 ( .A(p_input[88]), .B(p_input[72]), .Z(n6757) );
  XOR U6720 ( .A(n6758), .B(n6759), .Z(n6749) );
  AND U6721 ( .A(n6760), .B(n6761), .Z(n6759) );
  XOR U6722 ( .A(n6758), .B(n6609), .Z(n6761) );
  XNOR U6723 ( .A(p_input[103]), .B(n6762), .Z(n6609) );
  AND U6724 ( .A(n298), .B(n6763), .Z(n6762) );
  XOR U6725 ( .A(p_input[119]), .B(p_input[103]), .Z(n6763) );
  XNOR U6726 ( .A(n6606), .B(n6758), .Z(n6760) );
  XOR U6727 ( .A(n6764), .B(n6765), .Z(n6606) );
  AND U6728 ( .A(n296), .B(n6766), .Z(n6765) );
  XOR U6729 ( .A(p_input[87]), .B(p_input[71]), .Z(n6766) );
  XOR U6730 ( .A(n6767), .B(n6768), .Z(n6758) );
  AND U6731 ( .A(n6769), .B(n6770), .Z(n6768) );
  XOR U6732 ( .A(n6767), .B(n6621), .Z(n6770) );
  XNOR U6733 ( .A(p_input[102]), .B(n6771), .Z(n6621) );
  AND U6734 ( .A(n298), .B(n6772), .Z(n6771) );
  XOR U6735 ( .A(p_input[118]), .B(p_input[102]), .Z(n6772) );
  XNOR U6736 ( .A(n6618), .B(n6767), .Z(n6769) );
  XOR U6737 ( .A(n6773), .B(n6774), .Z(n6618) );
  AND U6738 ( .A(n296), .B(n6775), .Z(n6774) );
  XOR U6739 ( .A(p_input[86]), .B(p_input[70]), .Z(n6775) );
  XOR U6740 ( .A(n6776), .B(n6777), .Z(n6767) );
  AND U6741 ( .A(n6778), .B(n6779), .Z(n6777) );
  XOR U6742 ( .A(n6776), .B(n6633), .Z(n6779) );
  XNOR U6743 ( .A(p_input[101]), .B(n6780), .Z(n6633) );
  AND U6744 ( .A(n298), .B(n6781), .Z(n6780) );
  XOR U6745 ( .A(p_input[117]), .B(p_input[101]), .Z(n6781) );
  XNOR U6746 ( .A(n6630), .B(n6776), .Z(n6778) );
  XOR U6747 ( .A(n6782), .B(n6783), .Z(n6630) );
  AND U6748 ( .A(n296), .B(n6784), .Z(n6783) );
  XOR U6749 ( .A(p_input[85]), .B(p_input[69]), .Z(n6784) );
  XOR U6750 ( .A(n6785), .B(n6786), .Z(n6776) );
  AND U6751 ( .A(n6787), .B(n6788), .Z(n6786) );
  XOR U6752 ( .A(n6785), .B(n6645), .Z(n6788) );
  XNOR U6753 ( .A(p_input[100]), .B(n6789), .Z(n6645) );
  AND U6754 ( .A(n298), .B(n6790), .Z(n6789) );
  XOR U6755 ( .A(p_input[116]), .B(p_input[100]), .Z(n6790) );
  XNOR U6756 ( .A(n6642), .B(n6785), .Z(n6787) );
  XOR U6757 ( .A(n6791), .B(n6792), .Z(n6642) );
  AND U6758 ( .A(n296), .B(n6793), .Z(n6792) );
  XOR U6759 ( .A(p_input[84]), .B(p_input[68]), .Z(n6793) );
  XOR U6760 ( .A(n6794), .B(n6795), .Z(n6785) );
  AND U6761 ( .A(n6796), .B(n6797), .Z(n6795) );
  XOR U6762 ( .A(n6657), .B(n6794), .Z(n6797) );
  XNOR U6763 ( .A(p_input[99]), .B(n6798), .Z(n6657) );
  AND U6764 ( .A(n298), .B(n6799), .Z(n6798) );
  XOR U6765 ( .A(p_input[99]), .B(p_input[115]), .Z(n6799) );
  XNOR U6766 ( .A(n6794), .B(n6654), .Z(n6796) );
  XOR U6767 ( .A(n6800), .B(n6801), .Z(n6654) );
  AND U6768 ( .A(n296), .B(n6802), .Z(n6801) );
  XOR U6769 ( .A(p_input[83]), .B(p_input[67]), .Z(n6802) );
  XOR U6770 ( .A(n6803), .B(n6804), .Z(n6794) );
  AND U6771 ( .A(n6805), .B(n6806), .Z(n6804) );
  XOR U6772 ( .A(n6803), .B(n6669), .Z(n6806) );
  XNOR U6773 ( .A(p_input[98]), .B(n6807), .Z(n6669) );
  AND U6774 ( .A(n298), .B(n6808), .Z(n6807) );
  XOR U6775 ( .A(p_input[98]), .B(p_input[114]), .Z(n6808) );
  XNOR U6776 ( .A(n6666), .B(n6803), .Z(n6805) );
  XOR U6777 ( .A(n6809), .B(n6810), .Z(n6666) );
  AND U6778 ( .A(n296), .B(n6811), .Z(n6810) );
  XOR U6779 ( .A(p_input[82]), .B(p_input[66]), .Z(n6811) );
  XOR U6780 ( .A(n6812), .B(n6813), .Z(n6803) );
  AND U6781 ( .A(n6814), .B(n6815), .Z(n6813) );
  XNOR U6782 ( .A(n6816), .B(n6682), .Z(n6815) );
  XNOR U6783 ( .A(p_input[97]), .B(n6817), .Z(n6682) );
  AND U6784 ( .A(n298), .B(n6818), .Z(n6817) );
  XNOR U6785 ( .A(n6819), .B(p_input[113]), .Z(n6818) );
  IV U6786 ( .A(p_input[97]), .Z(n6819) );
  XNOR U6787 ( .A(n6679), .B(n6812), .Z(n6814) );
  XNOR U6788 ( .A(p_input[65]), .B(n6820), .Z(n6679) );
  AND U6789 ( .A(n296), .B(n6821), .Z(n6820) );
  XOR U6790 ( .A(p_input[81]), .B(p_input[65]), .Z(n6821) );
  IV U6791 ( .A(n6816), .Z(n6812) );
  AND U6792 ( .A(n6687), .B(n6690), .Z(n6816) );
  XOR U6793 ( .A(p_input[96]), .B(n6822), .Z(n6690) );
  AND U6794 ( .A(n298), .B(n6823), .Z(n6822) );
  XOR U6795 ( .A(p_input[96]), .B(p_input[112]), .Z(n6823) );
  XOR U6796 ( .A(n6824), .B(n6825), .Z(n298) );
  AND U6797 ( .A(n6826), .B(n6827), .Z(n6825) );
  XNOR U6798 ( .A(p_input[127]), .B(n6824), .Z(n6827) );
  XOR U6799 ( .A(n6824), .B(p_input[111]), .Z(n6826) );
  XOR U6800 ( .A(n6828), .B(n6829), .Z(n6824) );
  AND U6801 ( .A(n6830), .B(n6831), .Z(n6829) );
  XNOR U6802 ( .A(p_input[126]), .B(n6828), .Z(n6831) );
  XOR U6803 ( .A(n6828), .B(p_input[110]), .Z(n6830) );
  XOR U6804 ( .A(n6832), .B(n6833), .Z(n6828) );
  AND U6805 ( .A(n6834), .B(n6835), .Z(n6833) );
  XNOR U6806 ( .A(p_input[125]), .B(n6832), .Z(n6835) );
  XOR U6807 ( .A(n6832), .B(p_input[109]), .Z(n6834) );
  XOR U6808 ( .A(n6836), .B(n6837), .Z(n6832) );
  AND U6809 ( .A(n6838), .B(n6839), .Z(n6837) );
  XNOR U6810 ( .A(p_input[124]), .B(n6836), .Z(n6839) );
  XOR U6811 ( .A(n6836), .B(p_input[108]), .Z(n6838) );
  XOR U6812 ( .A(n6840), .B(n6841), .Z(n6836) );
  AND U6813 ( .A(n6842), .B(n6843), .Z(n6841) );
  XNOR U6814 ( .A(p_input[123]), .B(n6840), .Z(n6843) );
  XOR U6815 ( .A(n6840), .B(p_input[107]), .Z(n6842) );
  XOR U6816 ( .A(n6844), .B(n6845), .Z(n6840) );
  AND U6817 ( .A(n6846), .B(n6847), .Z(n6845) );
  XNOR U6818 ( .A(p_input[122]), .B(n6844), .Z(n6847) );
  XOR U6819 ( .A(n6844), .B(p_input[106]), .Z(n6846) );
  XOR U6820 ( .A(n6848), .B(n6849), .Z(n6844) );
  AND U6821 ( .A(n6850), .B(n6851), .Z(n6849) );
  XNOR U6822 ( .A(p_input[121]), .B(n6848), .Z(n6851) );
  XOR U6823 ( .A(n6848), .B(p_input[105]), .Z(n6850) );
  XOR U6824 ( .A(n6852), .B(n6853), .Z(n6848) );
  AND U6825 ( .A(n6854), .B(n6855), .Z(n6853) );
  XNOR U6826 ( .A(p_input[120]), .B(n6852), .Z(n6855) );
  XOR U6827 ( .A(n6852), .B(p_input[104]), .Z(n6854) );
  XOR U6828 ( .A(n6856), .B(n6857), .Z(n6852) );
  AND U6829 ( .A(n6858), .B(n6859), .Z(n6857) );
  XNOR U6830 ( .A(p_input[119]), .B(n6856), .Z(n6859) );
  XOR U6831 ( .A(n6856), .B(p_input[103]), .Z(n6858) );
  XOR U6832 ( .A(n6860), .B(n6861), .Z(n6856) );
  AND U6833 ( .A(n6862), .B(n6863), .Z(n6861) );
  XNOR U6834 ( .A(p_input[118]), .B(n6860), .Z(n6863) );
  XOR U6835 ( .A(n6860), .B(p_input[102]), .Z(n6862) );
  XOR U6836 ( .A(n6864), .B(n6865), .Z(n6860) );
  AND U6837 ( .A(n6866), .B(n6867), .Z(n6865) );
  XNOR U6838 ( .A(p_input[117]), .B(n6864), .Z(n6867) );
  XOR U6839 ( .A(n6864), .B(p_input[101]), .Z(n6866) );
  XOR U6840 ( .A(n6868), .B(n6869), .Z(n6864) );
  AND U6841 ( .A(n6870), .B(n6871), .Z(n6869) );
  XNOR U6842 ( .A(p_input[116]), .B(n6868), .Z(n6871) );
  XOR U6843 ( .A(n6868), .B(p_input[100]), .Z(n6870) );
  XOR U6844 ( .A(n6872), .B(n6873), .Z(n6868) );
  AND U6845 ( .A(n6874), .B(n6875), .Z(n6873) );
  XNOR U6846 ( .A(p_input[115]), .B(n6872), .Z(n6875) );
  XOR U6847 ( .A(n6872), .B(p_input[99]), .Z(n6874) );
  XOR U6848 ( .A(n6876), .B(n6877), .Z(n6872) );
  AND U6849 ( .A(n6878), .B(n6879), .Z(n6877) );
  XNOR U6850 ( .A(p_input[114]), .B(n6876), .Z(n6879) );
  XOR U6851 ( .A(n6876), .B(p_input[98]), .Z(n6878) );
  XNOR U6852 ( .A(n6880), .B(n6881), .Z(n6876) );
  AND U6853 ( .A(n6882), .B(n6883), .Z(n6881) );
  XOR U6854 ( .A(p_input[113]), .B(n6880), .Z(n6883) );
  XNOR U6855 ( .A(p_input[97]), .B(n6880), .Z(n6882) );
  AND U6856 ( .A(p_input[112]), .B(n6884), .Z(n6880) );
  IV U6857 ( .A(p_input[96]), .Z(n6884) );
  XNOR U6858 ( .A(p_input[64]), .B(n6885), .Z(n6687) );
  AND U6859 ( .A(n296), .B(n6886), .Z(n6885) );
  XOR U6860 ( .A(p_input[80]), .B(p_input[64]), .Z(n6886) );
  XOR U6861 ( .A(n6887), .B(n6888), .Z(n296) );
  AND U6862 ( .A(n6889), .B(n6890), .Z(n6888) );
  XNOR U6863 ( .A(p_input[95]), .B(n6887), .Z(n6890) );
  XOR U6864 ( .A(n6887), .B(p_input[79]), .Z(n6889) );
  XOR U6865 ( .A(n6891), .B(n6892), .Z(n6887) );
  AND U6866 ( .A(n6893), .B(n6894), .Z(n6892) );
  XNOR U6867 ( .A(p_input[94]), .B(n6891), .Z(n6894) );
  XNOR U6868 ( .A(n6891), .B(n6701), .Z(n6893) );
  IV U6869 ( .A(p_input[78]), .Z(n6701) );
  XOR U6870 ( .A(n6895), .B(n6896), .Z(n6891) );
  AND U6871 ( .A(n6897), .B(n6898), .Z(n6896) );
  XNOR U6872 ( .A(p_input[93]), .B(n6895), .Z(n6898) );
  XNOR U6873 ( .A(n6895), .B(n6710), .Z(n6897) );
  IV U6874 ( .A(p_input[77]), .Z(n6710) );
  XOR U6875 ( .A(n6899), .B(n6900), .Z(n6895) );
  AND U6876 ( .A(n6901), .B(n6902), .Z(n6900) );
  XNOR U6877 ( .A(p_input[92]), .B(n6899), .Z(n6902) );
  XNOR U6878 ( .A(n6899), .B(n6719), .Z(n6901) );
  IV U6879 ( .A(p_input[76]), .Z(n6719) );
  XOR U6880 ( .A(n6903), .B(n6904), .Z(n6899) );
  AND U6881 ( .A(n6905), .B(n6906), .Z(n6904) );
  XNOR U6882 ( .A(p_input[91]), .B(n6903), .Z(n6906) );
  XNOR U6883 ( .A(n6903), .B(n6728), .Z(n6905) );
  IV U6884 ( .A(p_input[75]), .Z(n6728) );
  XOR U6885 ( .A(n6907), .B(n6908), .Z(n6903) );
  AND U6886 ( .A(n6909), .B(n6910), .Z(n6908) );
  XNOR U6887 ( .A(p_input[90]), .B(n6907), .Z(n6910) );
  XNOR U6888 ( .A(n6907), .B(n6737), .Z(n6909) );
  IV U6889 ( .A(p_input[74]), .Z(n6737) );
  XOR U6890 ( .A(n6911), .B(n6912), .Z(n6907) );
  AND U6891 ( .A(n6913), .B(n6914), .Z(n6912) );
  XNOR U6892 ( .A(p_input[89]), .B(n6911), .Z(n6914) );
  XNOR U6893 ( .A(n6911), .B(n6746), .Z(n6913) );
  IV U6894 ( .A(p_input[73]), .Z(n6746) );
  XOR U6895 ( .A(n6915), .B(n6916), .Z(n6911) );
  AND U6896 ( .A(n6917), .B(n6918), .Z(n6916) );
  XNOR U6897 ( .A(p_input[88]), .B(n6915), .Z(n6918) );
  XNOR U6898 ( .A(n6915), .B(n6755), .Z(n6917) );
  IV U6899 ( .A(p_input[72]), .Z(n6755) );
  XOR U6900 ( .A(n6919), .B(n6920), .Z(n6915) );
  AND U6901 ( .A(n6921), .B(n6922), .Z(n6920) );
  XNOR U6902 ( .A(p_input[87]), .B(n6919), .Z(n6922) );
  XNOR U6903 ( .A(n6919), .B(n6764), .Z(n6921) );
  IV U6904 ( .A(p_input[71]), .Z(n6764) );
  XOR U6905 ( .A(n6923), .B(n6924), .Z(n6919) );
  AND U6906 ( .A(n6925), .B(n6926), .Z(n6924) );
  XNOR U6907 ( .A(p_input[86]), .B(n6923), .Z(n6926) );
  XNOR U6908 ( .A(n6923), .B(n6773), .Z(n6925) );
  IV U6909 ( .A(p_input[70]), .Z(n6773) );
  XOR U6910 ( .A(n6927), .B(n6928), .Z(n6923) );
  AND U6911 ( .A(n6929), .B(n6930), .Z(n6928) );
  XNOR U6912 ( .A(p_input[85]), .B(n6927), .Z(n6930) );
  XNOR U6913 ( .A(n6927), .B(n6782), .Z(n6929) );
  IV U6914 ( .A(p_input[69]), .Z(n6782) );
  XOR U6915 ( .A(n6931), .B(n6932), .Z(n6927) );
  AND U6916 ( .A(n6933), .B(n6934), .Z(n6932) );
  XNOR U6917 ( .A(p_input[84]), .B(n6931), .Z(n6934) );
  XNOR U6918 ( .A(n6931), .B(n6791), .Z(n6933) );
  IV U6919 ( .A(p_input[68]), .Z(n6791) );
  XOR U6920 ( .A(n6935), .B(n6936), .Z(n6931) );
  AND U6921 ( .A(n6937), .B(n6938), .Z(n6936) );
  XNOR U6922 ( .A(p_input[83]), .B(n6935), .Z(n6938) );
  XNOR U6923 ( .A(n6935), .B(n6800), .Z(n6937) );
  IV U6924 ( .A(p_input[67]), .Z(n6800) );
  XOR U6925 ( .A(n6939), .B(n6940), .Z(n6935) );
  AND U6926 ( .A(n6941), .B(n6942), .Z(n6940) );
  XNOR U6927 ( .A(p_input[82]), .B(n6939), .Z(n6942) );
  XNOR U6928 ( .A(n6939), .B(n6809), .Z(n6941) );
  IV U6929 ( .A(p_input[66]), .Z(n6809) );
  XNOR U6930 ( .A(n6943), .B(n6944), .Z(n6939) );
  AND U6931 ( .A(n6945), .B(n6946), .Z(n6944) );
  XOR U6932 ( .A(p_input[81]), .B(n6943), .Z(n6946) );
  XNOR U6933 ( .A(p_input[65]), .B(n6943), .Z(n6945) );
  AND U6934 ( .A(p_input[80]), .B(n6947), .Z(n6943) );
  IV U6935 ( .A(p_input[64]), .Z(n6947) );
  XOR U6936 ( .A(n6948), .B(n6949), .Z(n6506) );
  AND U6937 ( .A(n199), .B(n6950), .Z(n6949) );
  XNOR U6938 ( .A(n6951), .B(n6948), .Z(n6950) );
  XOR U6939 ( .A(n6952), .B(n6953), .Z(n199) );
  AND U6940 ( .A(n6954), .B(n6955), .Z(n6953) );
  XNOR U6941 ( .A(n6517), .B(n6952), .Z(n6955) );
  AND U6942 ( .A(p_input[63]), .B(p_input[47]), .Z(n6517) );
  XOR U6943 ( .A(n6952), .B(n6516), .Z(n6954) );
  AND U6944 ( .A(p_input[15]), .B(p_input[31]), .Z(n6516) );
  XOR U6945 ( .A(n6956), .B(n6957), .Z(n6952) );
  AND U6946 ( .A(n6958), .B(n6959), .Z(n6957) );
  XOR U6947 ( .A(n6956), .B(n6529), .Z(n6959) );
  XNOR U6948 ( .A(p_input[46]), .B(n6960), .Z(n6529) );
  AND U6949 ( .A(n306), .B(n6961), .Z(n6960) );
  XOR U6950 ( .A(p_input[62]), .B(p_input[46]), .Z(n6961) );
  XNOR U6951 ( .A(n6526), .B(n6956), .Z(n6958) );
  XOR U6952 ( .A(n6962), .B(n6963), .Z(n6526) );
  AND U6953 ( .A(n303), .B(n6964), .Z(n6963) );
  XOR U6954 ( .A(p_input[30]), .B(p_input[14]), .Z(n6964) );
  XOR U6955 ( .A(n6965), .B(n6966), .Z(n6956) );
  AND U6956 ( .A(n6967), .B(n6968), .Z(n6966) );
  XOR U6957 ( .A(n6965), .B(n6541), .Z(n6968) );
  XNOR U6958 ( .A(p_input[45]), .B(n6969), .Z(n6541) );
  AND U6959 ( .A(n306), .B(n6970), .Z(n6969) );
  XOR U6960 ( .A(p_input[61]), .B(p_input[45]), .Z(n6970) );
  XNOR U6961 ( .A(n6538), .B(n6965), .Z(n6967) );
  XOR U6962 ( .A(n6971), .B(n6972), .Z(n6538) );
  AND U6963 ( .A(n303), .B(n6973), .Z(n6972) );
  XOR U6964 ( .A(p_input[29]), .B(p_input[13]), .Z(n6973) );
  XOR U6965 ( .A(n6974), .B(n6975), .Z(n6965) );
  AND U6966 ( .A(n6976), .B(n6977), .Z(n6975) );
  XOR U6967 ( .A(n6974), .B(n6553), .Z(n6977) );
  XNOR U6968 ( .A(p_input[44]), .B(n6978), .Z(n6553) );
  AND U6969 ( .A(n306), .B(n6979), .Z(n6978) );
  XOR U6970 ( .A(p_input[60]), .B(p_input[44]), .Z(n6979) );
  XNOR U6971 ( .A(n6550), .B(n6974), .Z(n6976) );
  XOR U6972 ( .A(n6980), .B(n6981), .Z(n6550) );
  AND U6973 ( .A(n303), .B(n6982), .Z(n6981) );
  XOR U6974 ( .A(p_input[28]), .B(p_input[12]), .Z(n6982) );
  XOR U6975 ( .A(n6983), .B(n6984), .Z(n6974) );
  AND U6976 ( .A(n6985), .B(n6986), .Z(n6984) );
  XOR U6977 ( .A(n6983), .B(n6565), .Z(n6986) );
  XNOR U6978 ( .A(p_input[43]), .B(n6987), .Z(n6565) );
  AND U6979 ( .A(n306), .B(n6988), .Z(n6987) );
  XOR U6980 ( .A(p_input[59]), .B(p_input[43]), .Z(n6988) );
  XNOR U6981 ( .A(n6562), .B(n6983), .Z(n6985) );
  XOR U6982 ( .A(n6989), .B(n6990), .Z(n6562) );
  AND U6983 ( .A(n303), .B(n6991), .Z(n6990) );
  XOR U6984 ( .A(p_input[27]), .B(p_input[11]), .Z(n6991) );
  XOR U6985 ( .A(n6992), .B(n6993), .Z(n6983) );
  AND U6986 ( .A(n6994), .B(n6995), .Z(n6993) );
  XOR U6987 ( .A(n6992), .B(n6577), .Z(n6995) );
  XNOR U6988 ( .A(p_input[42]), .B(n6996), .Z(n6577) );
  AND U6989 ( .A(n306), .B(n6997), .Z(n6996) );
  XOR U6990 ( .A(p_input[58]), .B(p_input[42]), .Z(n6997) );
  XNOR U6991 ( .A(n6574), .B(n6992), .Z(n6994) );
  XOR U6992 ( .A(n6998), .B(n6999), .Z(n6574) );
  AND U6993 ( .A(n303), .B(n7000), .Z(n6999) );
  XOR U6994 ( .A(p_input[26]), .B(p_input[10]), .Z(n7000) );
  XOR U6995 ( .A(n7001), .B(n7002), .Z(n6992) );
  AND U6996 ( .A(n7003), .B(n7004), .Z(n7002) );
  XOR U6997 ( .A(n7001), .B(n6589), .Z(n7004) );
  XNOR U6998 ( .A(p_input[41]), .B(n7005), .Z(n6589) );
  AND U6999 ( .A(n306), .B(n7006), .Z(n7005) );
  XOR U7000 ( .A(p_input[57]), .B(p_input[41]), .Z(n7006) );
  XNOR U7001 ( .A(n6586), .B(n7001), .Z(n7003) );
  XOR U7002 ( .A(n7007), .B(n7008), .Z(n6586) );
  AND U7003 ( .A(n303), .B(n7009), .Z(n7008) );
  XOR U7004 ( .A(p_input[9]), .B(p_input[25]), .Z(n7009) );
  XOR U7005 ( .A(n7010), .B(n7011), .Z(n7001) );
  AND U7006 ( .A(n7012), .B(n7013), .Z(n7011) );
  XOR U7007 ( .A(n7010), .B(n6601), .Z(n7013) );
  XNOR U7008 ( .A(p_input[40]), .B(n7014), .Z(n6601) );
  AND U7009 ( .A(n306), .B(n7015), .Z(n7014) );
  XOR U7010 ( .A(p_input[56]), .B(p_input[40]), .Z(n7015) );
  XNOR U7011 ( .A(n6598), .B(n7010), .Z(n7012) );
  XOR U7012 ( .A(n7016), .B(n7017), .Z(n6598) );
  AND U7013 ( .A(n303), .B(n7018), .Z(n7017) );
  XOR U7014 ( .A(p_input[8]), .B(p_input[24]), .Z(n7018) );
  XOR U7015 ( .A(n7019), .B(n7020), .Z(n7010) );
  AND U7016 ( .A(n7021), .B(n7022), .Z(n7020) );
  XOR U7017 ( .A(n7019), .B(n6613), .Z(n7022) );
  XNOR U7018 ( .A(p_input[39]), .B(n7023), .Z(n6613) );
  AND U7019 ( .A(n306), .B(n7024), .Z(n7023) );
  XOR U7020 ( .A(p_input[55]), .B(p_input[39]), .Z(n7024) );
  XNOR U7021 ( .A(n6610), .B(n7019), .Z(n7021) );
  XOR U7022 ( .A(n7025), .B(n7026), .Z(n6610) );
  AND U7023 ( .A(n303), .B(n7027), .Z(n7026) );
  XOR U7024 ( .A(p_input[7]), .B(p_input[23]), .Z(n7027) );
  XOR U7025 ( .A(n7028), .B(n7029), .Z(n7019) );
  AND U7026 ( .A(n7030), .B(n7031), .Z(n7029) );
  XOR U7027 ( .A(n7028), .B(n6625), .Z(n7031) );
  XNOR U7028 ( .A(p_input[38]), .B(n7032), .Z(n6625) );
  AND U7029 ( .A(n306), .B(n7033), .Z(n7032) );
  XOR U7030 ( .A(p_input[54]), .B(p_input[38]), .Z(n7033) );
  XNOR U7031 ( .A(n6622), .B(n7028), .Z(n7030) );
  XOR U7032 ( .A(n7034), .B(n7035), .Z(n6622) );
  AND U7033 ( .A(n303), .B(n7036), .Z(n7035) );
  XOR U7034 ( .A(p_input[6]), .B(p_input[22]), .Z(n7036) );
  XOR U7035 ( .A(n7037), .B(n7038), .Z(n7028) );
  AND U7036 ( .A(n7039), .B(n7040), .Z(n7038) );
  XOR U7037 ( .A(n7037), .B(n6637), .Z(n7040) );
  XNOR U7038 ( .A(p_input[37]), .B(n7041), .Z(n6637) );
  AND U7039 ( .A(n306), .B(n7042), .Z(n7041) );
  XOR U7040 ( .A(p_input[53]), .B(p_input[37]), .Z(n7042) );
  XNOR U7041 ( .A(n6634), .B(n7037), .Z(n7039) );
  XOR U7042 ( .A(n7043), .B(n7044), .Z(n6634) );
  AND U7043 ( .A(n303), .B(n7045), .Z(n7044) );
  XOR U7044 ( .A(p_input[5]), .B(p_input[21]), .Z(n7045) );
  XOR U7045 ( .A(n7046), .B(n7047), .Z(n7037) );
  AND U7046 ( .A(n7048), .B(n7049), .Z(n7047) );
  XOR U7047 ( .A(n7046), .B(n6649), .Z(n7049) );
  XNOR U7048 ( .A(p_input[36]), .B(n7050), .Z(n6649) );
  AND U7049 ( .A(n306), .B(n7051), .Z(n7050) );
  XOR U7050 ( .A(p_input[52]), .B(p_input[36]), .Z(n7051) );
  XNOR U7051 ( .A(n6646), .B(n7046), .Z(n7048) );
  XOR U7052 ( .A(n7052), .B(n7053), .Z(n6646) );
  AND U7053 ( .A(n303), .B(n7054), .Z(n7053) );
  XOR U7054 ( .A(p_input[4]), .B(p_input[20]), .Z(n7054) );
  XOR U7055 ( .A(n7055), .B(n7056), .Z(n7046) );
  AND U7056 ( .A(n7057), .B(n7058), .Z(n7056) );
  XOR U7057 ( .A(n6661), .B(n7055), .Z(n7058) );
  XNOR U7058 ( .A(p_input[35]), .B(n7059), .Z(n6661) );
  AND U7059 ( .A(n306), .B(n7060), .Z(n7059) );
  XOR U7060 ( .A(p_input[51]), .B(p_input[35]), .Z(n7060) );
  XNOR U7061 ( .A(n7055), .B(n6658), .Z(n7057) );
  XOR U7062 ( .A(n7061), .B(n7062), .Z(n6658) );
  AND U7063 ( .A(n303), .B(n7063), .Z(n7062) );
  XOR U7064 ( .A(p_input[3]), .B(p_input[19]), .Z(n7063) );
  XOR U7065 ( .A(n7064), .B(n7065), .Z(n7055) );
  AND U7066 ( .A(n7066), .B(n7067), .Z(n7065) );
  XOR U7067 ( .A(n7064), .B(n6673), .Z(n7067) );
  XNOR U7068 ( .A(p_input[34]), .B(n7068), .Z(n6673) );
  AND U7069 ( .A(n306), .B(n7069), .Z(n7068) );
  XOR U7070 ( .A(p_input[50]), .B(p_input[34]), .Z(n7069) );
  XNOR U7071 ( .A(n6670), .B(n7064), .Z(n7066) );
  XOR U7072 ( .A(n7070), .B(n7071), .Z(n6670) );
  AND U7073 ( .A(n303), .B(n7072), .Z(n7071) );
  XOR U7074 ( .A(p_input[2]), .B(p_input[18]), .Z(n7072) );
  XOR U7075 ( .A(n7073), .B(n7074), .Z(n7064) );
  AND U7076 ( .A(n7075), .B(n7076), .Z(n7074) );
  XNOR U7077 ( .A(n7077), .B(n6686), .Z(n7076) );
  XNOR U7078 ( .A(p_input[33]), .B(n7078), .Z(n6686) );
  AND U7079 ( .A(n306), .B(n7079), .Z(n7078) );
  XNOR U7080 ( .A(p_input[49]), .B(n7080), .Z(n7079) );
  IV U7081 ( .A(p_input[33]), .Z(n7080) );
  XNOR U7082 ( .A(n6683), .B(n7073), .Z(n7075) );
  XNOR U7083 ( .A(p_input[1]), .B(n7081), .Z(n6683) );
  AND U7084 ( .A(n303), .B(n7082), .Z(n7081) );
  XOR U7085 ( .A(p_input[1]), .B(p_input[17]), .Z(n7082) );
  IV U7086 ( .A(n7077), .Z(n7073) );
  AND U7087 ( .A(n6948), .B(n6951), .Z(n7077) );
  XOR U7088 ( .A(p_input[32]), .B(n7083), .Z(n6951) );
  AND U7089 ( .A(n306), .B(n7084), .Z(n7083) );
  XOR U7090 ( .A(p_input[48]), .B(p_input[32]), .Z(n7084) );
  XOR U7091 ( .A(n7085), .B(n7086), .Z(n306) );
  AND U7092 ( .A(n7087), .B(n7088), .Z(n7086) );
  XNOR U7093 ( .A(p_input[63]), .B(n7085), .Z(n7088) );
  XOR U7094 ( .A(n7085), .B(p_input[47]), .Z(n7087) );
  XOR U7095 ( .A(n7089), .B(n7090), .Z(n7085) );
  AND U7096 ( .A(n7091), .B(n7092), .Z(n7090) );
  XNOR U7097 ( .A(p_input[62]), .B(n7089), .Z(n7092) );
  XOR U7098 ( .A(n7089), .B(p_input[46]), .Z(n7091) );
  XOR U7099 ( .A(n7093), .B(n7094), .Z(n7089) );
  AND U7100 ( .A(n7095), .B(n7096), .Z(n7094) );
  XNOR U7101 ( .A(p_input[61]), .B(n7093), .Z(n7096) );
  XOR U7102 ( .A(n7093), .B(p_input[45]), .Z(n7095) );
  XOR U7103 ( .A(n7097), .B(n7098), .Z(n7093) );
  AND U7104 ( .A(n7099), .B(n7100), .Z(n7098) );
  XNOR U7105 ( .A(p_input[60]), .B(n7097), .Z(n7100) );
  XOR U7106 ( .A(n7097), .B(p_input[44]), .Z(n7099) );
  XOR U7107 ( .A(n7101), .B(n7102), .Z(n7097) );
  AND U7108 ( .A(n7103), .B(n7104), .Z(n7102) );
  XNOR U7109 ( .A(p_input[59]), .B(n7101), .Z(n7104) );
  XOR U7110 ( .A(n7101), .B(p_input[43]), .Z(n7103) );
  XOR U7111 ( .A(n7105), .B(n7106), .Z(n7101) );
  AND U7112 ( .A(n7107), .B(n7108), .Z(n7106) );
  XNOR U7113 ( .A(p_input[58]), .B(n7105), .Z(n7108) );
  XOR U7114 ( .A(n7105), .B(p_input[42]), .Z(n7107) );
  XOR U7115 ( .A(n7109), .B(n7110), .Z(n7105) );
  AND U7116 ( .A(n7111), .B(n7112), .Z(n7110) );
  XNOR U7117 ( .A(p_input[57]), .B(n7109), .Z(n7112) );
  XOR U7118 ( .A(n7109), .B(p_input[41]), .Z(n7111) );
  XOR U7119 ( .A(n7113), .B(n7114), .Z(n7109) );
  AND U7120 ( .A(n7115), .B(n7116), .Z(n7114) );
  XNOR U7121 ( .A(p_input[56]), .B(n7113), .Z(n7116) );
  XOR U7122 ( .A(n7113), .B(p_input[40]), .Z(n7115) );
  XOR U7123 ( .A(n7117), .B(n7118), .Z(n7113) );
  AND U7124 ( .A(n7119), .B(n7120), .Z(n7118) );
  XNOR U7125 ( .A(p_input[55]), .B(n7117), .Z(n7120) );
  XOR U7126 ( .A(n7117), .B(p_input[39]), .Z(n7119) );
  XOR U7127 ( .A(n7121), .B(n7122), .Z(n7117) );
  AND U7128 ( .A(n7123), .B(n7124), .Z(n7122) );
  XNOR U7129 ( .A(p_input[54]), .B(n7121), .Z(n7124) );
  XOR U7130 ( .A(n7121), .B(p_input[38]), .Z(n7123) );
  XOR U7131 ( .A(n7125), .B(n7126), .Z(n7121) );
  AND U7132 ( .A(n7127), .B(n7128), .Z(n7126) );
  XNOR U7133 ( .A(p_input[53]), .B(n7125), .Z(n7128) );
  XOR U7134 ( .A(n7125), .B(p_input[37]), .Z(n7127) );
  XOR U7135 ( .A(n7129), .B(n7130), .Z(n7125) );
  AND U7136 ( .A(n7131), .B(n7132), .Z(n7130) );
  XNOR U7137 ( .A(p_input[52]), .B(n7129), .Z(n7132) );
  XOR U7138 ( .A(n7129), .B(p_input[36]), .Z(n7131) );
  XOR U7139 ( .A(n7133), .B(n7134), .Z(n7129) );
  AND U7140 ( .A(n7135), .B(n7136), .Z(n7134) );
  XNOR U7141 ( .A(p_input[51]), .B(n7133), .Z(n7136) );
  XOR U7142 ( .A(n7133), .B(p_input[35]), .Z(n7135) );
  XOR U7143 ( .A(n7137), .B(n7138), .Z(n7133) );
  AND U7144 ( .A(n7139), .B(n7140), .Z(n7138) );
  XNOR U7145 ( .A(p_input[50]), .B(n7137), .Z(n7140) );
  XOR U7146 ( .A(n7137), .B(p_input[34]), .Z(n7139) );
  XNOR U7147 ( .A(n7141), .B(n7142), .Z(n7137) );
  AND U7148 ( .A(n7143), .B(n7144), .Z(n7142) );
  XOR U7149 ( .A(p_input[49]), .B(n7141), .Z(n7144) );
  XNOR U7150 ( .A(p_input[33]), .B(n7141), .Z(n7143) );
  AND U7151 ( .A(p_input[48]), .B(n7145), .Z(n7141) );
  IV U7152 ( .A(p_input[32]), .Z(n7145) );
  XNOR U7153 ( .A(p_input[0]), .B(n7146), .Z(n6948) );
  AND U7154 ( .A(n303), .B(n7147), .Z(n7146) );
  XOR U7155 ( .A(p_input[16]), .B(p_input[0]), .Z(n7147) );
  XOR U7156 ( .A(n7148), .B(n7149), .Z(n303) );
  AND U7157 ( .A(n7150), .B(n7151), .Z(n7149) );
  XNOR U7158 ( .A(p_input[31]), .B(n7148), .Z(n7151) );
  XOR U7159 ( .A(n7148), .B(p_input[15]), .Z(n7150) );
  XOR U7160 ( .A(n7152), .B(n7153), .Z(n7148) );
  AND U7161 ( .A(n7154), .B(n7155), .Z(n7153) );
  XNOR U7162 ( .A(p_input[30]), .B(n7152), .Z(n7155) );
  XNOR U7163 ( .A(n7152), .B(n6962), .Z(n7154) );
  IV U7164 ( .A(p_input[14]), .Z(n6962) );
  XOR U7165 ( .A(n7156), .B(n7157), .Z(n7152) );
  AND U7166 ( .A(n7158), .B(n7159), .Z(n7157) );
  XNOR U7167 ( .A(p_input[29]), .B(n7156), .Z(n7159) );
  XNOR U7168 ( .A(n7156), .B(n6971), .Z(n7158) );
  IV U7169 ( .A(p_input[13]), .Z(n6971) );
  XOR U7170 ( .A(n7160), .B(n7161), .Z(n7156) );
  AND U7171 ( .A(n7162), .B(n7163), .Z(n7161) );
  XNOR U7172 ( .A(p_input[28]), .B(n7160), .Z(n7163) );
  XNOR U7173 ( .A(n7160), .B(n6980), .Z(n7162) );
  IV U7174 ( .A(p_input[12]), .Z(n6980) );
  XOR U7175 ( .A(n7164), .B(n7165), .Z(n7160) );
  AND U7176 ( .A(n7166), .B(n7167), .Z(n7165) );
  XNOR U7177 ( .A(p_input[27]), .B(n7164), .Z(n7167) );
  XNOR U7178 ( .A(n7164), .B(n6989), .Z(n7166) );
  IV U7179 ( .A(p_input[11]), .Z(n6989) );
  XOR U7180 ( .A(n7168), .B(n7169), .Z(n7164) );
  AND U7181 ( .A(n7170), .B(n7171), .Z(n7169) );
  XNOR U7182 ( .A(p_input[26]), .B(n7168), .Z(n7171) );
  XNOR U7183 ( .A(n7168), .B(n6998), .Z(n7170) );
  IV U7184 ( .A(p_input[10]), .Z(n6998) );
  XOR U7185 ( .A(n7172), .B(n7173), .Z(n7168) );
  AND U7186 ( .A(n7174), .B(n7175), .Z(n7173) );
  XNOR U7187 ( .A(p_input[25]), .B(n7172), .Z(n7175) );
  XNOR U7188 ( .A(n7172), .B(n7007), .Z(n7174) );
  IV U7189 ( .A(p_input[9]), .Z(n7007) );
  XOR U7190 ( .A(n7176), .B(n7177), .Z(n7172) );
  AND U7191 ( .A(n7178), .B(n7179), .Z(n7177) );
  XNOR U7192 ( .A(p_input[24]), .B(n7176), .Z(n7179) );
  XNOR U7193 ( .A(n7176), .B(n7016), .Z(n7178) );
  IV U7194 ( .A(p_input[8]), .Z(n7016) );
  XOR U7195 ( .A(n7180), .B(n7181), .Z(n7176) );
  AND U7196 ( .A(n7182), .B(n7183), .Z(n7181) );
  XNOR U7197 ( .A(p_input[23]), .B(n7180), .Z(n7183) );
  XNOR U7198 ( .A(n7180), .B(n7025), .Z(n7182) );
  IV U7199 ( .A(p_input[7]), .Z(n7025) );
  XOR U7200 ( .A(n7184), .B(n7185), .Z(n7180) );
  AND U7201 ( .A(n7186), .B(n7187), .Z(n7185) );
  XNOR U7202 ( .A(p_input[22]), .B(n7184), .Z(n7187) );
  XNOR U7203 ( .A(n7184), .B(n7034), .Z(n7186) );
  IV U7204 ( .A(p_input[6]), .Z(n7034) );
  XOR U7205 ( .A(n7188), .B(n7189), .Z(n7184) );
  AND U7206 ( .A(n7190), .B(n7191), .Z(n7189) );
  XNOR U7207 ( .A(p_input[21]), .B(n7188), .Z(n7191) );
  XNOR U7208 ( .A(n7188), .B(n7043), .Z(n7190) );
  IV U7209 ( .A(p_input[5]), .Z(n7043) );
  XOR U7210 ( .A(n7192), .B(n7193), .Z(n7188) );
  AND U7211 ( .A(n7194), .B(n7195), .Z(n7193) );
  XNOR U7212 ( .A(p_input[20]), .B(n7192), .Z(n7195) );
  XNOR U7213 ( .A(n7192), .B(n7052), .Z(n7194) );
  IV U7214 ( .A(p_input[4]), .Z(n7052) );
  XOR U7215 ( .A(n7196), .B(n7197), .Z(n7192) );
  AND U7216 ( .A(n7198), .B(n7199), .Z(n7197) );
  XNOR U7217 ( .A(p_input[19]), .B(n7196), .Z(n7199) );
  XNOR U7218 ( .A(n7196), .B(n7061), .Z(n7198) );
  IV U7219 ( .A(p_input[3]), .Z(n7061) );
  XOR U7220 ( .A(n7200), .B(n7201), .Z(n7196) );
  AND U7221 ( .A(n7202), .B(n7203), .Z(n7201) );
  XNOR U7222 ( .A(p_input[18]), .B(n7200), .Z(n7203) );
  XNOR U7223 ( .A(n7200), .B(n7070), .Z(n7202) );
  IV U7224 ( .A(p_input[2]), .Z(n7070) );
  XNOR U7225 ( .A(n7204), .B(n7205), .Z(n7200) );
  AND U7226 ( .A(n7206), .B(n7207), .Z(n7205) );
  XOR U7227 ( .A(p_input[17]), .B(n7204), .Z(n7207) );
  XNOR U7228 ( .A(p_input[1]), .B(n7204), .Z(n7206) );
  AND U7229 ( .A(p_input[16]), .B(n7208), .Z(n7204) );
  IV U7230 ( .A(p_input[0]), .Z(n7208) );
endmodule

